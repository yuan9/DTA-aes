
module aes_sbox_4 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559;

  OAI221X4 U28 ( .A0(n40), .A1(n553), .B0(n58), .B1(n547), .C0(n137), .Y(n136)
         );
  OAI221X4 U35 ( .A0(n145), .A1(n547), .B0(n28), .B1(n553), .C0(n146), .Y(n144) );
  OAI221X4 U38 ( .A0(n65), .A1(n553), .B0(n31), .B1(n539), .C0(n149), .Y(n143)
         );
  OAI221X4 U70 ( .A0(n46), .A1(n553), .B0(n63), .B1(n547), .C0(n200), .Y(n194)
         );
  OAI221X4 U103 ( .A0(n553), .A1(n87), .B0(n545), .B1(n104), .C0(n246), .Y(
        n235) );
  OAI221X4 U180 ( .A0(n553), .A1(n113), .B0(n88), .B1(n547), .C0(n320), .Y(
        n319) );
  OAI32X4 U188 ( .A0(n544), .A1(n63), .A2(n325), .B0(n37), .B1(n553), .Y(n324)
         );
  OAI221X4 U268 ( .A0(a[3]), .A1(n120), .B0(n201), .B1(n553), .C0(n363), .Y(
        n362) );
  NAND2X1 U1 ( .A(n56), .B(n535), .Y(n229) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X2 U3 ( .A(n66), .B(n71), .Y(n138) );
  AOI221XL U4 ( .A0(n559), .A1(n115), .B0(n554), .B1(n116), .C0(n117), .Y(n107) );
  AOI221X1 U5 ( .A0(n61), .A1(n556), .B0(n550), .B1(n147), .C0(n159), .Y(n153)
         );
  NAND2X2 U6 ( .A(n540), .B(n181), .Y(n113) );
  OAI221XL U7 ( .A0(n38), .A1(n539), .B0(n547), .B1(n183), .C0(n184), .Y(n176)
         );
  NAND2X2 U8 ( .A(a[3]), .B(n66), .Y(n181) );
  OAI221XL U9 ( .A0(n41), .A1(n547), .B0(n546), .B1(n181), .C0(n256), .Y(n255)
         );
  NAND2X1 U10 ( .A(n535), .B(n181), .Y(n102) );
  AOI221X1 U11 ( .A0(n551), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(n290) );
  NAND2X1 U12 ( .A(n536), .B(n75), .Y(n110) );
  NAND2X2 U13 ( .A(a[0]), .B(n26), .Y(n156) );
  NAND2X2 U14 ( .A(n75), .B(n26), .Y(n154) );
  NAND2X1 U15 ( .A(n39), .B(n535), .Y(n142) );
  NAND2X1 U16 ( .A(n535), .B(n542), .Y(n120) );
  NAND2X2 U17 ( .A(n66), .B(n538), .Y(n116) );
  OAI221XL U18 ( .A0(n43), .A1(n547), .B0(n546), .B1(n34), .C0(n365), .Y(n361)
         );
  AOI222X1 U19 ( .A0(n56), .A1(n543), .B0(n60), .B1(n555), .C0(n551), .C1(n71), 
        .Y(n356) );
  NAND2X1 U20 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U21 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI22XL U22 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  AOI22XL U23 ( .A0(n542), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  AOI222XL U24 ( .A0(n164), .A1(n550), .B0(a[2]), .B1(n227), .C0(n559), .C1(
        n228), .Y(n226) );
  AOI221XL U25 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357)
         );
  AOI33XL U26 ( .A0(a[3]), .A1(n543), .A2(n19), .B0(n185), .B1(n181), .B2(a[2]), .Y(n184) );
  CLKINVX3 U27 ( .A(a[2]), .Y(n73) );
  OAI222X4 U29 ( .A0(n546), .A1(n118), .B0(n119), .B1(n547), .C0(a[4]), .C1(
        n120), .Y(n117) );
  AOI21XL U30 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  NAND2X1 U31 ( .A(n535), .B(a[4]), .Y(n224) );
  NAND2X1 U32 ( .A(a[4]), .B(n538), .Y(n263) );
  CLKINVX3 U33 ( .A(a[4]), .Y(n66) );
  AOI22XL U34 ( .A0(n554), .A1(a[3]), .B0(n542), .B1(n66), .Y(n292) );
  NAND2X1 U36 ( .A(a[3]), .B(n538), .Y(n103) );
  NAND2X2 U37 ( .A(n535), .B(a[3]), .Y(n115) );
  NAND2XL U39 ( .A(n558), .B(a[3]), .Y(n259) );
  NAND2X2 U40 ( .A(a[3]), .B(a[4]), .Y(n111) );
  CLKINVX3 U41 ( .A(n539), .Y(n559) );
  CLKINVX3 U42 ( .A(n94), .Y(n543) );
  NAND2X1 U43 ( .A(n53), .B(n558), .Y(n288) );
  INVX1 U44 ( .A(n325), .Y(n34) );
  NOR2X1 U45 ( .A(n53), .B(n70), .Y(n326) );
  NAND2X1 U46 ( .A(n113), .B(n538), .Y(n214) );
  NOR2X1 U47 ( .A(n538), .B(n39), .Y(n325) );
  CLKINVX3 U48 ( .A(n557), .Y(n552) );
  NAND2X1 U49 ( .A(n56), .B(n538), .Y(n233) );
  NAND2X1 U50 ( .A(n46), .B(n538), .Y(n209) );
  NAND2X1 U51 ( .A(n138), .B(n538), .Y(n223) );
  NAND2X1 U52 ( .A(n50), .B(n538), .Y(n301) );
  NAND2X1 U53 ( .A(n541), .B(n268), .Y(n212) );
  NAND2X1 U54 ( .A(n39), .B(n538), .Y(n248) );
  INVX1 U55 ( .A(n102), .Y(n61) );
  NAND2X1 U56 ( .A(n147), .B(n214), .Y(n207) );
  INVX1 U57 ( .A(n541), .Y(n53) );
  INVX1 U58 ( .A(n168), .Y(n62) );
  INVX1 U59 ( .A(n182), .Y(n57) );
  INVX1 U60 ( .A(n116), .Y(n64) );
  INVX1 U61 ( .A(n230), .Y(n69) );
  CLKINVX3 U62 ( .A(n94), .Y(n542) );
  BUFX3 U63 ( .A(n74), .Y(n538) );
  NOR2X1 U64 ( .A(n540), .B(n538), .Y(n124) );
  NAND2X1 U65 ( .A(n50), .B(n535), .Y(n147) );
  NAND2X1 U66 ( .A(n538), .B(n71), .Y(n118) );
  CLKINVX3 U67 ( .A(n111), .Y(n39) );
  NAND2X1 U68 ( .A(n535), .B(n113), .Y(n165) );
  NAND2X1 U69 ( .A(n535), .B(n71), .Y(n230) );
  NAND2X1 U71 ( .A(n181), .B(n538), .Y(n166) );
  NAND2X1 U72 ( .A(n535), .B(n138), .Y(n182) );
  NAND2X1 U73 ( .A(n224), .B(n268), .Y(n141) );
  INVX1 U74 ( .A(n540), .Y(n46) );
  NAND2X1 U75 ( .A(n115), .B(n223), .Y(n306) );
  NAND2BX1 U76 ( .AN(n124), .B(n263), .Y(n196) );
  NAND2X1 U77 ( .A(n115), .B(n209), .Y(n210) );
  NAND2X1 U78 ( .A(n111), .B(n147), .Y(n96) );
  NAND2X1 U79 ( .A(n224), .B(n233), .Y(n104) );
  INVX1 U80 ( .A(n103), .Y(n68) );
  CLKINVX3 U81 ( .A(n536), .Y(n26) );
  CLKINVX3 U82 ( .A(n108), .Y(n22) );
  NAND2X1 U83 ( .A(n535), .B(n66), .Y(n337) );
  NAND2BX1 U84 ( .AN(n93), .B(n540), .Y(n299) );
  INVX1 U85 ( .A(n156), .Y(n24) );
  BUFX3 U86 ( .A(a[1]), .Y(n535) );
  OAI22X1 U87 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  NAND2X1 U88 ( .A(a[7]), .B(a[2]), .Y(n94) );
  NAND2X1 U89 ( .A(n536), .B(a[0]), .Y(n108) );
  NAND2X1 U90 ( .A(n59), .B(n543), .Y(n114) );
  INVX1 U91 ( .A(n238), .Y(n15) );
  INVX1 U92 ( .A(n326), .Y(n52) );
  INVX1 U93 ( .A(n288), .Y(n14) );
  CLKINVX3 U94 ( .A(n82), .Y(n558) );
  INVX1 U95 ( .A(n207), .Y(n48) );
  NOR2X1 U96 ( .A(n552), .B(n325), .Y(n199) );
  NOR2X1 U97 ( .A(n49), .B(n62), .Y(n247) );
  NOR2BX1 U98 ( .AN(n214), .B(n69), .Y(n88) );
  AOI22X1 U99 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  OAI221XL U100 ( .A0(n36), .A1(n552), .B0(n121), .B1(n544), .C0(n140), .Y(
        n135) );
  INVX1 U101 ( .A(n85), .Y(n36) );
  NOR2X1 U102 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U104 ( .A(n222), .B(n543), .Y(n162) );
  NAND2X1 U105 ( .A(n34), .B(n223), .Y(n183) );
  NAND2X1 U106 ( .A(n51), .B(n559), .Y(n238) );
  INVX1 U107 ( .A(n301), .Y(n49) );
  NAND2X1 U108 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U109 ( .A(n233), .Y(n55) );
  INVX1 U110 ( .A(n223), .Y(n59) );
  NOR2X1 U111 ( .A(n57), .B(n55), .Y(n197) );
  INVX1 U112 ( .A(n248), .Y(n37) );
  INVX1 U113 ( .A(n127), .Y(n35) );
  NOR2X1 U114 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U115 ( .A(n212), .Y(n41) );
  NOR2X1 U116 ( .A(n62), .B(n55), .Y(n145) );
  INVX1 U117 ( .A(n209), .Y(n45) );
  INVX1 U118 ( .A(n234), .Y(n54) );
  CLKINVX3 U119 ( .A(n113), .Y(n50) );
  CLKINVX8 U120 ( .A(n548), .Y(n547) );
  NAND2X1 U121 ( .A(n63), .B(n538), .Y(n243) );
  AOI22X1 U122 ( .A0(n347), .A1(n26), .B0(n558), .B1(n90), .Y(n343) );
  OAI221XL U123 ( .A0(n58), .A1(n547), .B0(n98), .B1(n545), .C0(n18), .Y(n347)
         );
  INVX1 U124 ( .A(n199), .Y(n18) );
  NOR2X1 U125 ( .A(n39), .B(n57), .Y(n179) );
  OAI22X1 U126 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U127 ( .A0(n559), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U128 ( .A0(n11), .A1(n538), .B0(n27), .B1(n559), .C0(n307), .Y(n302) );
  OAI22X1 U129 ( .A0(n64), .A1(n546), .B0(n552), .B1(n306), .Y(n304) );
  NAND2X1 U130 ( .A(n229), .B(n248), .Y(n87) );
  NOR2X1 U131 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U132 ( .A0(n94), .A1(n207), .B0(n547), .B1(n541), .Y(n242) );
  NAND3X1 U133 ( .A(n541), .B(n113), .C(n543), .Y(n89) );
  NAND2X1 U134 ( .A(n214), .B(n142), .Y(n90) );
  NAND2X1 U135 ( .A(n541), .B(n166), .Y(n311) );
  AOI22X1 U136 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U137 ( .A0(n98), .A1(n547), .B0(n30), .B1(n544), .C0(n99), .Y(n91)
         );
  OAI221XL U138 ( .A0(n42), .A1(n547), .B0(n51), .B1(n545), .C0(n95), .Y(n92)
         );
  INVX1 U139 ( .A(n104), .Y(n30) );
  NOR2BX1 U140 ( .AN(n229), .B(n68), .Y(n164) );
  NAND2X1 U141 ( .A(n558), .B(n96), .Y(n187) );
  AOI22X1 U142 ( .A0(n49), .A1(n549), .B0(n558), .B1(n141), .Y(n140) );
  AOI22X1 U143 ( .A0(n551), .A1(n34), .B0(n48), .B1(n542), .Y(n169) );
  OAI211X1 U144 ( .A0(n326), .A1(n552), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U145 ( .A0(n550), .A1(n63), .B0(n247), .B1(n542), .Y(n334) );
  OAI221XL U146 ( .A0(n35), .A1(n547), .B0(n44), .B1(n545), .C0(n333), .Y(n332) );
  AOI22X1 U147 ( .A0(n35), .A1(n558), .B0(n39), .B1(n554), .Y(n333) );
  AOI22X1 U148 ( .A0(n164), .A1(n558), .B0(n129), .B1(n556), .Y(n163) );
  AOI22X1 U149 ( .A0(n29), .A1(n558), .B0(n222), .B1(n549), .Y(n221) );
  AOI22X1 U150 ( .A0(n550), .A1(n311), .B0(n50), .B1(n542), .Y(n350) );
  NOR2X1 U151 ( .A(n138), .B(n539), .Y(n97) );
  NAND2X1 U152 ( .A(n243), .B(n142), .Y(n127) );
  NAND2X1 U153 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U154 ( .A(n138), .Y(n56) );
  NAND2X1 U155 ( .A(n229), .B(n209), .Y(n260) );
  INVX1 U156 ( .A(n118), .Y(n70) );
  INVX1 U157 ( .A(n120), .Y(n4) );
  NOR2X1 U158 ( .A(n64), .B(n124), .Y(n121) );
  AOI21X1 U159 ( .A0(n301), .A1(n337), .B0(n552), .Y(n336) );
  AND2X2 U160 ( .A(n165), .B(n166), .Y(n129) );
  NAND2X1 U161 ( .A(n541), .B(n214), .Y(n126) );
  OAI2BB2X1 U162 ( .B0(n547), .B1(n183), .A0N(n188), .A1N(n543), .Y(n335) );
  OAI31XL U163 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U164 ( .A0(n546), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U165 ( .A(n147), .Y(n47) );
  AOI221X1 U166 ( .A0(n126), .A1(n556), .B0(n127), .B1(n549), .C0(n128), .Y(
        n125) );
  OAI21XL U167 ( .A0(n539), .A1(n129), .B0(n130), .Y(n128) );
  OAI22X1 U168 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U169 ( .A0(n61), .A1(n549), .B0(n559), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U170 ( .A0(n559), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U171 ( .A(n116), .B(n229), .Y(n244) );
  AOI2BB2X1 U172 ( .B0(n11), .B1(n538), .A0N(n539), .A1N(n247), .Y(n246) );
  INVX1 U173 ( .A(n337), .Y(n65) );
  AOI22X1 U174 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  AOI2BB2X1 U175 ( .B0(n542), .B1(n87), .A0N(n547), .A1N(n121), .Y(n149) );
  OAI221XL U176 ( .A0(n31), .A1(n539), .B0(n553), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U177 ( .B0(n88), .B1(n542), .A0N(n547), .A1N(n197), .Y(n279) );
  INVX1 U178 ( .A(n166), .Y(n60) );
  INVX1 U179 ( .A(n208), .Y(n29) );
  INVX1 U181 ( .A(n299), .Y(n11) );
  NOR2X1 U182 ( .A(n547), .B(n538), .Y(n202) );
  INVX1 U183 ( .A(n100), .Y(n33) );
  INVX1 U184 ( .A(n228), .Y(n51) );
  OAI2BB1X1 U185 ( .A0N(n142), .A1N(n549), .B0(n187), .Y(n186) );
  AOI221XL U186 ( .A0(n550), .A1(n247), .B0(n212), .B1(n543), .C0(n266), .Y(
        n265) );
  OAI21XL U187 ( .A0(n165), .A1(n552), .B0(n187), .Y(n266) );
  NAND2BX1 U189 ( .AN(n97), .B(n206), .Y(n205) );
  OAI221XL U190 ( .A0(n539), .A1(n196), .B0(n197), .B1(n547), .C0(n198), .Y(
        n195) );
  AOI222X1 U191 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n543), 
        .Y(n198) );
  INVX1 U192 ( .A(n306), .Y(n58) );
  INVX1 U193 ( .A(n196), .Y(n31) );
  INVX1 U194 ( .A(n158), .Y(n42) );
  OAI221XL U195 ( .A0(n308), .A1(n553), .B0(n547), .B1(n165), .C0(n162), .Y(
        n307) );
  NOR2X1 U196 ( .A(n69), .B(n68), .Y(n308) );
  INVX1 U197 ( .A(n210), .Y(n44) );
  AOI211X1 U198 ( .A0(n554), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  INVX1 U199 ( .A(n141), .Y(n27) );
  INVX1 U200 ( .A(n96), .Y(n40) );
  INVX1 U201 ( .A(n148), .Y(n28) );
  CLKINVX3 U202 ( .A(n557), .Y(n553) );
  INVX1 U203 ( .A(n167), .Y(n32) );
  AOI31X1 U204 ( .A0(n102), .A1(n138), .A2(n559), .B0(n8), .Y(n137) );
  INVX1 U205 ( .A(n89), .Y(n8) );
  INVX1 U206 ( .A(n185), .Y(n19) );
  INVX1 U207 ( .A(n543), .Y(n544) );
  INVX1 U208 ( .A(n543), .Y(n545) );
  INVX1 U209 ( .A(n543), .Y(n546) );
  CLKINVX3 U210 ( .A(n110), .Y(n23) );
  NAND2X1 U211 ( .A(n116), .B(n142), .Y(n85) );
  INVX1 U212 ( .A(n154), .Y(n25) );
  OAI22X1 U213 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI211X1 U214 ( .A0(n39), .A1(n543), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U215 ( .A0(n553), .A1(n116), .B0(n73), .B1(n230), .C0(n547), .C1(
        n102), .Y(n275) );
  OAI21XL U216 ( .A0(n66), .A1(n552), .B0(n259), .Y(n257) );
  AOI221X1 U217 ( .A0(n56), .A1(n4), .B0(n551), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI221XL U218 ( .A0(n535), .A1(n259), .B0(n545), .B1(n214), .C0(n287), .Y(
        n293) );
  AOI31X1 U219 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI211X1 U220 ( .A0(n536), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  AOI22X1 U221 ( .A0(n536), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  AOI21X1 U222 ( .A0(n356), .A1(n357), .B0(n536), .Y(n355) );
  BUFX3 U223 ( .A(n82), .Y(n539) );
  NAND2X1 U224 ( .A(n73), .B(n20), .Y(n82) );
  AOI211X1 U225 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  INVX1 U226 ( .A(n284), .Y(n10) );
  OAI22X1 U227 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  OAI221XL U228 ( .A0(n67), .A1(n553), .B0(n546), .B1(n541), .C0(n294), .Y(
        n282) );
  AOI211X1 U229 ( .A0(n48), .A1(n559), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U230 ( .A(n114), .Y(n6) );
  AOI21X1 U231 ( .A0(n224), .A1(n243), .B0(n547), .Y(n295) );
  INVX1 U232 ( .A(n93), .Y(n548) );
  AOI22X1 U233 ( .A0(n348), .A1(n26), .B0(n536), .B1(n349), .Y(n342) );
  OAI221XL U234 ( .A0(n539), .A1(n166), .B0(n286), .B1(n547), .C0(n351), .Y(
        n348) );
  OAI211X1 U235 ( .A0(n88), .A1(n552), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U236 ( .B0(n542), .B1(n196), .A0N(n552), .A1N(n179), .Y(n351) );
  NAND2X1 U237 ( .A(n111), .B(n538), .Y(n268) );
  NAND2X1 U238 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U239 ( .A(n263), .B(n142), .Y(n100) );
  NAND2X1 U240 ( .A(n224), .B(n301), .Y(n148) );
  OAI21XL U241 ( .A0(n321), .A1(n539), .B0(n322), .Y(n318) );
  AOI31X1 U242 ( .A0(n541), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  OAI21XL U243 ( .A0(n73), .A1(n301), .B0(n552), .Y(n323) );
  CLKINVX3 U244 ( .A(n181), .Y(n63) );
  AOI21X1 U245 ( .A0(n539), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U246 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  NOR2BX1 U247 ( .AN(n263), .B(n61), .Y(n321) );
  AOI22X1 U248 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  OAI221XL U249 ( .A0(n66), .A1(n539), .B0(n61), .B1(n553), .C0(n84), .Y(n81)
         );
  OAI221XL U250 ( .A0(n86), .A1(n87), .B0(n88), .B1(n553), .C0(n89), .Y(n80)
         );
  AOI22X1 U251 ( .A0(n549), .A1(n85), .B0(n41), .B1(n542), .Y(n84) );
  NAND2X1 U252 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U253 ( .A0(n558), .A1(n66), .B0(n542), .B1(n147), .Y(n146) );
  AOI31X1 U254 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U255 ( .A0(n148), .A1(n73), .B0(n29), .B1(n556), .Y(n300) );
  OAI221XL U256 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  AOI222XL U257 ( .A0(n551), .A1(n210), .B0(n211), .B1(n212), .C0(n559), .C1(
        n540), .Y(n191) );
  AOI211X1 U258 ( .A0(n45), .A1(n543), .B0(n204), .C0(n205), .Y(n192) );
  AOI22X1 U259 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  AOI22X1 U260 ( .A0(n542), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  NAND2X1 U261 ( .A(n263), .B(n337), .Y(n167) );
  NAND2X1 U262 ( .A(n224), .B(n118), .Y(n208) );
  OAI21XL U263 ( .A0(n547), .A1(n540), .B0(n120), .Y(n276) );
  NAND2X1 U264 ( .A(n103), .B(n165), .Y(n188) );
  NAND2X1 U265 ( .A(n63), .B(n535), .Y(n168) );
  OAI21XL U266 ( .A0(n73), .A1(n214), .B0(n552), .Y(n211) );
  OAI21XL U267 ( .A0(n73), .A1(n243), .B0(n552), .Y(n245) );
  AOI21X1 U269 ( .A0(n263), .A1(n182), .B0(n547), .Y(n305) );
  INVX1 U270 ( .A(n535), .Y(n74) );
  NAND2X1 U271 ( .A(n558), .B(n535), .Y(n206) );
  XNOR2X1 U272 ( .A(n20), .B(n535), .Y(n185) );
  NAND2X1 U273 ( .A(n542), .B(n540), .Y(n130) );
  AOI21X1 U274 ( .A0(n90), .A1(n73), .B0(n559), .Y(n86) );
  AOI221X1 U275 ( .A0(n551), .A1(n111), .B0(n47), .B1(n543), .C0(n112), .Y(
        n109) );
  OAI221XL U276 ( .A0(n539), .A1(n113), .B0(n44), .B1(n553), .C0(n114), .Y(
        n112) );
  AOI221XL U277 ( .A0(n550), .A1(n230), .B0(n559), .B1(n126), .C0(n231), .Y(
        n225) );
  OAI22X1 U278 ( .A0(n35), .A1(n544), .B0(n552), .B1(n540), .Y(n231) );
  AOI21X1 U279 ( .A0(n558), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U280 ( .A0(n102), .A1(n103), .B0(n552), .Y(n101) );
  OAI221XL U281 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  AOI211X1 U282 ( .A0(n559), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  AOI211X1 U283 ( .A0(n543), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  AOI22X1 U284 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  AOI221X1 U285 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76)
         );
  OAI221XL U286 ( .A0(n539), .A1(n115), .B0(n121), .B1(n547), .C0(n122), .Y(
        n105) );
  INVX1 U287 ( .A(n125), .Y(n7) );
  OAI22X1 U288 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  XNOR2X1 U289 ( .A(n73), .B(n535), .Y(n161) );
  AOI211X1 U290 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U291 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI221XL U292 ( .A0(n54), .A1(n547), .B0(n33), .B1(n546), .C0(n232), .Y(n217) );
  OAI22X1 U293 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI211X1 U294 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  OAI22X1 U295 ( .A0(n544), .A1(n71), .B0(n37), .B1(n552), .Y(n157) );
  NAND2X1 U296 ( .A(n62), .B(n554), .Y(n287) );
  OAI221XL U297 ( .A0(n61), .A1(n553), .B0(n547), .B1(n260), .C0(n261), .Y(
        n254) );
  AOI21X1 U298 ( .A0(n33), .A1(n558), .B0(n262), .Y(n261) );
  AOI21X1 U299 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  OAI221XL U300 ( .A0(n63), .A1(n547), .B0(n546), .B1(n116), .C0(n178), .Y(
        n177) );
  AOI21X1 U301 ( .A0(n179), .A1(n555), .B0(n180), .Y(n178) );
  AOI21X1 U302 ( .A0(n181), .A1(n182), .B0(n539), .Y(n180) );
  INVX1 U303 ( .A(n260), .Y(n43) );
  AOI21X1 U304 ( .A0(n50), .A1(n558), .B0(n366), .Y(n365) );
  OAI32X1 U305 ( .A0(n553), .A1(n56), .A2(n53), .B0(n544), .B1(n103), .Y(n366)
         );
  AOI221X1 U306 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131) );
  OAI221XL U307 ( .A0(n56), .A1(n547), .B0(n32), .B1(n545), .C0(n163), .Y(n151) );
  OAI221XL U308 ( .A0(n539), .A1(n168), .B0(n164), .B1(n553), .C0(n169), .Y(
        n150) );
  OAI22X1 U309 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  OAI221XL U310 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  AOI221X1 U311 ( .A0(n559), .A1(n52), .B0(n550), .B1(n123), .C0(n324), .Y(
        n316) );
  AOI22X1 U312 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  AOI221X1 U313 ( .A0(n321), .A1(n554), .B0(n543), .B1(n311), .C0(n327), .Y(
        n315) );
  AOI211X1 U314 ( .A0(n201), .A1(n559), .B0(n202), .C0(n203), .Y(n200) );
  AOI21X1 U315 ( .A0(n111), .A1(n541), .B0(n545), .Y(n203) );
  OAI21XL U316 ( .A0(n539), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U317 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U318 ( .A(n162), .Y(n5) );
  NOR2BX1 U319 ( .AN(n263), .B(n47), .Y(n201) );
  OAI222X1 U320 ( .A0(n553), .A1(n207), .B0(n181), .B1(n120), .C0(n547), .C1(
        n208), .Y(n204) );
  OAI222X1 U321 ( .A0(n553), .A1(n167), .B0(n339), .B1(n539), .C0(n547), .C1(
        n34), .Y(n338) );
  AOI21X1 U322 ( .A0(n540), .A1(n538), .B0(n65), .Y(n339) );
  OAI221XL U323 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  AOI221X1 U324 ( .A0(n46), .A1(n543), .B0(n556), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI22X1 U325 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  AOI221X1 U326 ( .A0(n4), .A1(n71), .B0(n555), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI221XL U327 ( .A0(n539), .A1(n209), .B0(n547), .B1(n103), .C0(n288), .Y(
        n327) );
  OAI221XL U328 ( .A0(n547), .A1(n116), .B0(n321), .B1(n545), .C0(n359), .Y(
        n354) );
  AOI31X1 U329 ( .A0(n559), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  AOI21X1 U330 ( .A0(n115), .A1(n243), .B0(n552), .Y(n360) );
  BUFX3 U331 ( .A(n139), .Y(n541) );
  NAND2X1 U332 ( .A(n535), .B(n540), .Y(n139) );
  OAI2BB1X1 U333 ( .A0N(n223), .A1N(n224), .B0(n555), .Y(n220) );
  AOI32X1 U334 ( .A0(n34), .A1(n181), .A2(n559), .B0(n555), .B1(n233), .Y(n232) );
  AOI31X1 U335 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  AOI22X1 U336 ( .A0(n57), .A1(n548), .B0(n555), .B1(n113), .Y(n239) );
  AOI31X1 U337 ( .A0(n114), .A1(n206), .A2(n273), .B0(n536), .Y(n272) );
  AOI2BB2X1 U338 ( .B0(n70), .B1(n554), .A0N(n90), .A1N(n547), .Y(n273) );
  XOR2X1 U339 ( .A(n536), .B(n535), .Y(n358) );
  INVX1 U340 ( .A(n83), .Y(n557) );
  INVX1 U341 ( .A(n83), .Y(n554) );
  INVX1 U342 ( .A(n93), .Y(n551) );
  INVX1 U343 ( .A(n93), .Y(n550) );
  INVX1 U344 ( .A(n93), .Y(n549) );
  INVX1 U345 ( .A(n83), .Y(n555) );
  INVX1 U346 ( .A(n83), .Y(n556) );
  INVX1 U347 ( .A(n115), .Y(n67) );
  CLKINVX3 U348 ( .A(n537), .Y(n21) );
  OAI22X1 U349 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  AOI2BB2X1 U350 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  AOI22X1 U351 ( .A0(n536), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U352 ( .A0(n46), .A1(n553), .B0(n547), .B1(n116), .C0(n267), .Y(
        n264) );
  CLKINVX3 U353 ( .A(a[3]), .Y(n71) );
  OAI22X1 U354 ( .A0(n537), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  AOI211X1 U355 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  OAI22X1 U356 ( .A0(n340), .A1(n21), .B0(n537), .B1(n341), .Y(d[0]) );
  AOI22X1 U357 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  INVX1 U358 ( .A(n249), .Y(d[3]) );
  AOI22X1 U359 ( .A0(n250), .A1(n21), .B0(n537), .B1(n251), .Y(n249) );
  AOI22X1 U360 ( .A0(n536), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  AOI211X1 U361 ( .A0(n55), .A1(n559), .B0(n271), .C0(n272), .Y(n270) );
  OAI222X1 U362 ( .A0(n547), .A1(n141), .B0(n553), .B1(n263), .C0(n29), .C1(
        n544), .Y(n277) );
  AOI211X1 U363 ( .A0(n60), .A1(n543), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U364 ( .A(n547), .B(n39), .C(n61), .Y(n364) );
  INVX1 U365 ( .A(n259), .Y(n13) );
  BUFX3 U366 ( .A(n213), .Y(n540) );
  NAND2X1 U367 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U368 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U369 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U370 ( .A(n161), .Y(n72) );
  OAI2BB2X1 U371 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  NOR2X1 U372 ( .A(n549), .B(n556), .Y(n309) );
  OAI21XL U373 ( .A0(n537), .A1(n131), .B0(n132), .Y(d[6]) );
  OAI2BB1X1 U374 ( .A0N(n133), .A1N(n134), .B0(n537), .Y(n132) );
  OAI21XL U375 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  OAI2BB1X1 U376 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  OAI22X1 U377 ( .A0(n537), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  AOI211X1 U378 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  INVX1 U379 ( .A(n170), .Y(d[5]) );
  AOI22X1 U380 ( .A0(n171), .A1(n21), .B0(n537), .B1(n172), .Y(n170) );
  INVX1 U381 ( .A(n312), .Y(d[1]) );
  AOI22X1 U382 ( .A0(n537), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  NAND2X1 U383 ( .A(n138), .B(n102), .Y(n227) );
  OAI32X1 U384 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  NOR2X1 U385 ( .A(n60), .B(n62), .Y(n119) );
  AOI211X1 U386 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U387 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U388 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U389 ( .A(a[5]), .Y(n536) );
  INVX1 U390 ( .A(n87), .Y(n38) );
  CLKINVX3 U391 ( .A(a[0]), .Y(n75) );
  BUFX3 U392 ( .A(a[6]), .Y(n537) );
endmodule


module aes_sbox_3 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555;

  OAI221X4 U28 ( .A0(n40), .A1(n550), .B0(n58), .B1(n544), .C0(n137), .Y(n136)
         );
  OAI221X4 U35 ( .A0(n145), .A1(n544), .B0(n28), .B1(n550), .C0(n146), .Y(n144) );
  OAI221X4 U38 ( .A0(n65), .A1(n550), .B0(n31), .B1(n535), .C0(n149), .Y(n143)
         );
  OAI221X4 U70 ( .A0(n46), .A1(n550), .B0(n63), .B1(n544), .C0(n200), .Y(n194)
         );
  OAI221X4 U103 ( .A0(n550), .A1(n87), .B0(n540), .B1(n104), .C0(n246), .Y(
        n235) );
  OAI221X4 U166 ( .A0(n308), .A1(n550), .B0(n544), .B1(n165), .C0(n162), .Y(
        n307) );
  OAI221X4 U180 ( .A0(n550), .A1(n113), .B0(n88), .B1(n544), .C0(n320), .Y(
        n319) );
  OAI32X4 U188 ( .A0(n94), .A1(n63), .A2(n325), .B0(n37), .B1(n550), .Y(n324)
         );
  NAND2X4 U285 ( .A(a[3]), .B(n66), .Y(n181) );
  NAND2X2 U1 ( .A(n66), .B(n71), .Y(n138) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n56), .B(n531), .Y(n229) );
  NAND2X2 U4 ( .A(n536), .B(n181), .Y(n113) );
  OAI221XL U5 ( .A0(n41), .A1(n544), .B0(n542), .B1(n181), .C0(n256), .Y(n255)
         );
  NAND2X1 U6 ( .A(n531), .B(n181), .Y(n102) );
  NAND2X1 U7 ( .A(n532), .B(n75), .Y(n110) );
  NAND2X2 U8 ( .A(n66), .B(n534), .Y(n116) );
  NAND2X1 U9 ( .A(n39), .B(n531), .Y(n142) );
  OAI222X1 U10 ( .A0(n542), .A1(n118), .B0(n119), .B1(n544), .C0(a[4]), .C1(
        n120), .Y(n117) );
  AOI221XL U11 ( .A0(n4), .A1(n71), .B0(n553), .B1(n113), .C0(n186), .Y(n174)
         );
  AOI211X1 U12 ( .A0(n539), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  NAND2X2 U13 ( .A(a[0]), .B(n26), .Y(n156) );
  NAND2X2 U14 ( .A(n75), .B(n26), .Y(n154) );
  OAI221XL U15 ( .A0(a[3]), .A1(n120), .B0(n201), .B1(n550), .C0(n363), .Y(
        n362) );
  NAND2X1 U16 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U17 ( .A(a[7]), .B(n73), .Y(n93) );
  CLKINVX3 U18 ( .A(a[2]), .Y(n73) );
  AOI33X1 U19 ( .A0(a[3]), .A1(n539), .A2(n19), .B0(n185), .B1(n181), .B2(a[2]), .Y(n184) );
  AOI221X1 U20 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357)
         );
  AOI21XL U21 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  NAND2X1 U22 ( .A(n531), .B(a[4]), .Y(n224) );
  NAND2X1 U23 ( .A(a[4]), .B(n534), .Y(n263) );
  CLKINVX3 U24 ( .A(a[4]), .Y(n66) );
  AOI22XL U25 ( .A0(n553), .A1(a[3]), .B0(n538), .B1(n66), .Y(n292) );
  NAND2X1 U26 ( .A(a[3]), .B(n534), .Y(n103) );
  NAND2X2 U27 ( .A(n531), .B(a[3]), .Y(n115) );
  NAND2XL U29 ( .A(n16), .B(a[3]), .Y(n259) );
  NAND2X2 U30 ( .A(a[3]), .B(a[4]), .Y(n111) );
  CLKINVX3 U31 ( .A(n541), .Y(n539) );
  NAND2X1 U32 ( .A(n53), .B(n555), .Y(n288) );
  INVX1 U33 ( .A(n325), .Y(n34) );
  NOR2X1 U34 ( .A(n53), .B(n70), .Y(n326) );
  NAND2X1 U36 ( .A(n113), .B(n534), .Y(n214) );
  NOR2X1 U37 ( .A(n534), .B(n39), .Y(n325) );
  CLKINVX3 U39 ( .A(n554), .Y(n549) );
  CLKINVX3 U40 ( .A(n540), .Y(n538) );
  NAND2X1 U41 ( .A(n56), .B(n534), .Y(n233) );
  NAND2X1 U42 ( .A(n46), .B(n534), .Y(n209) );
  NAND2X1 U43 ( .A(n138), .B(n534), .Y(n223) );
  NAND2X1 U44 ( .A(n39), .B(n534), .Y(n248) );
  NAND2X1 U45 ( .A(n537), .B(n268), .Y(n212) );
  NAND2X1 U46 ( .A(n50), .B(n534), .Y(n301) );
  NAND2X1 U47 ( .A(n229), .B(n248), .Y(n87) );
  NAND2X1 U48 ( .A(n147), .B(n214), .Y(n207) );
  INVX1 U49 ( .A(n537), .Y(n53) );
  INVX1 U50 ( .A(n182), .Y(n57) );
  INVX1 U51 ( .A(n116), .Y(n64) );
  INVX1 U52 ( .A(n102), .Y(n61) );
  INVX1 U53 ( .A(n168), .Y(n62) );
  INVX1 U54 ( .A(n230), .Y(n69) );
  NOR2X1 U55 ( .A(n536), .B(n534), .Y(n124) );
  NAND2X1 U56 ( .A(n50), .B(n531), .Y(n147) );
  NAND2X1 U57 ( .A(n534), .B(n71), .Y(n118) );
  NAND2X1 U58 ( .A(n531), .B(n113), .Y(n165) );
  NAND2X1 U59 ( .A(n181), .B(n534), .Y(n166) );
  NAND2X1 U60 ( .A(n531), .B(n138), .Y(n182) );
  NAND2X1 U61 ( .A(n224), .B(n268), .Y(n141) );
  INVX1 U62 ( .A(n536), .Y(n46) );
  NAND2BX1 U63 ( .AN(n124), .B(n263), .Y(n196) );
  NAND2X1 U64 ( .A(n115), .B(n223), .Y(n306) );
  NAND2X1 U65 ( .A(n115), .B(n209), .Y(n210) );
  NAND2X1 U66 ( .A(n111), .B(n147), .Y(n96) );
  BUFX3 U67 ( .A(n74), .Y(n534) );
  NAND2X1 U68 ( .A(n263), .B(n142), .Y(n100) );
  INVX1 U69 ( .A(n103), .Y(n68) );
  CLKINVX3 U71 ( .A(n532), .Y(n26) );
  CLKINVX3 U72 ( .A(n111), .Y(n39) );
  NAND2X1 U73 ( .A(n531), .B(n71), .Y(n230) );
  CLKINVX3 U74 ( .A(n108), .Y(n22) );
  NAND2X1 U75 ( .A(n531), .B(n66), .Y(n337) );
  NAND2BX1 U76 ( .AN(n93), .B(n536), .Y(n299) );
  NAND2X1 U77 ( .A(n224), .B(n233), .Y(n104) );
  INVX1 U78 ( .A(n156), .Y(n24) );
  BUFX3 U79 ( .A(a[1]), .Y(n531) );
  NAND2X1 U80 ( .A(a[7]), .B(a[2]), .Y(n94) );
  NAND2X1 U81 ( .A(n532), .B(a[0]), .Y(n108) );
  NAND2X1 U82 ( .A(n59), .B(n539), .Y(n114) );
  INVX1 U83 ( .A(n238), .Y(n15) );
  INVX1 U84 ( .A(n326), .Y(n52) );
  INVX1 U85 ( .A(n288), .Y(n14) );
  NOR2X1 U86 ( .A(n549), .B(n325), .Y(n199) );
  NOR2X1 U87 ( .A(n49), .B(n62), .Y(n247) );
  NOR2BX1 U88 ( .AN(n214), .B(n69), .Y(n88) );
  AOI22X1 U89 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  OAI221XL U90 ( .A0(n36), .A1(n549), .B0(n121), .B1(n94), .C0(n140), .Y(n135)
         );
  INVX1 U91 ( .A(n85), .Y(n36) );
  NOR2X1 U92 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U93 ( .A(n222), .B(n539), .Y(n162) );
  NAND2X1 U94 ( .A(n34), .B(n223), .Y(n183) );
  NAND2X1 U95 ( .A(n51), .B(n555), .Y(n238) );
  INVX1 U96 ( .A(n301), .Y(n49) );
  INVX1 U97 ( .A(n233), .Y(n55) );
  INVX1 U98 ( .A(n223), .Y(n59) );
  NOR2X1 U99 ( .A(n57), .B(n55), .Y(n197) );
  INVX1 U100 ( .A(n248), .Y(n37) );
  INVX1 U101 ( .A(n127), .Y(n35) );
  INVX1 U102 ( .A(n207), .Y(n48) );
  INVX1 U104 ( .A(n212), .Y(n41) );
  INVX1 U105 ( .A(n87), .Y(n38) );
  INVX4 U106 ( .A(n535), .Y(n555) );
  NAND2X1 U107 ( .A(n34), .B(n248), .Y(n123) );
  NOR2X1 U108 ( .A(n59), .B(n69), .Y(n98) );
  NOR2X1 U109 ( .A(n62), .B(n55), .Y(n145) );
  INVX1 U110 ( .A(n209), .Y(n45) );
  NAND2X1 U111 ( .A(n63), .B(n534), .Y(n243) );
  NOR2X1 U112 ( .A(n39), .B(n57), .Y(n179) );
  OAI22X1 U113 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U114 ( .A0(n555), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U115 ( .A0(n11), .A1(n534), .B0(n27), .B1(n555), .C0(n307), .Y(n302) );
  OAI22X1 U116 ( .A0(n64), .A1(n542), .B0(n549), .B1(n306), .Y(n304) );
  NOR2X1 U117 ( .A(n46), .B(n57), .Y(n222) );
  CLKINVX3 U118 ( .A(n113), .Y(n50) );
  OAI22X1 U119 ( .A0(n541), .A1(n207), .B0(n544), .B1(n537), .Y(n242) );
  NAND3X1 U120 ( .A(n537), .B(n113), .C(n539), .Y(n89) );
  NAND2X1 U121 ( .A(n214), .B(n142), .Y(n90) );
  AOI22X1 U122 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U123 ( .A0(n98), .A1(n544), .B0(n30), .B1(n540), .C0(n99), .Y(n91)
         );
  OAI221XL U124 ( .A0(n42), .A1(n544), .B0(n51), .B1(n542), .C0(n95), .Y(n92)
         );
  INVX1 U125 ( .A(n104), .Y(n30) );
  NOR2BX1 U126 ( .AN(n229), .B(n68), .Y(n164) );
  NAND2X1 U127 ( .A(n555), .B(n96), .Y(n187) );
  AOI22X1 U128 ( .A0(n49), .A1(n547), .B0(n555), .B1(n141), .Y(n140) );
  AOI22X1 U129 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U130 ( .A0(n35), .A1(n544), .B0(n44), .B1(n542), .C0(n333), .Y(n332) );
  OAI211X1 U131 ( .A0(n326), .A1(n549), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U132 ( .A0(n35), .A1(n555), .B0(n39), .B1(n551), .Y(n333) );
  AOI22X1 U133 ( .A0(n548), .A1(n63), .B0(n247), .B1(n538), .Y(n334) );
  NOR2X1 U134 ( .A(n138), .B(n535), .Y(n97) );
  NAND2X1 U135 ( .A(n243), .B(n142), .Y(n127) );
  NAND2X1 U136 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U137 ( .A(n138), .Y(n56) );
  INVX1 U138 ( .A(n118), .Y(n70) );
  INVX1 U139 ( .A(n120), .Y(n4) );
  AND2X2 U140 ( .A(n165), .B(n166), .Y(n129) );
  NAND2X1 U141 ( .A(n537), .B(n214), .Y(n126) );
  NAND2X1 U142 ( .A(n138), .B(n102), .Y(n227) );
  INVX1 U143 ( .A(n284), .Y(n10) );
  OAI31XL U144 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U145 ( .A0(n540), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U146 ( .A(n147), .Y(n47) );
  OAI22X1 U147 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U148 ( .A0(n61), .A1(n546), .B0(n555), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U149 ( .A0(n555), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U150 ( .A(n116), .B(n229), .Y(n244) );
  AOI2BB2X1 U151 ( .B0(n11), .B1(n534), .A0N(n535), .A1N(n247), .Y(n246) );
  INVX1 U152 ( .A(n337), .Y(n65) );
  CLKINVX8 U153 ( .A(n545), .Y(n544) );
  AOI22X1 U154 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  AOI2BB2X1 U155 ( .B0(n538), .B1(n87), .A0N(n544), .A1N(n121), .Y(n149) );
  INVX1 U156 ( .A(n166), .Y(n60) );
  INVX1 U157 ( .A(n299), .Y(n11) );
  NOR2X1 U158 ( .A(n544), .B(n534), .Y(n202) );
  INVX1 U159 ( .A(n228), .Y(n51) );
  AOI221XL U160 ( .A0(n547), .A1(n247), .B0(n212), .B1(n539), .C0(n266), .Y(
        n265) );
  OAI21XL U161 ( .A0(n165), .A1(n549), .B0(n187), .Y(n266) );
  NAND2BX1 U162 ( .AN(n97), .B(n206), .Y(n205) );
  OAI221XL U163 ( .A0(n535), .A1(n196), .B0(n197), .B1(n544), .C0(n198), .Y(
        n195) );
  AOI222X1 U164 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n539), 
        .Y(n198) );
  NOR2X1 U165 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U167 ( .A0(n56), .A1(n544), .B0(n32), .B1(n540), .C0(n163), .Y(n151) );
  INVX1 U168 ( .A(n167), .Y(n32) );
  AOI22X1 U169 ( .A0(n164), .A1(n555), .B0(n129), .B1(n551), .Y(n163) );
  AOI211X1 U170 ( .A0(n555), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  AOI21X1 U171 ( .A0(n301), .A1(n337), .B0(n549), .Y(n336) );
  OAI2BB2X1 U172 ( .B0(n544), .B1(n183), .A0N(n188), .A1N(n539), .Y(n335) );
  INVX1 U173 ( .A(n210), .Y(n44) );
  OAI221XL U174 ( .A0(n535), .A1(n168), .B0(n164), .B1(n550), .C0(n169), .Y(
        n150) );
  AOI22X1 U175 ( .A0(n547), .A1(n34), .B0(n48), .B1(n538), .Y(n169) );
  AOI211X1 U176 ( .A0(n553), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  INVX1 U177 ( .A(n96), .Y(n40) );
  INVX1 U178 ( .A(n148), .Y(n28) );
  CLKINVX3 U179 ( .A(n554), .Y(n550) );
  AOI31X1 U181 ( .A0(n102), .A1(n138), .A2(n555), .B0(n8), .Y(n137) );
  INVX1 U182 ( .A(n89), .Y(n8) );
  INVX1 U183 ( .A(n185), .Y(n19) );
  INVX1 U184 ( .A(n543), .Y(n541) );
  INVX1 U185 ( .A(n125), .Y(n7) );
  AOI221X1 U186 ( .A0(n126), .A1(n551), .B0(n127), .B1(n548), .C0(n128), .Y(
        n125) );
  OAI21XL U187 ( .A0(n535), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U189 ( .A(n535), .Y(n16) );
  INVX1 U190 ( .A(n539), .Y(n542) );
  AOI22X1 U191 ( .A0(n347), .A1(n26), .B0(n16), .B1(n90), .Y(n343) );
  OAI221XL U192 ( .A0(n58), .A1(n544), .B0(n98), .B1(n94), .C0(n18), .Y(n347)
         );
  INVX1 U193 ( .A(n199), .Y(n18) );
  CLKINVX3 U194 ( .A(n110), .Y(n23) );
  NAND2X1 U195 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U196 ( .A(n537), .B(n166), .Y(n311) );
  AOI22X1 U197 ( .A0(n546), .A1(n311), .B0(n50), .B1(n538), .Y(n350) );
  INVX1 U198 ( .A(n154), .Y(n25) );
  NAND2X1 U199 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U200 ( .A(n64), .B(n124), .Y(n121) );
  INVX1 U201 ( .A(n208), .Y(n29) );
  INVX1 U202 ( .A(n100), .Y(n33) );
  INVX1 U203 ( .A(n306), .Y(n58) );
  INVX1 U204 ( .A(n196), .Y(n31) );
  INVX1 U205 ( .A(n158), .Y(n42) );
  INVX1 U206 ( .A(n141), .Y(n27) );
  NAND2X2 U207 ( .A(n531), .B(n538), .Y(n120) );
  AOI22X1 U208 ( .A0(n348), .A1(n26), .B0(n532), .B1(n349), .Y(n342) );
  OAI221XL U209 ( .A0(n535), .A1(n166), .B0(n286), .B1(n544), .C0(n351), .Y(
        n348) );
  OAI211X1 U210 ( .A0(n88), .A1(n549), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U211 ( .B0(n538), .B1(n196), .A0N(n549), .A1N(n179), .Y(n351) );
  AOI22X1 U212 ( .A0(n532), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U213 ( .A0(n544), .A1(n141), .B0(n550), .B1(n263), .C0(n29), .C1(
        n541), .Y(n277) );
  OAI221XL U214 ( .A0(n31), .A1(n535), .B0(n550), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U215 ( .B0(n88), .B1(n538), .A0N(n544), .A1N(n197), .Y(n279) );
  OAI22X1 U216 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U217 ( .A0(n547), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U218 ( .A0(n56), .A1(n4), .B0(n546), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U219 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U220 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U221 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U222 ( .A0(n61), .A1(n552), .B0(n546), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U223 ( .A0(n541), .A1(n71), .B0(n37), .B1(n549), .Y(n157) );
  NAND2X1 U224 ( .A(n111), .B(n534), .Y(n268) );
  OAI22X1 U225 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U226 ( .A0(n547), .A1(n111), .B0(n47), .B1(n539), .C0(n112), .Y(
        n109) );
  AOI221X1 U227 ( .A0(n555), .A1(n115), .B0(n553), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U228 ( .A0(n535), .A1(n113), .B0(n44), .B1(n550), .C0(n114), .Y(
        n112) );
  NAND2X1 U229 ( .A(n224), .B(n301), .Y(n148) );
  OAI21XL U230 ( .A0(n321), .A1(n535), .B0(n322), .Y(n318) );
  AOI31X1 U231 ( .A0(n537), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  OAI21XL U232 ( .A0(n73), .A1(n301), .B0(n549), .Y(n323) );
  CLKINVX3 U233 ( .A(n181), .Y(n63) );
  NOR2BX1 U234 ( .AN(n263), .B(n61), .Y(n321) );
  AOI22X1 U235 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  OAI221XL U236 ( .A0(n66), .A1(n535), .B0(n61), .B1(n550), .C0(n84), .Y(n81)
         );
  OAI221XL U237 ( .A0(n86), .A1(n87), .B0(n88), .B1(n550), .C0(n89), .Y(n80)
         );
  AOI22X1 U238 ( .A0(n546), .A1(n85), .B0(n41), .B1(n538), .Y(n84) );
  NAND2X1 U239 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U240 ( .A0(n555), .A1(n66), .B0(n538), .B1(n147), .Y(n146) );
  OAI221XL U241 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  AOI222X1 U242 ( .A0(n547), .A1(n210), .B0(n211), .B1(n212), .C0(n555), .C1(
        n536), .Y(n191) );
  AOI211X1 U243 ( .A0(n45), .A1(n539), .B0(n204), .C0(n205), .Y(n192) );
  AOI22X1 U244 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  AOI22X1 U245 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U246 ( .A0(n63), .A1(n544), .B0(n542), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U247 ( .A0(n38), .A1(n535), .B0(n544), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U248 ( .A0(n179), .A1(n551), .B0(n180), .Y(n178) );
  NAND2X1 U249 ( .A(n263), .B(n337), .Y(n167) );
  NAND2X1 U250 ( .A(n224), .B(n118), .Y(n208) );
  OAI21XL U251 ( .A0(n544), .A1(n536), .B0(n120), .Y(n276) );
  NAND2X1 U252 ( .A(n103), .B(n165), .Y(n188) );
  NAND2X1 U253 ( .A(n63), .B(n531), .Y(n168) );
  AOI21X1 U254 ( .A0(n224), .A1(n243), .B0(n544), .Y(n295) );
  OAI21XL U255 ( .A0(n73), .A1(n214), .B0(n549), .Y(n211) );
  OAI21XL U256 ( .A0(n73), .A1(n243), .B0(n549), .Y(n245) );
  AOI21X1 U257 ( .A0(n263), .A1(n182), .B0(n544), .Y(n305) );
  INVX1 U258 ( .A(n531), .Y(n74) );
  OAI21XL U259 ( .A0(n66), .A1(n549), .B0(n259), .Y(n257) );
  NAND2X1 U260 ( .A(n555), .B(n531), .Y(n206) );
  XNOR2X1 U261 ( .A(n20), .B(n531), .Y(n185) );
  NAND2X1 U262 ( .A(n538), .B(n536), .Y(n130) );
  AOI21X1 U263 ( .A0(n90), .A1(n73), .B0(n555), .Y(n86) );
  AOI21X1 U264 ( .A0(n16), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U265 ( .A0(n102), .A1(n103), .B0(n549), .Y(n101) );
  AOI211X1 U266 ( .A0(n39), .A1(n539), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U267 ( .A0(n550), .A1(n116), .B0(n73), .B1(n230), .C0(n544), .C1(
        n102), .Y(n275) );
  XNOR2X1 U268 ( .A(n73), .B(n531), .Y(n161) );
  AOI211X1 U269 ( .A0(n55), .A1(n555), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U270 ( .A0(n114), .A1(n206), .A2(n273), .B0(n532), .Y(n272) );
  OAI22X1 U271 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U272 ( .B0(n70), .B1(n551), .A0N(n90), .A1N(n544), .Y(n273) );
  NAND2X1 U273 ( .A(n62), .B(n553), .Y(n287) );
  OAI221XL U274 ( .A0(n61), .A1(n550), .B0(n544), .B1(n260), .C0(n261), .Y(
        n254) );
  AOI21X1 U275 ( .A0(n33), .A1(n555), .B0(n262), .Y(n261) );
  AOI21X1 U276 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI21X1 U277 ( .A0(n50), .A1(n16), .B0(n366), .Y(n365) );
  OAI32X1 U278 ( .A0(n550), .A1(n56), .A2(n53), .B0(n94), .B1(n103), .Y(n366)
         );
  OAI221XL U279 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  AOI221XL U280 ( .A0(n555), .A1(n52), .B0(n548), .B1(n123), .C0(n324), .Y(
        n316) );
  AOI22X1 U281 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  AOI221X1 U282 ( .A0(n321), .A1(n552), .B0(n539), .B1(n311), .C0(n327), .Y(
        n315) );
  AOI211X1 U283 ( .A0(n201), .A1(n555), .B0(n202), .C0(n203), .Y(n200) );
  AOI21X1 U284 ( .A0(n111), .A1(n537), .B0(n540), .Y(n203) );
  OAI21XL U286 ( .A0(n535), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U287 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U288 ( .A(n162), .Y(n5) );
  NOR2BX1 U289 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U290 ( .A(n82), .Y(n535) );
  NAND2X1 U291 ( .A(n73), .B(n20), .Y(n82) );
  OAI222X1 U292 ( .A0(n550), .A1(n207), .B0(n181), .B1(n120), .C0(n544), .C1(
        n208), .Y(n204) );
  OAI222X1 U293 ( .A0(n550), .A1(n167), .B0(n339), .B1(n535), .C0(n544), .C1(
        n34), .Y(n338) );
  AOI21X1 U294 ( .A0(n536), .A1(n534), .B0(n65), .Y(n339) );
  OAI2BB1X1 U295 ( .A0N(n142), .A1N(n548), .B0(n187), .Y(n186) );
  AOI221X1 U296 ( .A0(n46), .A1(n539), .B0(n552), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U297 ( .A0(n535), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U298 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  OAI221XL U299 ( .A0(n535), .A1(n209), .B0(n544), .B1(n103), .C0(n288), .Y(
        n327) );
  OAI221XL U300 ( .A0(n531), .A1(n259), .B0(n94), .B1(n214), .C0(n287), .Y(
        n293) );
  OAI221XL U301 ( .A0(n54), .A1(n544), .B0(n33), .B1(n94), .C0(n232), .Y(n217)
         );
  INVX1 U302 ( .A(n234), .Y(n54) );
  AOI32X1 U303 ( .A0(n34), .A1(n181), .A2(n555), .B0(n551), .B1(n233), .Y(n232) );
  BUFX3 U304 ( .A(n139), .Y(n537) );
  NAND2X1 U305 ( .A(n531), .B(n536), .Y(n139) );
  AOI211X1 U306 ( .A0(n60), .A1(n539), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U307 ( .A(n544), .B(n39), .C(n61), .Y(n364) );
  INVX1 U308 ( .A(n259), .Y(n13) );
  OAI221XL U309 ( .A0(n67), .A1(n550), .B0(n542), .B1(n537), .C0(n294), .Y(
        n282) );
  INVX1 U310 ( .A(n115), .Y(n67) );
  AOI211X1 U311 ( .A0(n48), .A1(n555), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U312 ( .A(n114), .Y(n6) );
  AOI211X1 U313 ( .A0(n532), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  AOI21X1 U314 ( .A0(n356), .A1(n357), .B0(n532), .Y(n355) );
  OAI221XL U315 ( .A0(n544), .A1(n116), .B0(n321), .B1(n540), .C0(n359), .Y(
        n354) );
  AOI222X1 U316 ( .A0(n56), .A1(n539), .B0(n60), .B1(n553), .C0(n548), .C1(n71), .Y(n356) );
  AOI31X1 U317 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U318 ( .A0N(n223), .A1N(n224), .B0(n552), .Y(n220) );
  AOI22X1 U319 ( .A0(n29), .A1(n16), .B0(n222), .B1(n548), .Y(n221) );
  AOI31X1 U320 ( .A0(n555), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  AOI21X1 U321 ( .A0(n115), .A1(n243), .B0(n549), .Y(n360) );
  AOI31X1 U322 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  AOI22X1 U323 ( .A0(n57), .A1(n545), .B0(n552), .B1(n113), .Y(n239) );
  AOI31X1 U324 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U325 ( .A0(n148), .A1(n73), .B0(n29), .B1(n552), .Y(n300) );
  INVX1 U326 ( .A(n83), .Y(n553) );
  INVX1 U327 ( .A(n93), .Y(n545) );
  INVX1 U328 ( .A(n543), .Y(n540) );
  INVX1 U329 ( .A(n94), .Y(n543) );
  INVX1 U330 ( .A(n83), .Y(n554) );
  INVX1 U331 ( .A(n93), .Y(n546) );
  INVX1 U332 ( .A(n93), .Y(n547) );
  INVX1 U333 ( .A(n93), .Y(n548) );
  NAND2X1 U334 ( .A(n115), .B(n268), .Y(n158) );
  AOI21X1 U335 ( .A0(n181), .A1(n182), .B0(n535), .Y(n180) );
  AOI22X1 U336 ( .A0(n538), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  XOR2X1 U337 ( .A(n532), .B(n531), .Y(n358) );
  INVX1 U338 ( .A(n83), .Y(n551) );
  INVX1 U339 ( .A(n83), .Y(n552) );
  CLKINVX3 U340 ( .A(n533), .Y(n21) );
  OAI22X1 U341 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  AOI2BB2X1 U342 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  AOI22X1 U343 ( .A0(n532), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U344 ( .A0(n46), .A1(n550), .B0(n544), .B1(n116), .C0(n267), .Y(
        n264) );
  CLKINVX3 U345 ( .A(a[3]), .Y(n71) );
  OAI22X1 U346 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U347 ( .A0(n548), .A1(n230), .B0(n555), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U348 ( .A0(n164), .A1(n546), .B0(a[2]), .B1(n227), .C0(n555), .C1(
        n228), .Y(n226) );
  OAI22X1 U349 ( .A0(n35), .A1(n541), .B0(n549), .B1(n536), .Y(n231) );
  OAI22X1 U350 ( .A0(n340), .A1(n21), .B0(n533), .B1(n341), .Y(d[0]) );
  AOI22X1 U351 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U352 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  OAI22X1 U353 ( .A0(n533), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  AOI211X1 U354 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U355 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  OAI22X1 U356 ( .A0(n533), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  AOI211X1 U357 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U358 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI21XL U359 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  OAI2BB1X1 U360 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI221X1 U361 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76)
         );
  INVX1 U362 ( .A(n312), .Y(d[1]) );
  AOI22X1 U363 ( .A0(n533), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U364 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  INVX1 U365 ( .A(n249), .Y(d[3]) );
  AOI22X1 U366 ( .A0(n250), .A1(n21), .B0(n533), .B1(n251), .Y(n249) );
  OAI22X1 U367 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  INVX1 U368 ( .A(n170), .Y(d[5]) );
  AOI22X1 U369 ( .A0(n171), .A1(n21), .B0(n533), .B1(n172), .Y(n170) );
  OAI221XL U370 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  AOI22X1 U371 ( .A0(n532), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U372 ( .A0(n43), .A1(n544), .B0(n542), .B1(n34), .C0(n365), .Y(n361) );
  INVX1 U373 ( .A(n260), .Y(n43) );
  OAI21XL U374 ( .A0(n533), .A1(n131), .B0(n132), .Y(d[6]) );
  OAI2BB1X1 U375 ( .A0N(n133), .A1N(n134), .B0(n533), .Y(n132) );
  AOI221X1 U376 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n536) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI221XL U383 ( .A0(n535), .A1(n115), .B0(n121), .B1(n544), .C0(n122), .Y(
        n105) );
  AOI22X1 U384 ( .A0(n538), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  OAI2BB2X1 U385 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  NOR2X1 U386 ( .A(n547), .B(n553), .Y(n309) );
  AOI22X1 U387 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U388 ( .A(a[0]), .Y(n75) );
  AOI211X1 U389 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U390 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U391 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U392 ( .A(a[5]), .Y(n532) );
  BUFX3 U393 ( .A(a[6]), .Y(n533) );
endmodule


module aes_rcon ( clk, kld, out );
  output [31:0] out;
  input clk, kld;
  wire   N44, N45, N46, N47, N48, N49, N51, N55, n14, n6, n7, n8, n9, n11, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n32, n33, n34;
  wire   [3:0] rcnt;
  assign out[0] = 1'b0;
  assign out[1] = 1'b0;
  assign out[2] = 1'b0;
  assign out[3] = 1'b0;
  assign out[4] = 1'b0;
  assign out[5] = 1'b0;
  assign out[6] = 1'b0;
  assign out[7] = 1'b0;
  assign out[8] = 1'b0;
  assign out[9] = 1'b0;
  assign out[10] = 1'b0;
  assign out[11] = 1'b0;
  assign out[12] = 1'b0;
  assign out[13] = 1'b0;
  assign out[14] = 1'b0;
  assign out[15] = 1'b0;
  assign out[16] = 1'b0;
  assign out[17] = 1'b0;
  assign out[18] = 1'b0;
  assign out[19] = 1'b0;
  assign out[20] = 1'b0;
  assign out[21] = 1'b0;
  assign out[22] = 1'b0;
  assign out[23] = 1'b0;

  DFFTRX1 \out_reg[30]  ( .D(n14), .RN(n7), .CK(clk), .Q(out[30]) );
  DFFHQX1 \out_reg[24]  ( .D(N44), .CK(clk), .Q(out[24]) );
  DFFHQX1 \out_reg[31]  ( .D(N51), .CK(clk), .Q(out[31]) );
  DFFHQX1 \out_reg[27]  ( .D(N47), .CK(clk), .Q(out[27]) );
  DFFHQX1 \out_reg[26]  ( .D(N46), .CK(clk), .Q(out[26]) );
  DFFHQX1 \out_reg[25]  ( .D(N45), .CK(clk), .Q(out[25]) );
  DFFHQX1 \out_reg[29]  ( .D(N49), .CK(clk), .Q(out[29]) );
  DFFHQX1 \out_reg[28]  ( .D(N48), .CK(clk), .Q(out[28]) );
  DFFTRX1 \rcnt_reg[1]  ( .D(n14), .RN(n34), .CK(clk), .Q(rcnt[1]) );
  DFFX1 \rcnt_reg[3]  ( .D(N55), .CK(clk), .Q(n30), .QN(n11) );
  DFFTRX1 \rcnt_reg[2]  ( .D(n8), .RN(n34), .CK(clk), .Q(rcnt[2]), .QN(n33) );
  JKFFX1 \rcnt_reg[0]  ( .J(n34), .K(1'b1), .CK(clk), .Q(rcnt[0]), .QN(n32) );
  XOR2X1 U3 ( .A(rcnt[1]), .B(rcnt[0]), .Y(n14) );
  NAND4X1 U4 ( .A(n22), .B(rcnt[0]), .C(n8), .D(n34), .Y(n15) );
  INVX1 U5 ( .A(kld), .Y(n34) );
  NOR2X1 U6 ( .A(n22), .B(n14), .Y(n21) );
  OAI21XL U7 ( .A0(n9), .A1(n33), .B0(n25), .Y(n27) );
  INVX1 U8 ( .A(n14), .Y(n9) );
  NAND3X1 U9 ( .A(n14), .B(n32), .C(n22), .Y(n17) );
  NAND2X1 U10 ( .A(n18), .B(n34), .Y(n20) );
  OAI22X1 U11 ( .A0(n14), .A1(n15), .B0(n6), .B1(n20), .Y(N48) );
  INVX1 U12 ( .A(n21), .Y(n6) );
  NAND4X1 U13 ( .A(n28), .B(n27), .C(n34), .D(n11), .Y(n16) );
  NOR3X1 U14 ( .A(n17), .B(kld), .C(n18), .Y(N51) );
  OAI21XL U15 ( .A0(N44), .A1(n11), .B0(n16), .Y(N55) );
  OAI2BB1X1 U16 ( .A0N(n27), .A1N(n28), .B0(n34), .Y(N44) );
  INVX1 U17 ( .A(n18), .Y(n8) );
  INVX1 U18 ( .A(n15), .Y(n7) );
  OAI31X1 U19 ( .A0(n27), .A1(kld), .A2(n28), .B0(n16), .Y(N45) );
  NAND2X1 U20 ( .A(rcnt[1]), .B(rcnt[0]), .Y(n25) );
  NOR4BX1 U21 ( .AN(n19), .B(rcnt[0]), .C(kld), .D(n14), .Y(N49) );
  XOR2X1 U22 ( .A(rcnt[2]), .B(n30), .Y(n19) );
  XOR2X1 U23 ( .A(n25), .B(rcnt[2]), .Y(n18) );
  XNOR2X1 U24 ( .A(n30), .B(n26), .Y(n22) );
  NOR2X1 U25 ( .A(n25), .B(n33), .Y(n26) );
  AOI21X1 U26 ( .A0(n17), .A1(n23), .B0(n20), .Y(N47) );
  NAND2X1 U27 ( .A(n21), .B(rcnt[0]), .Y(n23) );
  XNOR2X1 U28 ( .A(n32), .B(n29), .Y(n28) );
  XOR2X1 U29 ( .A(rcnt[2]), .B(rcnt[1]), .Y(n29) );
  NOR2X1 U30 ( .A(n24), .B(n20), .Y(N46) );
  AOI32X1 U31 ( .A0(rcnt[0]), .A1(n14), .A2(n22), .B0(n21), .B1(n32), .Y(n24)
         );
endmodule


module aes_sbox_1 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915;

  OAI221X4 U28 ( .A0(n882), .A1(n550), .B0(n864), .B1(n544), .C0(n785), .Y(
        n786) );
  OAI221X4 U35 ( .A0(n777), .A1(n544), .B0(n894), .B1(n550), .C0(n776), .Y(
        n778) );
  OAI221X4 U38 ( .A0(n857), .A1(n550), .B0(n891), .B1(n535), .C0(n773), .Y(
        n779) );
  OAI221X4 U70 ( .A0(n876), .A1(n550), .B0(n859), .B1(n544), .C0(n722), .Y(
        n728) );
  OAI221X4 U103 ( .A0(n550), .A1(n835), .B0(n540), .B1(n818), .C0(n676), .Y(
        n687) );
  OAI221X4 U166 ( .A0(n614), .A1(n550), .B0(n544), .B1(n757), .C0(n760), .Y(
        n615) );
  OAI221X4 U180 ( .A0(n550), .A1(n809), .B0(n834), .B1(n544), .C0(n602), .Y(
        n603) );
  OAI32X4 U188 ( .A0(n828), .A1(n859), .A2(n597), .B0(n885), .B1(n550), .Y(
        n598) );
  NAND2X4 U285 ( .A(a[3]), .B(n856), .Y(n741) );
  NAND2X2 U1 ( .A(n856), .B(n851), .Y(n784) );
  INVX1 U2 ( .A(a[7]), .Y(n902) );
  NAND2X1 U3 ( .A(n866), .B(n531), .Y(n693) );
  NAND2X2 U4 ( .A(n536), .B(n741), .Y(n809) );
  OAI221XL U5 ( .A0(n881), .A1(n544), .B0(n542), .B1(n741), .C0(n666), .Y(n667) );
  NAND2X1 U6 ( .A(n531), .B(n741), .Y(n820) );
  NAND2X1 U7 ( .A(n532), .B(n847), .Y(n812) );
  NAND2X2 U8 ( .A(n856), .B(n534), .Y(n806) );
  NAND2X1 U9 ( .A(n883), .B(n531), .Y(n780) );
  OAI222X1 U10 ( .A0(n542), .A1(n804), .B0(n803), .B1(n544), .C0(a[4]), .C1(
        n802), .Y(n805) );
  AOI221XL U11 ( .A0(n915), .A1(n851), .B0(n551), .B1(n809), .C0(n736), .Y(
        n748) );
  AOI211X1 U12 ( .A0(n539), .A1(n851), .B0(n584), .C0(n646), .Y(n594) );
  NAND2X2 U13 ( .A(a[0]), .B(n896), .Y(n766) );
  NAND2X2 U14 ( .A(n847), .B(n896), .Y(n768) );
  OAI221XL U15 ( .A0(a[3]), .A1(n802), .B0(n721), .B1(n550), .C0(n559), .Y(
        n560) );
  NAND2X1 U16 ( .A(a[2]), .B(n902), .Y(n839) );
  NAND2X1 U17 ( .A(a[7]), .B(n849), .Y(n829) );
  CLKINVX3 U18 ( .A(a[2]), .Y(n849) );
  AOI33X1 U19 ( .A0(a[3]), .A1(n539), .A2(n903), .B0(n737), .B1(n741), .B2(
        a[2]), .Y(n738) );
  AOI221X1 U20 ( .A0(n857), .A1(a[2]), .B0(n825), .B1(n564), .C0(n915), .Y(
        n565) );
  AOI21XL U21 ( .A0(n915), .A1(a[4]), .B0(n906), .Y(n602) );
  NAND2X1 U22 ( .A(n531), .B(a[4]), .Y(n698) );
  NAND2X1 U23 ( .A(a[4]), .B(n534), .Y(n659) );
  CLKINVX3 U24 ( .A(a[4]), .Y(n856) );
  AOI22XL U25 ( .A0(n551), .A1(a[3]), .B0(n538), .B1(n856), .Y(n630) );
  NAND2X1 U26 ( .A(a[3]), .B(n534), .Y(n819) );
  NAND2X2 U27 ( .A(n531), .B(a[3]), .Y(n807) );
  NAND2XL U29 ( .A(n905), .B(a[3]), .Y(n663) );
  NAND2X2 U30 ( .A(a[3]), .B(a[4]), .Y(n811) );
  CLKINVX3 U31 ( .A(n541), .Y(n539) );
  NAND2X1 U32 ( .A(n869), .B(n555), .Y(n634) );
  INVX1 U33 ( .A(n597), .Y(n888) );
  NOR2X1 U34 ( .A(n869), .B(n852), .Y(n596) );
  NAND2X1 U36 ( .A(n809), .B(n534), .Y(n708) );
  NOR2X1 U37 ( .A(n534), .B(n883), .Y(n597) );
  CLKINVX3 U39 ( .A(n554), .Y(n549) );
  CLKINVX3 U40 ( .A(n540), .Y(n538) );
  NAND2X1 U41 ( .A(n866), .B(n534), .Y(n689) );
  NAND2X1 U42 ( .A(n876), .B(n534), .Y(n713) );
  NAND2X1 U43 ( .A(n784), .B(n534), .Y(n699) );
  NAND2X1 U44 ( .A(n883), .B(n534), .Y(n674) );
  NAND2X1 U45 ( .A(n537), .B(n654), .Y(n710) );
  NAND2X1 U46 ( .A(n872), .B(n534), .Y(n621) );
  NAND2X1 U47 ( .A(n693), .B(n674), .Y(n835) );
  NAND2X1 U48 ( .A(n775), .B(n708), .Y(n715) );
  INVX1 U49 ( .A(n537), .Y(n869) );
  INVX1 U50 ( .A(n740), .Y(n865) );
  INVX1 U51 ( .A(n806), .Y(n858) );
  INVX1 U52 ( .A(n820), .Y(n861) );
  INVX1 U53 ( .A(n754), .Y(n860) );
  INVX1 U54 ( .A(n692), .Y(n853) );
  NOR2X1 U55 ( .A(n536), .B(n534), .Y(n798) );
  NAND2X1 U56 ( .A(n872), .B(n531), .Y(n775) );
  NAND2X1 U57 ( .A(n534), .B(n851), .Y(n804) );
  NAND2X1 U58 ( .A(n531), .B(n809), .Y(n757) );
  NAND2X1 U59 ( .A(n741), .B(n534), .Y(n756) );
  NAND2X1 U60 ( .A(n531), .B(n784), .Y(n740) );
  NAND2X1 U61 ( .A(n698), .B(n654), .Y(n781) );
  INVX1 U62 ( .A(n536), .Y(n876) );
  NAND2BX1 U63 ( .AN(n798), .B(n659), .Y(n726) );
  NAND2X1 U64 ( .A(n807), .B(n699), .Y(n616) );
  NAND2X1 U65 ( .A(n807), .B(n713), .Y(n712) );
  NAND2X1 U66 ( .A(n811), .B(n775), .Y(n826) );
  BUFX3 U67 ( .A(n848), .Y(n534) );
  NAND2X1 U68 ( .A(n659), .B(n780), .Y(n822) );
  INVX1 U69 ( .A(n819), .Y(n854) );
  CLKINVX3 U71 ( .A(n532), .Y(n896) );
  CLKINVX3 U72 ( .A(n811), .Y(n883) );
  NAND2X1 U73 ( .A(n531), .B(n851), .Y(n692) );
  CLKINVX3 U74 ( .A(n814), .Y(n900) );
  NAND2X1 U75 ( .A(n531), .B(n856), .Y(n585) );
  NAND2BX1 U76 ( .AN(n829), .B(n536), .Y(n623) );
  NAND2X1 U77 ( .A(n698), .B(n689), .Y(n818) );
  INVX1 U78 ( .A(n766), .Y(n898) );
  BUFX3 U79 ( .A(a[1]), .Y(n531) );
  NAND2X1 U80 ( .A(a[7]), .B(a[2]), .Y(n828) );
  NAND2X1 U81 ( .A(n532), .B(a[0]), .Y(n814) );
  NAND2X1 U82 ( .A(n863), .B(n539), .Y(n808) );
  INVX1 U83 ( .A(n684), .Y(n906) );
  INVX1 U84 ( .A(n596), .Y(n870) );
  INVX1 U85 ( .A(n634), .Y(n907) );
  NOR2X1 U86 ( .A(n549), .B(n597), .Y(n723) );
  NOR2X1 U87 ( .A(n873), .B(n860), .Y(n675) );
  NOR2BX1 U88 ( .AN(n708), .B(n853), .Y(n834) );
  AOI22X1 U89 ( .A0(n899), .A1(n787), .B0(n897), .B1(n786), .Y(n788) );
  OAI221XL U90 ( .A0(n886), .A1(n549), .B0(n801), .B1(n828), .C0(n782), .Y(
        n787) );
  INVX1 U91 ( .A(n837), .Y(n886) );
  NOR2X1 U92 ( .A(n872), .B(n861), .Y(n636) );
  NAND2X1 U93 ( .A(n700), .B(n539), .Y(n760) );
  NAND2X1 U94 ( .A(n888), .B(n699), .Y(n739) );
  NAND2X1 U95 ( .A(n871), .B(n555), .Y(n684) );
  INVX1 U96 ( .A(n621), .Y(n873) );
  INVX1 U97 ( .A(n689), .Y(n867) );
  INVX1 U98 ( .A(n699), .Y(n863) );
  NOR2X1 U99 ( .A(n865), .B(n867), .Y(n725) );
  INVX1 U100 ( .A(n674), .Y(n885) );
  INVX1 U101 ( .A(n795), .Y(n887) );
  INVX1 U102 ( .A(n715), .Y(n874) );
  INVX1 U104 ( .A(n710), .Y(n881) );
  INVX1 U105 ( .A(n835), .Y(n884) );
  INVX4 U106 ( .A(n535), .Y(n555) );
  NAND2X1 U107 ( .A(n888), .B(n674), .Y(n799) );
  NOR2X1 U108 ( .A(n863), .B(n853), .Y(n824) );
  NOR2X1 U109 ( .A(n860), .B(n867), .Y(n777) );
  INVX1 U110 ( .A(n713), .Y(n877) );
  NAND2X1 U111 ( .A(n859), .B(n534), .Y(n679) );
  NOR2X1 U112 ( .A(n883), .B(n865), .Y(n743) );
  OAI22X1 U113 ( .A0(n620), .A1(n768), .B0(n619), .B1(n812), .Y(n625) );
  AOI211X1 U114 ( .A0(n555), .A1(n820), .B0(n618), .C0(n617), .Y(n619) );
  AOI221X1 U115 ( .A0(n909), .A1(n534), .B0(n895), .B1(n555), .C0(n615), .Y(
        n620) );
  OAI22X1 U116 ( .A0(n858), .A1(n542), .B0(n549), .B1(n616), .Y(n618) );
  NOR2X1 U117 ( .A(n876), .B(n865), .Y(n700) );
  CLKINVX3 U118 ( .A(n809), .Y(n872) );
  OAI22X1 U119 ( .A0(n541), .A1(n715), .B0(n544), .B1(n537), .Y(n680) );
  NAND3X1 U120 ( .A(n537), .B(n809), .C(n539), .Y(n833) );
  NAND2X1 U121 ( .A(n708), .B(n780), .Y(n832) );
  AOI22X1 U122 ( .A0(n898), .A1(n831), .B0(n899), .B1(n830), .Y(n844) );
  OAI221XL U123 ( .A0(n824), .A1(n544), .B0(n892), .B1(n540), .C0(n823), .Y(
        n831) );
  OAI221XL U124 ( .A0(n880), .A1(n544), .B0(n871), .B1(n542), .C0(n827), .Y(
        n830) );
  INVX1 U125 ( .A(n818), .Y(n892) );
  NOR2BX1 U126 ( .AN(n693), .B(n854), .Y(n758) );
  NAND2X1 U127 ( .A(n555), .B(n826), .Y(n735) );
  AOI22X1 U128 ( .A0(n873), .A1(n547), .B0(n555), .B1(n781), .Y(n782) );
  AOI22X1 U129 ( .A0(n899), .A1(n591), .B0(n900), .B1(n590), .Y(n592) );
  OAI221XL U130 ( .A0(n887), .A1(n544), .B0(n878), .B1(n542), .C0(n589), .Y(
        n590) );
  OAI211X1 U131 ( .A0(n596), .A1(n549), .B0(n634), .C0(n588), .Y(n591) );
  AOI22X1 U132 ( .A0(n887), .A1(n555), .B0(n883), .B1(n553), .Y(n589) );
  AOI22X1 U133 ( .A0(n548), .A1(n859), .B0(n675), .B1(n538), .Y(n588) );
  NOR2X1 U134 ( .A(n784), .B(n535), .Y(n825) );
  NAND2X1 U135 ( .A(n679), .B(n780), .Y(n795) );
  NAND2X1 U136 ( .A(n693), .B(n679), .Y(n688) );
  CLKINVX3 U137 ( .A(n784), .Y(n866) );
  INVX1 U138 ( .A(n804), .Y(n852) );
  INVX1 U139 ( .A(n802), .Y(n915) );
  AND2X2 U140 ( .A(n757), .B(n756), .Y(n793) );
  NAND2X1 U141 ( .A(n537), .B(n708), .Y(n796) );
  NAND2X1 U142 ( .A(n784), .B(n820), .Y(n695) );
  INVX1 U143 ( .A(n638), .Y(n910) );
  OAI31XL U144 ( .A0(n720), .A1(n907), .A2(n637), .B0(n897), .Y(n638) );
  OAI21XL U145 ( .A0(n540), .A1(n636), .B0(n635), .Y(n637) );
  INVX1 U146 ( .A(n775), .Y(n875) );
  OAI22X1 U147 ( .A0(n682), .A1(n812), .B0(n681), .B1(n768), .Y(n686) );
  AOI222X1 U148 ( .A0(n861), .A1(n546), .B0(n555), .B1(n678), .C0(n677), .C1(
        n710), .Y(n682) );
  AOI211X1 U149 ( .A0(n555), .A1(n688), .B0(n680), .C0(n723), .Y(n681) );
  NAND2X1 U150 ( .A(n806), .B(n693), .Y(n678) );
  INVX1 U151 ( .A(n585), .Y(n857) );
  CLKINVX8 U152 ( .A(n545), .Y(n544) );
  AOI22X1 U153 ( .A0(n898), .A1(n779), .B0(n900), .B1(n778), .Y(n789) );
  AOI2BB2X1 U154 ( .B0(n538), .B1(n835), .A0N(n544), .A1N(n801), .Y(n773) );
  INVX1 U155 ( .A(n756), .Y(n862) );
  INVX1 U156 ( .A(n623), .Y(n909) );
  NOR2X1 U157 ( .A(n544), .B(n534), .Y(n720) );
  INVX1 U158 ( .A(n694), .Y(n871) );
  AOI221XL U159 ( .A0(n547), .A1(n675), .B0(n710), .B1(n539), .C0(n656), .Y(
        n657) );
  OAI21XL U160 ( .A0(n757), .A1(n549), .B0(n735), .Y(n656) );
  NAND2BX1 U161 ( .AN(n825), .B(n716), .Y(n717) );
  OAI221XL U162 ( .A0(n535), .A1(n726), .B0(n725), .B1(n544), .C0(n724), .Y(
        n727) );
  AOI222X1 U163 ( .A0(n915), .A1(n809), .B0(n723), .B1(n872), .C0(n885), .C1(
        n539), .Y(n724) );
  NOR2X1 U164 ( .A(n853), .B(n854), .Y(n614) );
  OAI221XL U165 ( .A0(n866), .A1(n544), .B0(n890), .B1(n540), .C0(n759), .Y(
        n771) );
  INVX1 U167 ( .A(n755), .Y(n890) );
  AOI22X1 U168 ( .A0(n758), .A1(n555), .B0(n793), .B1(n551), .Y(n759) );
  AOI211X1 U169 ( .A0(n555), .A1(n616), .B0(n587), .C0(n586), .Y(n593) );
  AOI21X1 U170 ( .A0(n621), .A1(n585), .B0(n549), .Y(n586) );
  OAI2BB2X1 U171 ( .B0(n544), .B1(n739), .A0N(n734), .A1N(n539), .Y(n587) );
  AOI2BB2X1 U172 ( .B0(n909), .B1(n534), .A0N(n535), .A1N(n675), .Y(n676) );
  INVX1 U173 ( .A(n712), .Y(n878) );
  OAI221XL U174 ( .A0(n535), .A1(n754), .B0(n758), .B1(n550), .C0(n753), .Y(
        n772) );
  AOI22X1 U175 ( .A0(n547), .A1(n888), .B0(n874), .B1(n538), .Y(n753) );
  AOI211X1 U176 ( .A0(n553), .A1(n826), .B0(n907), .C0(n825), .Y(n827) );
  INVX1 U177 ( .A(n826), .Y(n882) );
  INVX1 U178 ( .A(n774), .Y(n894) );
  CLKINVX3 U179 ( .A(n554), .Y(n550) );
  AOI31X1 U181 ( .A0(n820), .A1(n784), .A2(n555), .B0(n911), .Y(n785) );
  INVX1 U182 ( .A(n833), .Y(n911) );
  INVX1 U183 ( .A(n737), .Y(n903) );
  INVX1 U184 ( .A(n543), .Y(n541) );
  INVX1 U185 ( .A(n797), .Y(n912) );
  AOI221X1 U186 ( .A0(n796), .A1(n551), .B0(n795), .B1(n548), .C0(n794), .Y(
        n797) );
  OAI21XL U187 ( .A0(n535), .A1(n793), .B0(n792), .Y(n794) );
  INVX1 U189 ( .A(n535), .Y(n905) );
  INVX1 U190 ( .A(n539), .Y(n542) );
  AOI22X1 U191 ( .A0(n575), .A1(n896), .B0(n905), .B1(n832), .Y(n579) );
  OAI221XL U192 ( .A0(n864), .A1(n544), .B0(n824), .B1(n828), .C0(n904), .Y(
        n575) );
  INVX1 U193 ( .A(n723), .Y(n904) );
  CLKINVX3 U194 ( .A(n812), .Y(n899) );
  NAND2X1 U195 ( .A(n806), .B(n780), .Y(n837) );
  NAND2X1 U196 ( .A(n537), .B(n756), .Y(n611) );
  AOI22X1 U197 ( .A0(n546), .A1(n611), .B0(n872), .B1(n538), .Y(n572) );
  INVX1 U198 ( .A(n768), .Y(n897) );
  NAND2X1 U199 ( .A(n693), .B(n713), .Y(n662) );
  NOR2X1 U200 ( .A(n858), .B(n798), .Y(n801) );
  INVX1 U201 ( .A(n714), .Y(n893) );
  INVX1 U202 ( .A(n822), .Y(n889) );
  INVX1 U203 ( .A(n616), .Y(n864) );
  INVX1 U204 ( .A(n726), .Y(n891) );
  INVX1 U205 ( .A(n764), .Y(n880) );
  INVX1 U206 ( .A(n781), .Y(n895) );
  NAND2X2 U207 ( .A(n531), .B(n538), .Y(n802) );
  AOI22X1 U208 ( .A0(n574), .A1(n896), .B0(n532), .B1(n573), .Y(n580) );
  OAI221XL U209 ( .A0(n535), .A1(n756), .B0(n636), .B1(n544), .C0(n571), .Y(
        n574) );
  OAI211X1 U210 ( .A0(n834), .A1(n549), .B0(n735), .C0(n572), .Y(n573) );
  AOI2BB2X1 U211 ( .B0(n538), .B1(n726), .A0N(n549), .A1N(n743), .Y(n571) );
  AOI22X1 U212 ( .A0(n532), .A1(n645), .B0(n644), .B1(n896), .Y(n653) );
  OAI222X1 U213 ( .A0(n544), .A1(n781), .B0(n550), .B1(n659), .C0(n893), .C1(
        n541), .Y(n645) );
  OAI221XL U214 ( .A0(n891), .A1(n535), .B0(n550), .B1(n818), .C0(n643), .Y(
        n644) );
  AOI2BB2X1 U215 ( .B0(n834), .B1(n538), .A0N(n544), .A1N(n725), .Y(n643) );
  OAI22X1 U216 ( .A0(n633), .A1(n812), .B0(n632), .B1(n766), .Y(n639) );
  AOI221XL U217 ( .A0(n547), .A1(n739), .B0(n798), .B1(n849), .C0(n631), .Y(
        n632) );
  AOI221XL U218 ( .A0(n866), .A1(n915), .B0(n546), .B1(n712), .C0(n629), .Y(
        n633) );
  OAI32X1 U219 ( .A0(n737), .A1(n859), .A2(n849), .B0(n630), .B1(n903), .Y(
        n631) );
  OAI22X1 U220 ( .A0(n769), .A1(n768), .B0(n767), .B1(n766), .Y(n770) );
  AOI211X1 U221 ( .A0(n880), .A1(n849), .B0(n765), .C0(n906), .Y(n767) );
  AOI221XL U222 ( .A0(n861), .A1(n552), .B0(n546), .B1(n775), .C0(n763), .Y(
        n769) );
  OAI22X1 U223 ( .A0(n541), .A1(n851), .B0(n885), .B1(n549), .Y(n765) );
  NAND2X1 U224 ( .A(n811), .B(n534), .Y(n654) );
  OAI22X1 U225 ( .A0(n815), .A1(n814), .B0(n813), .B1(n812), .Y(n816) );
  AOI221XL U226 ( .A0(n547), .A1(n811), .B0(n875), .B1(n539), .C0(n810), .Y(
        n813) );
  AOI221X1 U227 ( .A0(n555), .A1(n807), .B0(n551), .B1(n806), .C0(n805), .Y(
        n815) );
  OAI221XL U228 ( .A0(n535), .A1(n809), .B0(n878), .B1(n550), .C0(n808), .Y(
        n810) );
  NAND2X1 U229 ( .A(n698), .B(n621), .Y(n774) );
  OAI21XL U230 ( .A0(n601), .A1(n535), .B0(n600), .Y(n604) );
  AOI31X1 U231 ( .A0(n537), .A1(n741), .A2(n599), .B0(n909), .Y(n600) );
  OAI21XL U232 ( .A0(n849), .A1(n621), .B0(n549), .Y(n599) );
  CLKINVX3 U233 ( .A(n741), .Y(n859) );
  NOR2BX1 U234 ( .AN(n659), .B(n861), .Y(n601) );
  AOI22X1 U235 ( .A0(n900), .A1(n842), .B0(n897), .B1(n841), .Y(n843) );
  OAI221XL U236 ( .A0(n856), .A1(n535), .B0(n861), .B1(n550), .C0(n838), .Y(
        n841) );
  OAI221XL U237 ( .A0(n836), .A1(n835), .B0(n834), .B1(n550), .C0(n833), .Y(
        n842) );
  AOI22X1 U238 ( .A0(n546), .A1(n837), .B0(n881), .B1(n538), .Y(n838) );
  NAND2X1 U239 ( .A(n807), .B(n708), .Y(n694) );
  AOI22X1 U240 ( .A0(n555), .A1(n856), .B0(n538), .B1(n775), .Y(n776) );
  OAI221XL U241 ( .A0(n731), .A1(n768), .B0(n730), .B1(n766), .C0(n729), .Y(
        n751) );
  AOI222X1 U242 ( .A0(n547), .A1(n712), .B0(n711), .B1(n710), .C0(n555), .C1(
        n536), .Y(n731) );
  AOI211X1 U243 ( .A0(n877), .A1(n539), .B0(n718), .C0(n717), .Y(n730) );
  AOI22X1 U244 ( .A0(n899), .A1(n728), .B0(n900), .B1(n727), .Y(n729) );
  AOI22X1 U245 ( .A0(n899), .A1(n746), .B0(n898), .B1(n745), .Y(n747) );
  OAI221XL U246 ( .A0(n859), .A1(n544), .B0(n542), .B1(n806), .C0(n744), .Y(
        n745) );
  OAI221XL U247 ( .A0(n884), .A1(n535), .B0(n544), .B1(n739), .C0(n738), .Y(
        n746) );
  AOI21X1 U248 ( .A0(n743), .A1(n551), .B0(n742), .Y(n744) );
  NAND2X1 U249 ( .A(n659), .B(n585), .Y(n755) );
  NAND2X1 U250 ( .A(n698), .B(n804), .Y(n714) );
  OAI21XL U251 ( .A0(n544), .A1(n536), .B0(n802), .Y(n646) );
  NAND2X1 U252 ( .A(n819), .B(n757), .Y(n734) );
  NAND2X1 U253 ( .A(n859), .B(n531), .Y(n754) );
  AOI21X1 U254 ( .A0(n698), .A1(n679), .B0(n544), .Y(n627) );
  OAI21XL U255 ( .A0(n849), .A1(n708), .B0(n549), .Y(n711) );
  OAI21XL U256 ( .A0(n849), .A1(n679), .B0(n549), .Y(n677) );
  AOI21X1 U257 ( .A0(n659), .A1(n740), .B0(n544), .Y(n617) );
  INVX1 U258 ( .A(n531), .Y(n848) );
  OAI21XL U259 ( .A0(n856), .A1(n549), .B0(n663), .Y(n665) );
  NAND2X1 U260 ( .A(n555), .B(n531), .Y(n716) );
  XNOR2X1 U261 ( .A(n902), .B(n531), .Y(n737) );
  NAND2X1 U262 ( .A(n538), .B(n536), .Y(n792) );
  AOI21X1 U263 ( .A0(n832), .A1(n849), .B0(n555), .Y(n836) );
  AOI21X1 U264 ( .A0(n905), .A1(n822), .B0(n821), .Y(n823) );
  AOI21X1 U265 ( .A0(n820), .A1(n819), .B0(n549), .Y(n821) );
  AOI211X1 U266 ( .A0(n883), .A1(n539), .B0(n647), .C0(n646), .Y(n648) );
  OAI222X1 U267 ( .A0(n550), .A1(n806), .B0(n849), .B1(n692), .C0(n544), .C1(
        n820), .Y(n647) );
  XNOR2X1 U268 ( .A(n849), .B(n531), .Y(n761) );
  AOI211X1 U269 ( .A0(n867), .A1(n555), .B0(n651), .C0(n650), .Y(n652) );
  AOI31X1 U270 ( .A0(n808), .A1(n716), .A2(n649), .B0(n532), .Y(n650) );
  OAI22X1 U271 ( .A0(n856), .A1(n802), .B0(n648), .B1(n896), .Y(n651) );
  AOI2BB2X1 U272 ( .B0(n852), .B1(n553), .A0N(n832), .A1N(n544), .Y(n649) );
  NAND2X1 U273 ( .A(n860), .B(n551), .Y(n635) );
  OAI221XL U274 ( .A0(n861), .A1(n550), .B0(n544), .B1(n662), .C0(n661), .Y(
        n668) );
  AOI21X1 U275 ( .A0(n889), .A1(n555), .B0(n660), .Y(n661) );
  AOI21X1 U276 ( .A0(n689), .A1(n757), .B0(n902), .Y(n660) );
  AOI21X1 U277 ( .A0(n872), .A1(n905), .B0(n556), .Y(n557) );
  OAI32X1 U278 ( .A0(n550), .A1(n866), .A2(n869), .B0(n828), .B1(n819), .Y(
        n556) );
  OAI221XL U279 ( .A0(n607), .A1(n766), .B0(n606), .B1(n768), .C0(n605), .Y(
        n608) );
  AOI221XL U280 ( .A0(n555), .A1(n870), .B0(n548), .B1(n799), .C0(n598), .Y(
        n606) );
  AOI22X1 U281 ( .A0(n900), .A1(n604), .B0(n899), .B1(n603), .Y(n605) );
  AOI221X1 U282 ( .A0(n601), .A1(n552), .B0(n539), .B1(n611), .C0(n595), .Y(
        n607) );
  AOI211X1 U283 ( .A0(n721), .A1(n555), .B0(n720), .C0(n719), .Y(n722) );
  AOI21X1 U284 ( .A0(n811), .A1(n537), .B0(n540), .Y(n719) );
  OAI21XL U286 ( .A0(n535), .A1(n804), .B0(n762), .Y(n763) );
  AOI31X1 U287 ( .A0(n811), .A1(n902), .A2(n761), .B0(n914), .Y(n762) );
  INVX1 U288 ( .A(n760), .Y(n914) );
  NOR2BX1 U289 ( .AN(n659), .B(n875), .Y(n721) );
  BUFX3 U290 ( .A(n840), .Y(n535) );
  NAND2X1 U291 ( .A(n849), .B(n902), .Y(n840) );
  OAI222X1 U292 ( .A0(n550), .A1(n715), .B0(n741), .B1(n802), .C0(n544), .C1(
        n714), .Y(n718) );
  OAI222X1 U293 ( .A0(n550), .A1(n755), .B0(n583), .B1(n535), .C0(n544), .C1(
        n888), .Y(n584) );
  AOI21X1 U294 ( .A0(n536), .A1(n534), .B0(n857), .Y(n583) );
  OAI2BB1X1 U295 ( .A0N(n780), .A1N(n548), .B0(n735), .Y(n736) );
  AOI221X1 U296 ( .A0(n876), .A1(n539), .B0(n552), .B1(n734), .C0(n733), .Y(
        n749) );
  AOI21X1 U297 ( .A0(n535), .A1(n732), .B0(n798), .Y(n733) );
  OAI21XL U298 ( .A0(n860), .A1(n852), .B0(n849), .Y(n732) );
  OAI221XL U299 ( .A0(n535), .A1(n713), .B0(n544), .B1(n819), .C0(n634), .Y(
        n595) );
  OAI221XL U300 ( .A0(n531), .A1(n663), .B0(n828), .B1(n708), .C0(n635), .Y(
        n629) );
  OAI221XL U301 ( .A0(n868), .A1(n544), .B0(n889), .B1(n828), .C0(n690), .Y(
        n705) );
  INVX1 U302 ( .A(n688), .Y(n868) );
  AOI32X1 U303 ( .A0(n888), .A1(n741), .A2(n555), .B0(n553), .B1(n689), .Y(
        n690) );
  BUFX3 U304 ( .A(n783), .Y(n537) );
  NAND2X1 U305 ( .A(n531), .B(n536), .Y(n783) );
  AOI211X1 U306 ( .A0(n862), .A1(n539), .B0(n908), .C0(n558), .Y(n559) );
  NOR3X1 U307 ( .A(n544), .B(n883), .C(n861), .Y(n558) );
  INVX1 U308 ( .A(n663), .Y(n908) );
  OAI221XL U309 ( .A0(n855), .A1(n550), .B0(n542), .B1(n537), .C0(n628), .Y(
        n640) );
  INVX1 U310 ( .A(n807), .Y(n855) );
  AOI211X1 U311 ( .A0(n874), .A1(n555), .B0(n913), .C0(n627), .Y(n628) );
  INVX1 U312 ( .A(n808), .Y(n913) );
  AOI211X1 U313 ( .A0(n532), .A1(n568), .B0(n847), .C0(n567), .Y(n569) );
  AOI21X1 U314 ( .A0(n566), .A1(n565), .B0(n532), .Y(n567) );
  OAI221XL U315 ( .A0(n544), .A1(n806), .B0(n601), .B1(n540), .C0(n563), .Y(
        n568) );
  AOI222X1 U316 ( .A0(n866), .A1(n539), .B0(n862), .B1(n553), .C0(n548), .C1(
        n851), .Y(n566) );
  AOI31X1 U317 ( .A0(n702), .A1(n792), .A2(n701), .B0(n814), .Y(n703) );
  OAI2BB1X1 U318 ( .A0N(n699), .A1N(n698), .B0(n552), .Y(n702) );
  AOI22X1 U319 ( .A0(n893), .A1(n905), .B0(n700), .B1(n548), .Y(n701) );
  AOI31X1 U320 ( .A0(n555), .A1(n564), .A2(n883), .B0(n562), .Y(n563) );
  AOI21X1 U321 ( .A0(n807), .A1(n679), .B0(n549), .Y(n562) );
  AOI31X1 U322 ( .A0(n684), .A1(n792), .A2(n683), .B0(n766), .Y(n685) );
  AOI22X1 U323 ( .A0(n865), .A1(n545), .B0(n552), .B1(n809), .Y(n683) );
  AOI31X1 U324 ( .A0(n760), .A1(n623), .A2(n622), .B0(n766), .Y(n624) );
  AOI22X1 U325 ( .A0(n774), .A1(n849), .B0(n893), .B1(n552), .Y(n622) );
  INVX1 U326 ( .A(n839), .Y(n553) );
  INVX1 U327 ( .A(n829), .Y(n545) );
  INVX1 U328 ( .A(n543), .Y(n540) );
  INVX1 U329 ( .A(n828), .Y(n543) );
  INVX1 U330 ( .A(n839), .Y(n554) );
  INVX1 U331 ( .A(n829), .Y(n546) );
  INVX1 U332 ( .A(n829), .Y(n547) );
  INVX1 U333 ( .A(n829), .Y(n548) );
  NAND2X1 U334 ( .A(n807), .B(n654), .Y(n764) );
  AOI21X1 U335 ( .A0(n741), .A1(n740), .B0(n535), .Y(n742) );
  AOI22X1 U336 ( .A0(n538), .A1(n764), .B0(n872), .B1(n902), .Y(n655) );
  XOR2X1 U337 ( .A(n532), .B(n531), .Y(n564) );
  INVX1 U338 ( .A(n839), .Y(n551) );
  INVX1 U339 ( .A(n839), .Y(n552) );
  CLKINVX3 U340 ( .A(n533), .Y(n901) );
  OAI22X1 U341 ( .A0(a[0]), .A1(n670), .B0(n669), .B1(n847), .Y(n671) );
  AOI2BB2X1 U342 ( .B0(n658), .B1(n896), .A0N(n896), .A1N(n657), .Y(n670) );
  AOI22X1 U343 ( .A0(n532), .A1(n668), .B0(n667), .B1(n896), .Y(n669) );
  OAI221XL U344 ( .A0(n876), .A1(n550), .B0(n544), .B1(n806), .C0(n655), .Y(
        n658) );
  CLKINVX3 U345 ( .A(a[3]), .Y(n851) );
  OAI22X1 U346 ( .A0(n697), .A1(n766), .B0(n696), .B1(n768), .Y(n704) );
  AOI221X1 U347 ( .A0(n548), .A1(n692), .B0(n555), .B1(n796), .C0(n691), .Y(
        n697) );
  AOI222X1 U348 ( .A0(n758), .A1(n546), .B0(a[2]), .B1(n695), .C0(n555), .C1(
        n694), .Y(n696) );
  OAI22X1 U349 ( .A0(n887), .A1(n541), .B0(n549), .B1(n536), .Y(n691) );
  OAI22X1 U350 ( .A0(n582), .A1(n901), .B0(n533), .B1(n581), .Y(d[0]) );
  AOI22X1 U351 ( .A0(n580), .A1(a[0]), .B0(n579), .B1(n578), .Y(n581) );
  AOI31X1 U352 ( .A0(n716), .A1(n847), .A2(n570), .B0(n569), .Y(n582) );
  OAI22X1 U353 ( .A0(n533), .A1(n707), .B0(n706), .B1(n901), .Y(d[4]) );
  AOI211X1 U354 ( .A0(n900), .A1(n687), .B0(n686), .C0(n685), .Y(n707) );
  AOI211X1 U355 ( .A0(n899), .A1(n705), .B0(n704), .C0(n703), .Y(n706) );
  OAI22X1 U356 ( .A0(n533), .A1(n642), .B0(n641), .B1(n901), .Y(d[2]) );
  AOI211X1 U357 ( .A0(n900), .A1(n626), .B0(n625), .C0(n624), .Y(n642) );
  AOI211X1 U358 ( .A0(n900), .A1(n640), .B0(n639), .C0(n910), .Y(n641) );
  OAI21XL U359 ( .A0(n846), .A1(n901), .B0(n845), .Y(d[7]) );
  OAI2BB1X1 U360 ( .A0N(n844), .A1N(n843), .B0(n901), .Y(n845) );
  AOI221X1 U361 ( .A0(n898), .A1(n912), .B0(n897), .B1(n817), .C0(n816), .Y(
        n846) );
  INVX1 U362 ( .A(n610), .Y(d[1]) );
  AOI22X1 U363 ( .A0(n533), .A1(n609), .B0(n608), .B1(n901), .Y(n610) );
  OAI221XL U364 ( .A0(n594), .A1(n766), .B0(n593), .B1(n768), .C0(n592), .Y(
        n609) );
  INVX1 U365 ( .A(n673), .Y(d[3]) );
  AOI22X1 U366 ( .A0(n672), .A1(n901), .B0(n533), .B1(n671), .Y(n673) );
  OAI22X1 U367 ( .A0(a[0]), .A1(n653), .B0(n652), .B1(n847), .Y(n672) );
  INVX1 U368 ( .A(n752), .Y(d[5]) );
  AOI22X1 U369 ( .A0(n751), .A1(n901), .B0(n533), .B1(n750), .Y(n752) );
  OAI221XL U370 ( .A0(n749), .A1(n814), .B0(n748), .B1(n768), .C0(n747), .Y(
        n750) );
  AOI22X1 U371 ( .A0(n532), .A1(n561), .B0(n560), .B1(n896), .Y(n570) );
  OAI221XL U372 ( .A0(n879), .A1(n544), .B0(n542), .B1(n888), .C0(n557), .Y(
        n561) );
  INVX1 U373 ( .A(n662), .Y(n879) );
  OAI21XL U374 ( .A0(n533), .A1(n791), .B0(n790), .Y(d[6]) );
  OAI2BB1X1 U375 ( .A0N(n789), .A1N(n788), .B0(n533), .Y(n790) );
  AOI221X1 U376 ( .A0(n899), .A1(n772), .B0(n900), .B1(n771), .C0(n770), .Y(
        n791) );
  NOR2X1 U377 ( .A(n862), .B(n860), .Y(n803) );
  BUFX3 U378 ( .A(n709), .Y(n536) );
  NAND2X1 U379 ( .A(a[4]), .B(n851), .Y(n709) );
  AOI221X1 U380 ( .A0(n915), .A1(n784), .B0(n850), .B1(n665), .C0(n664), .Y(
        n666) );
  NOR3X1 U381 ( .A(n850), .B(a[7]), .C(n859), .Y(n664) );
  INVX1 U382 ( .A(n761), .Y(n850) );
  OAI221XL U383 ( .A0(n535), .A1(n807), .B0(n801), .B1(n544), .C0(n800), .Y(
        n817) );
  AOI22X1 U384 ( .A0(n538), .A1(n799), .B0(n798), .B1(a[2]), .Y(n800) );
  OAI2BB2X1 U385 ( .B0(n613), .B1(n612), .A0N(n743), .A1N(n613), .Y(n626) );
  NOR2X1 U386 ( .A(n547), .B(n553), .Y(n613) );
  AOI22X1 U387 ( .A0(n881), .A1(n849), .B0(a[2]), .B1(n611), .Y(n612) );
  CLKINVX3 U388 ( .A(a[0]), .Y(n847) );
  AOI211X1 U389 ( .A0(n723), .A1(n577), .B0(n576), .C0(a[0]), .Y(n578) );
  NAND2X1 U390 ( .A(n780), .B(n804), .Y(n577) );
  AOI21X1 U391 ( .A0(n802), .A1(n623), .B0(n896), .Y(n576) );
  BUFX3 U392 ( .A(a[5]), .Y(n532) );
  BUFX3 U393 ( .A(a[6]), .Y(n533) );
endmodule


module aes_sbox_2 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915;

  OAI221X4 U28 ( .A0(n882), .A1(n550), .B0(n864), .B1(n544), .C0(n785), .Y(
        n786) );
  OAI221X4 U35 ( .A0(n777), .A1(n544), .B0(n894), .B1(n550), .C0(n776), .Y(
        n778) );
  OAI221X4 U38 ( .A0(n857), .A1(n550), .B0(n891), .B1(n535), .C0(n773), .Y(
        n779) );
  OAI221X4 U70 ( .A0(n876), .A1(n550), .B0(n859), .B1(n544), .C0(n722), .Y(
        n728) );
  OAI221X4 U103 ( .A0(n550), .A1(n835), .B0(n540), .B1(n818), .C0(n676), .Y(
        n687) );
  OAI221X4 U166 ( .A0(n614), .A1(n550), .B0(n544), .B1(n757), .C0(n760), .Y(
        n615) );
  OAI221X4 U180 ( .A0(n550), .A1(n809), .B0(n834), .B1(n544), .C0(n602), .Y(
        n603) );
  OAI32X4 U188 ( .A0(n828), .A1(n859), .A2(n597), .B0(n885), .B1(n550), .Y(
        n598) );
  NAND2X4 U285 ( .A(a[3]), .B(n856), .Y(n741) );
  NAND2X2 U1 ( .A(n856), .B(n851), .Y(n784) );
  INVX1 U2 ( .A(a[7]), .Y(n902) );
  NAND2X1 U3 ( .A(n866), .B(n531), .Y(n693) );
  NAND2X2 U4 ( .A(n536), .B(n741), .Y(n809) );
  OAI221XL U5 ( .A0(n881), .A1(n544), .B0(n542), .B1(n741), .C0(n666), .Y(n667) );
  NAND2X1 U6 ( .A(n531), .B(n741), .Y(n820) );
  NAND2X1 U7 ( .A(n532), .B(n847), .Y(n812) );
  NAND2X2 U8 ( .A(n856), .B(n534), .Y(n806) );
  NAND2X1 U9 ( .A(n883), .B(n531), .Y(n780) );
  OAI222X1 U10 ( .A0(n542), .A1(n804), .B0(n803), .B1(n544), .C0(a[4]), .C1(
        n802), .Y(n805) );
  AOI221XL U11 ( .A0(n915), .A1(n851), .B0(n551), .B1(n809), .C0(n736), .Y(
        n748) );
  AOI211X1 U12 ( .A0(n539), .A1(n851), .B0(n584), .C0(n646), .Y(n594) );
  NAND2X2 U13 ( .A(a[0]), .B(n896), .Y(n766) );
  NAND2X2 U14 ( .A(n847), .B(n896), .Y(n768) );
  OAI221XL U15 ( .A0(a[3]), .A1(n802), .B0(n721), .B1(n550), .C0(n559), .Y(
        n560) );
  NAND2X1 U16 ( .A(a[2]), .B(n902), .Y(n839) );
  NAND2X1 U17 ( .A(a[7]), .B(n849), .Y(n829) );
  CLKINVX3 U18 ( .A(a[2]), .Y(n849) );
  AOI33X1 U19 ( .A0(a[3]), .A1(n539), .A2(n903), .B0(n737), .B1(n741), .B2(
        a[2]), .Y(n738) );
  AOI221X1 U20 ( .A0(n857), .A1(a[2]), .B0(n825), .B1(n564), .C0(n915), .Y(
        n565) );
  AOI21XL U21 ( .A0(n915), .A1(a[4]), .B0(n906), .Y(n602) );
  NAND2X1 U22 ( .A(n531), .B(a[4]), .Y(n698) );
  NAND2X1 U23 ( .A(a[4]), .B(n534), .Y(n659) );
  CLKINVX3 U24 ( .A(a[4]), .Y(n856) );
  AOI22XL U25 ( .A0(n551), .A1(a[3]), .B0(n538), .B1(n856), .Y(n630) );
  NAND2X1 U26 ( .A(a[3]), .B(n534), .Y(n819) );
  NAND2X2 U27 ( .A(n531), .B(a[3]), .Y(n807) );
  NAND2XL U29 ( .A(n905), .B(a[3]), .Y(n663) );
  NAND2X2 U30 ( .A(a[3]), .B(a[4]), .Y(n811) );
  CLKINVX3 U31 ( .A(n541), .Y(n539) );
  NAND2X1 U32 ( .A(n869), .B(n555), .Y(n634) );
  INVX1 U33 ( .A(n597), .Y(n888) );
  NOR2X1 U34 ( .A(n869), .B(n852), .Y(n596) );
  NAND2X1 U36 ( .A(n809), .B(n534), .Y(n708) );
  NOR2X1 U37 ( .A(n534), .B(n883), .Y(n597) );
  CLKINVX3 U39 ( .A(n554), .Y(n549) );
  CLKINVX3 U40 ( .A(n540), .Y(n538) );
  NAND2X1 U41 ( .A(n866), .B(n534), .Y(n689) );
  NAND2X1 U42 ( .A(n876), .B(n534), .Y(n713) );
  NAND2X1 U43 ( .A(n784), .B(n534), .Y(n699) );
  NAND2X1 U44 ( .A(n883), .B(n534), .Y(n674) );
  NAND2X1 U45 ( .A(n537), .B(n654), .Y(n710) );
  NAND2X1 U46 ( .A(n872), .B(n534), .Y(n621) );
  NAND2X1 U47 ( .A(n693), .B(n674), .Y(n835) );
  NAND2X1 U48 ( .A(n775), .B(n708), .Y(n715) );
  INVX1 U49 ( .A(n537), .Y(n869) );
  INVX1 U50 ( .A(n740), .Y(n865) );
  INVX1 U51 ( .A(n806), .Y(n858) );
  INVX1 U52 ( .A(n820), .Y(n861) );
  INVX1 U53 ( .A(n754), .Y(n860) );
  INVX1 U54 ( .A(n692), .Y(n853) );
  NOR2X1 U55 ( .A(n536), .B(n534), .Y(n798) );
  NAND2X1 U56 ( .A(n872), .B(n531), .Y(n775) );
  NAND2X1 U57 ( .A(n534), .B(n851), .Y(n804) );
  NAND2X1 U58 ( .A(n531), .B(n809), .Y(n757) );
  NAND2X1 U59 ( .A(n741), .B(n534), .Y(n756) );
  NAND2X1 U60 ( .A(n531), .B(n784), .Y(n740) );
  NAND2X1 U61 ( .A(n698), .B(n654), .Y(n781) );
  INVX1 U62 ( .A(n536), .Y(n876) );
  NAND2BX1 U63 ( .AN(n798), .B(n659), .Y(n726) );
  NAND2X1 U64 ( .A(n807), .B(n699), .Y(n616) );
  NAND2X1 U65 ( .A(n807), .B(n713), .Y(n712) );
  NAND2X1 U66 ( .A(n811), .B(n775), .Y(n826) );
  BUFX3 U67 ( .A(n848), .Y(n534) );
  NAND2X1 U68 ( .A(n659), .B(n780), .Y(n822) );
  INVX1 U69 ( .A(n819), .Y(n854) );
  CLKINVX3 U71 ( .A(n532), .Y(n896) );
  CLKINVX3 U72 ( .A(n811), .Y(n883) );
  NAND2X1 U73 ( .A(n531), .B(n851), .Y(n692) );
  CLKINVX3 U74 ( .A(n814), .Y(n900) );
  NAND2X1 U75 ( .A(n531), .B(n856), .Y(n585) );
  NAND2BX1 U76 ( .AN(n829), .B(n536), .Y(n623) );
  NAND2X1 U77 ( .A(n698), .B(n689), .Y(n818) );
  INVX1 U78 ( .A(n766), .Y(n898) );
  BUFX3 U79 ( .A(a[1]), .Y(n531) );
  NAND2X1 U80 ( .A(a[7]), .B(a[2]), .Y(n828) );
  NAND2X1 U81 ( .A(n532), .B(a[0]), .Y(n814) );
  NAND2X1 U82 ( .A(n863), .B(n539), .Y(n808) );
  INVX1 U83 ( .A(n684), .Y(n906) );
  INVX1 U84 ( .A(n596), .Y(n870) );
  INVX1 U85 ( .A(n634), .Y(n907) );
  NOR2X1 U86 ( .A(n549), .B(n597), .Y(n723) );
  NOR2X1 U87 ( .A(n873), .B(n860), .Y(n675) );
  NOR2BX1 U88 ( .AN(n708), .B(n853), .Y(n834) );
  AOI22X1 U89 ( .A0(n899), .A1(n787), .B0(n897), .B1(n786), .Y(n788) );
  OAI221XL U90 ( .A0(n886), .A1(n549), .B0(n801), .B1(n828), .C0(n782), .Y(
        n787) );
  INVX1 U91 ( .A(n837), .Y(n886) );
  NOR2X1 U92 ( .A(n872), .B(n861), .Y(n636) );
  NAND2X1 U93 ( .A(n700), .B(n539), .Y(n760) );
  NAND2X1 U94 ( .A(n888), .B(n699), .Y(n739) );
  NAND2X1 U95 ( .A(n871), .B(n555), .Y(n684) );
  INVX1 U96 ( .A(n621), .Y(n873) );
  INVX1 U97 ( .A(n689), .Y(n867) );
  INVX1 U98 ( .A(n699), .Y(n863) );
  NOR2X1 U99 ( .A(n865), .B(n867), .Y(n725) );
  INVX1 U100 ( .A(n674), .Y(n885) );
  INVX1 U101 ( .A(n795), .Y(n887) );
  INVX1 U102 ( .A(n715), .Y(n874) );
  INVX1 U104 ( .A(n710), .Y(n881) );
  INVX1 U105 ( .A(n835), .Y(n884) );
  INVX4 U106 ( .A(n535), .Y(n555) );
  NAND2X1 U107 ( .A(n888), .B(n674), .Y(n799) );
  NOR2X1 U108 ( .A(n863), .B(n853), .Y(n824) );
  NOR2X1 U109 ( .A(n860), .B(n867), .Y(n777) );
  INVX1 U110 ( .A(n713), .Y(n877) );
  NAND2X1 U111 ( .A(n859), .B(n534), .Y(n679) );
  NOR2X1 U112 ( .A(n883), .B(n865), .Y(n743) );
  OAI22X1 U113 ( .A0(n620), .A1(n768), .B0(n619), .B1(n812), .Y(n625) );
  AOI211X1 U114 ( .A0(n555), .A1(n820), .B0(n618), .C0(n617), .Y(n619) );
  AOI221X1 U115 ( .A0(n909), .A1(n534), .B0(n895), .B1(n555), .C0(n615), .Y(
        n620) );
  OAI22X1 U116 ( .A0(n858), .A1(n542), .B0(n549), .B1(n616), .Y(n618) );
  NOR2X1 U117 ( .A(n876), .B(n865), .Y(n700) );
  CLKINVX3 U118 ( .A(n809), .Y(n872) );
  OAI22X1 U119 ( .A0(n541), .A1(n715), .B0(n544), .B1(n537), .Y(n680) );
  NAND3X1 U120 ( .A(n537), .B(n809), .C(n539), .Y(n833) );
  NAND2X1 U121 ( .A(n708), .B(n780), .Y(n832) );
  AOI22X1 U122 ( .A0(n898), .A1(n831), .B0(n899), .B1(n830), .Y(n844) );
  OAI221XL U123 ( .A0(n824), .A1(n544), .B0(n892), .B1(n540), .C0(n823), .Y(
        n831) );
  OAI221XL U124 ( .A0(n880), .A1(n544), .B0(n871), .B1(n542), .C0(n827), .Y(
        n830) );
  INVX1 U125 ( .A(n818), .Y(n892) );
  NOR2BX1 U126 ( .AN(n693), .B(n854), .Y(n758) );
  NAND2X1 U127 ( .A(n555), .B(n826), .Y(n735) );
  AOI22X1 U128 ( .A0(n873), .A1(n547), .B0(n555), .B1(n781), .Y(n782) );
  AOI22X1 U129 ( .A0(n899), .A1(n591), .B0(n900), .B1(n590), .Y(n592) );
  OAI221XL U130 ( .A0(n887), .A1(n544), .B0(n878), .B1(n542), .C0(n589), .Y(
        n590) );
  OAI211X1 U131 ( .A0(n596), .A1(n549), .B0(n634), .C0(n588), .Y(n591) );
  AOI22X1 U132 ( .A0(n887), .A1(n555), .B0(n883), .B1(n553), .Y(n589) );
  AOI22X1 U133 ( .A0(n548), .A1(n859), .B0(n675), .B1(n538), .Y(n588) );
  NOR2X1 U134 ( .A(n784), .B(n535), .Y(n825) );
  NAND2X1 U135 ( .A(n679), .B(n780), .Y(n795) );
  NAND2X1 U136 ( .A(n693), .B(n679), .Y(n688) );
  CLKINVX3 U137 ( .A(n784), .Y(n866) );
  INVX1 U138 ( .A(n804), .Y(n852) );
  INVX1 U139 ( .A(n802), .Y(n915) );
  AND2X2 U140 ( .A(n757), .B(n756), .Y(n793) );
  NAND2X1 U141 ( .A(n537), .B(n708), .Y(n796) );
  NAND2X1 U142 ( .A(n784), .B(n820), .Y(n695) );
  INVX1 U143 ( .A(n638), .Y(n910) );
  OAI31XL U144 ( .A0(n720), .A1(n907), .A2(n637), .B0(n897), .Y(n638) );
  OAI21XL U145 ( .A0(n540), .A1(n636), .B0(n635), .Y(n637) );
  INVX1 U146 ( .A(n775), .Y(n875) );
  OAI22X1 U147 ( .A0(n682), .A1(n812), .B0(n681), .B1(n768), .Y(n686) );
  AOI222X1 U148 ( .A0(n861), .A1(n546), .B0(n555), .B1(n678), .C0(n677), .C1(
        n710), .Y(n682) );
  AOI211X1 U149 ( .A0(n555), .A1(n688), .B0(n680), .C0(n723), .Y(n681) );
  NAND2X1 U150 ( .A(n806), .B(n693), .Y(n678) );
  AOI2BB2X1 U151 ( .B0(n909), .B1(n534), .A0N(n535), .A1N(n675), .Y(n676) );
  INVX1 U152 ( .A(n585), .Y(n857) );
  CLKINVX8 U153 ( .A(n545), .Y(n544) );
  AOI22X1 U154 ( .A0(n898), .A1(n779), .B0(n900), .B1(n778), .Y(n789) );
  AOI2BB2X1 U155 ( .B0(n538), .B1(n835), .A0N(n544), .A1N(n801), .Y(n773) );
  INVX1 U156 ( .A(n756), .Y(n862) );
  INVX1 U157 ( .A(n623), .Y(n909) );
  NOR2X1 U158 ( .A(n544), .B(n534), .Y(n720) );
  INVX1 U159 ( .A(n694), .Y(n871) );
  AOI221XL U160 ( .A0(n547), .A1(n675), .B0(n710), .B1(n539), .C0(n656), .Y(
        n657) );
  OAI21XL U161 ( .A0(n757), .A1(n549), .B0(n735), .Y(n656) );
  NAND2BX1 U162 ( .AN(n825), .B(n716), .Y(n717) );
  OAI221XL U163 ( .A0(n535), .A1(n726), .B0(n725), .B1(n544), .C0(n724), .Y(
        n727) );
  AOI222X1 U164 ( .A0(n915), .A1(n809), .B0(n723), .B1(n872), .C0(n885), .C1(
        n539), .Y(n724) );
  NOR2X1 U165 ( .A(n853), .B(n854), .Y(n614) );
  OAI221XL U167 ( .A0(n866), .A1(n544), .B0(n890), .B1(n540), .C0(n759), .Y(
        n771) );
  INVX1 U168 ( .A(n755), .Y(n890) );
  AOI22X1 U169 ( .A0(n758), .A1(n555), .B0(n793), .B1(n551), .Y(n759) );
  AOI211X1 U170 ( .A0(n555), .A1(n616), .B0(n587), .C0(n586), .Y(n593) );
  AOI21X1 U171 ( .A0(n621), .A1(n585), .B0(n549), .Y(n586) );
  OAI2BB2X1 U172 ( .B0(n544), .B1(n739), .A0N(n734), .A1N(n539), .Y(n587) );
  INVX1 U173 ( .A(n712), .Y(n878) );
  OAI221XL U174 ( .A0(n535), .A1(n754), .B0(n758), .B1(n550), .C0(n753), .Y(
        n772) );
  AOI22X1 U175 ( .A0(n547), .A1(n888), .B0(n874), .B1(n538), .Y(n753) );
  AOI211X1 U176 ( .A0(n553), .A1(n826), .B0(n907), .C0(n825), .Y(n827) );
  INVX1 U177 ( .A(n826), .Y(n882) );
  INVX1 U178 ( .A(n774), .Y(n894) );
  CLKINVX3 U179 ( .A(n554), .Y(n550) );
  AOI31X1 U181 ( .A0(n820), .A1(n784), .A2(n555), .B0(n911), .Y(n785) );
  INVX1 U182 ( .A(n833), .Y(n911) );
  INVX1 U183 ( .A(n737), .Y(n903) );
  INVX1 U184 ( .A(n543), .Y(n541) );
  INVX1 U185 ( .A(n797), .Y(n912) );
  AOI221X1 U186 ( .A0(n796), .A1(n551), .B0(n795), .B1(n548), .C0(n794), .Y(
        n797) );
  OAI21XL U187 ( .A0(n535), .A1(n793), .B0(n792), .Y(n794) );
  INVX1 U189 ( .A(n535), .Y(n905) );
  INVX1 U190 ( .A(n539), .Y(n542) );
  AOI22X1 U191 ( .A0(n575), .A1(n896), .B0(n905), .B1(n832), .Y(n579) );
  OAI221XL U192 ( .A0(n864), .A1(n544), .B0(n824), .B1(n828), .C0(n904), .Y(
        n575) );
  INVX1 U193 ( .A(n723), .Y(n904) );
  CLKINVX3 U194 ( .A(n812), .Y(n899) );
  NAND2X1 U195 ( .A(n806), .B(n780), .Y(n837) );
  NAND2X1 U196 ( .A(n537), .B(n756), .Y(n611) );
  AOI22X1 U197 ( .A0(n546), .A1(n611), .B0(n872), .B1(n538), .Y(n572) );
  INVX1 U198 ( .A(n768), .Y(n897) );
  NAND2X1 U199 ( .A(n693), .B(n713), .Y(n662) );
  NOR2X1 U200 ( .A(n858), .B(n798), .Y(n801) );
  INVX1 U201 ( .A(n714), .Y(n893) );
  INVX1 U202 ( .A(n822), .Y(n889) );
  INVX1 U203 ( .A(n616), .Y(n864) );
  INVX1 U204 ( .A(n726), .Y(n891) );
  INVX1 U205 ( .A(n764), .Y(n880) );
  INVX1 U206 ( .A(n781), .Y(n895) );
  NAND2X2 U207 ( .A(n531), .B(n538), .Y(n802) );
  AOI22X1 U208 ( .A0(n574), .A1(n896), .B0(n532), .B1(n573), .Y(n580) );
  OAI221XL U209 ( .A0(n535), .A1(n756), .B0(n636), .B1(n544), .C0(n571), .Y(
        n574) );
  OAI211X1 U210 ( .A0(n834), .A1(n549), .B0(n735), .C0(n572), .Y(n573) );
  AOI2BB2X1 U211 ( .B0(n538), .B1(n726), .A0N(n549), .A1N(n743), .Y(n571) );
  AOI22X1 U212 ( .A0(n532), .A1(n645), .B0(n644), .B1(n896), .Y(n653) );
  OAI222X1 U213 ( .A0(n544), .A1(n781), .B0(n550), .B1(n659), .C0(n893), .C1(
        n541), .Y(n645) );
  OAI221XL U214 ( .A0(n891), .A1(n535), .B0(n550), .B1(n818), .C0(n643), .Y(
        n644) );
  AOI2BB2X1 U215 ( .B0(n834), .B1(n538), .A0N(n544), .A1N(n725), .Y(n643) );
  OAI22X1 U216 ( .A0(n633), .A1(n812), .B0(n632), .B1(n766), .Y(n639) );
  AOI221XL U217 ( .A0(n547), .A1(n739), .B0(n798), .B1(n849), .C0(n631), .Y(
        n632) );
  AOI221XL U218 ( .A0(n866), .A1(n915), .B0(n546), .B1(n712), .C0(n629), .Y(
        n633) );
  OAI32X1 U219 ( .A0(n737), .A1(n859), .A2(n849), .B0(n630), .B1(n903), .Y(
        n631) );
  OAI22X1 U220 ( .A0(n769), .A1(n768), .B0(n767), .B1(n766), .Y(n770) );
  AOI211X1 U221 ( .A0(n880), .A1(n849), .B0(n765), .C0(n906), .Y(n767) );
  AOI221XL U222 ( .A0(n861), .A1(n552), .B0(n546), .B1(n775), .C0(n763), .Y(
        n769) );
  OAI22X1 U223 ( .A0(n541), .A1(n851), .B0(n885), .B1(n549), .Y(n765) );
  NAND2X1 U224 ( .A(n811), .B(n534), .Y(n654) );
  OAI22X1 U225 ( .A0(n815), .A1(n814), .B0(n813), .B1(n812), .Y(n816) );
  AOI221XL U226 ( .A0(n547), .A1(n811), .B0(n875), .B1(n539), .C0(n810), .Y(
        n813) );
  AOI221X1 U227 ( .A0(n555), .A1(n807), .B0(n551), .B1(n806), .C0(n805), .Y(
        n815) );
  OAI221XL U228 ( .A0(n535), .A1(n809), .B0(n878), .B1(n550), .C0(n808), .Y(
        n810) );
  NAND2X1 U229 ( .A(n698), .B(n621), .Y(n774) );
  OAI21XL U230 ( .A0(n601), .A1(n535), .B0(n600), .Y(n604) );
  AOI31X1 U231 ( .A0(n537), .A1(n741), .A2(n599), .B0(n909), .Y(n600) );
  OAI21XL U232 ( .A0(n849), .A1(n621), .B0(n549), .Y(n599) );
  CLKINVX3 U233 ( .A(n741), .Y(n859) );
  NOR2BX1 U234 ( .AN(n659), .B(n861), .Y(n601) );
  AOI22X1 U235 ( .A0(n900), .A1(n842), .B0(n897), .B1(n841), .Y(n843) );
  OAI221XL U236 ( .A0(n856), .A1(n535), .B0(n861), .B1(n550), .C0(n838), .Y(
        n841) );
  OAI221XL U237 ( .A0(n836), .A1(n835), .B0(n834), .B1(n550), .C0(n833), .Y(
        n842) );
  AOI22X1 U238 ( .A0(n546), .A1(n837), .B0(n881), .B1(n538), .Y(n838) );
  NAND2X1 U239 ( .A(n807), .B(n708), .Y(n694) );
  AOI22X1 U240 ( .A0(n555), .A1(n856), .B0(n538), .B1(n775), .Y(n776) );
  OAI221XL U241 ( .A0(n731), .A1(n768), .B0(n730), .B1(n766), .C0(n729), .Y(
        n751) );
  AOI222X1 U242 ( .A0(n547), .A1(n712), .B0(n711), .B1(n710), .C0(n555), .C1(
        n536), .Y(n731) );
  AOI211X1 U243 ( .A0(n877), .A1(n539), .B0(n718), .C0(n717), .Y(n730) );
  AOI22X1 U244 ( .A0(n899), .A1(n728), .B0(n900), .B1(n727), .Y(n729) );
  AOI22X1 U245 ( .A0(n899), .A1(n746), .B0(n898), .B1(n745), .Y(n747) );
  OAI221XL U246 ( .A0(n859), .A1(n544), .B0(n542), .B1(n806), .C0(n744), .Y(
        n745) );
  OAI221XL U247 ( .A0(n884), .A1(n535), .B0(n544), .B1(n739), .C0(n738), .Y(
        n746) );
  AOI21X1 U248 ( .A0(n743), .A1(n551), .B0(n742), .Y(n744) );
  NAND2X1 U249 ( .A(n659), .B(n585), .Y(n755) );
  NAND2X1 U250 ( .A(n698), .B(n804), .Y(n714) );
  OAI21XL U251 ( .A0(n544), .A1(n536), .B0(n802), .Y(n646) );
  NAND2X1 U252 ( .A(n819), .B(n757), .Y(n734) );
  NAND2X1 U253 ( .A(n859), .B(n531), .Y(n754) );
  AOI21X1 U254 ( .A0(n698), .A1(n679), .B0(n544), .Y(n627) );
  OAI21XL U255 ( .A0(n849), .A1(n708), .B0(n549), .Y(n711) );
  OAI21XL U256 ( .A0(n849), .A1(n679), .B0(n549), .Y(n677) );
  AOI21X1 U257 ( .A0(n659), .A1(n740), .B0(n544), .Y(n617) );
  INVX1 U258 ( .A(n531), .Y(n848) );
  OAI21XL U259 ( .A0(n856), .A1(n549), .B0(n663), .Y(n665) );
  NAND2X1 U260 ( .A(n555), .B(n531), .Y(n716) );
  XNOR2X1 U261 ( .A(n902), .B(n531), .Y(n737) );
  NAND2X1 U262 ( .A(n538), .B(n536), .Y(n792) );
  AOI21X1 U263 ( .A0(n832), .A1(n849), .B0(n555), .Y(n836) );
  AOI21X1 U264 ( .A0(n905), .A1(n822), .B0(n821), .Y(n823) );
  AOI21X1 U265 ( .A0(n820), .A1(n819), .B0(n549), .Y(n821) );
  AOI211X1 U266 ( .A0(n883), .A1(n539), .B0(n647), .C0(n646), .Y(n648) );
  OAI222X1 U267 ( .A0(n550), .A1(n806), .B0(n849), .B1(n692), .C0(n544), .C1(
        n820), .Y(n647) );
  XNOR2X1 U268 ( .A(n849), .B(n531), .Y(n761) );
  AOI211X1 U269 ( .A0(n867), .A1(n555), .B0(n651), .C0(n650), .Y(n652) );
  AOI31X1 U270 ( .A0(n808), .A1(n716), .A2(n649), .B0(n532), .Y(n650) );
  OAI22X1 U271 ( .A0(n856), .A1(n802), .B0(n648), .B1(n896), .Y(n651) );
  AOI2BB2X1 U272 ( .B0(n852), .B1(n553), .A0N(n832), .A1N(n544), .Y(n649) );
  NAND2X1 U273 ( .A(n860), .B(n551), .Y(n635) );
  OAI221XL U274 ( .A0(n861), .A1(n550), .B0(n544), .B1(n662), .C0(n661), .Y(
        n668) );
  AOI21X1 U275 ( .A0(n889), .A1(n555), .B0(n660), .Y(n661) );
  AOI21X1 U276 ( .A0(n689), .A1(n757), .B0(n902), .Y(n660) );
  AOI21X1 U277 ( .A0(n872), .A1(n905), .B0(n556), .Y(n557) );
  OAI32X1 U278 ( .A0(n550), .A1(n866), .A2(n869), .B0(n828), .B1(n819), .Y(
        n556) );
  OAI221XL U279 ( .A0(n607), .A1(n766), .B0(n606), .B1(n768), .C0(n605), .Y(
        n608) );
  AOI221XL U280 ( .A0(n555), .A1(n870), .B0(n548), .B1(n799), .C0(n598), .Y(
        n606) );
  AOI22X1 U281 ( .A0(n900), .A1(n604), .B0(n899), .B1(n603), .Y(n605) );
  AOI221X1 U282 ( .A0(n601), .A1(n552), .B0(n539), .B1(n611), .C0(n595), .Y(
        n607) );
  AOI211X1 U283 ( .A0(n721), .A1(n555), .B0(n720), .C0(n719), .Y(n722) );
  AOI21X1 U284 ( .A0(n811), .A1(n537), .B0(n540), .Y(n719) );
  OAI21XL U286 ( .A0(n535), .A1(n804), .B0(n762), .Y(n763) );
  AOI31X1 U287 ( .A0(n811), .A1(n902), .A2(n761), .B0(n914), .Y(n762) );
  INVX1 U288 ( .A(n760), .Y(n914) );
  NOR2BX1 U289 ( .AN(n659), .B(n875), .Y(n721) );
  BUFX3 U290 ( .A(n840), .Y(n535) );
  NAND2X1 U291 ( .A(n849), .B(n902), .Y(n840) );
  OAI222X1 U292 ( .A0(n550), .A1(n715), .B0(n741), .B1(n802), .C0(n544), .C1(
        n714), .Y(n718) );
  OAI222X1 U293 ( .A0(n550), .A1(n755), .B0(n583), .B1(n535), .C0(n544), .C1(
        n888), .Y(n584) );
  AOI21X1 U294 ( .A0(n536), .A1(n534), .B0(n857), .Y(n583) );
  OAI2BB1X1 U295 ( .A0N(n780), .A1N(n548), .B0(n735), .Y(n736) );
  AOI221X1 U296 ( .A0(n876), .A1(n539), .B0(n552), .B1(n734), .C0(n733), .Y(
        n749) );
  AOI21X1 U297 ( .A0(n535), .A1(n732), .B0(n798), .Y(n733) );
  OAI21XL U298 ( .A0(n860), .A1(n852), .B0(n849), .Y(n732) );
  OAI221XL U299 ( .A0(n535), .A1(n713), .B0(n544), .B1(n819), .C0(n634), .Y(
        n595) );
  OAI221XL U300 ( .A0(n531), .A1(n663), .B0(n828), .B1(n708), .C0(n635), .Y(
        n629) );
  OAI221XL U301 ( .A0(n868), .A1(n544), .B0(n889), .B1(n828), .C0(n690), .Y(
        n705) );
  INVX1 U302 ( .A(n688), .Y(n868) );
  AOI32X1 U303 ( .A0(n888), .A1(n741), .A2(n555), .B0(n553), .B1(n689), .Y(
        n690) );
  BUFX3 U304 ( .A(n783), .Y(n537) );
  NAND2X1 U305 ( .A(n531), .B(n536), .Y(n783) );
  AOI211X1 U306 ( .A0(n862), .A1(n539), .B0(n908), .C0(n558), .Y(n559) );
  NOR3X1 U307 ( .A(n544), .B(n883), .C(n861), .Y(n558) );
  INVX1 U308 ( .A(n663), .Y(n908) );
  OAI221XL U309 ( .A0(n855), .A1(n550), .B0(n542), .B1(n537), .C0(n628), .Y(
        n640) );
  INVX1 U310 ( .A(n807), .Y(n855) );
  AOI211X1 U311 ( .A0(n874), .A1(n555), .B0(n913), .C0(n627), .Y(n628) );
  INVX1 U312 ( .A(n808), .Y(n913) );
  AOI211X1 U313 ( .A0(n532), .A1(n568), .B0(n847), .C0(n567), .Y(n569) );
  AOI21X1 U314 ( .A0(n566), .A1(n565), .B0(n532), .Y(n567) );
  OAI221XL U315 ( .A0(n544), .A1(n806), .B0(n601), .B1(n540), .C0(n563), .Y(
        n568) );
  AOI222X1 U316 ( .A0(n866), .A1(n539), .B0(n862), .B1(n553), .C0(n548), .C1(
        n851), .Y(n566) );
  AOI31X1 U317 ( .A0(n702), .A1(n792), .A2(n701), .B0(n814), .Y(n703) );
  OAI2BB1X1 U318 ( .A0N(n699), .A1N(n698), .B0(n552), .Y(n702) );
  AOI22X1 U319 ( .A0(n893), .A1(n905), .B0(n700), .B1(n548), .Y(n701) );
  AOI31X1 U320 ( .A0(n555), .A1(n564), .A2(n883), .B0(n562), .Y(n563) );
  AOI21X1 U321 ( .A0(n807), .A1(n679), .B0(n549), .Y(n562) );
  AOI31X1 U322 ( .A0(n684), .A1(n792), .A2(n683), .B0(n766), .Y(n685) );
  AOI22X1 U323 ( .A0(n865), .A1(n545), .B0(n552), .B1(n809), .Y(n683) );
  AOI31X1 U324 ( .A0(n760), .A1(n623), .A2(n622), .B0(n766), .Y(n624) );
  AOI22X1 U325 ( .A0(n774), .A1(n849), .B0(n893), .B1(n552), .Y(n622) );
  INVX1 U326 ( .A(n839), .Y(n553) );
  INVX1 U327 ( .A(n829), .Y(n545) );
  INVX1 U328 ( .A(n543), .Y(n540) );
  INVX1 U329 ( .A(n828), .Y(n543) );
  INVX1 U330 ( .A(n839), .Y(n554) );
  INVX1 U331 ( .A(n829), .Y(n546) );
  INVX1 U332 ( .A(n829), .Y(n547) );
  INVX1 U333 ( .A(n829), .Y(n548) );
  NAND2X1 U334 ( .A(n807), .B(n654), .Y(n764) );
  AOI21X1 U335 ( .A0(n741), .A1(n740), .B0(n535), .Y(n742) );
  AOI22X1 U336 ( .A0(n538), .A1(n764), .B0(n872), .B1(n902), .Y(n655) );
  XOR2X1 U337 ( .A(n532), .B(n531), .Y(n564) );
  INVX1 U338 ( .A(n839), .Y(n551) );
  INVX1 U339 ( .A(n839), .Y(n552) );
  CLKINVX3 U340 ( .A(n533), .Y(n901) );
  OAI22X1 U341 ( .A0(a[0]), .A1(n670), .B0(n669), .B1(n847), .Y(n671) );
  AOI2BB2X1 U342 ( .B0(n658), .B1(n896), .A0N(n896), .A1N(n657), .Y(n670) );
  AOI22X1 U343 ( .A0(n532), .A1(n668), .B0(n667), .B1(n896), .Y(n669) );
  OAI221XL U344 ( .A0(n876), .A1(n550), .B0(n544), .B1(n806), .C0(n655), .Y(
        n658) );
  CLKINVX3 U345 ( .A(a[3]), .Y(n851) );
  OAI22X1 U346 ( .A0(n697), .A1(n766), .B0(n696), .B1(n768), .Y(n704) );
  AOI221X1 U347 ( .A0(n548), .A1(n692), .B0(n555), .B1(n796), .C0(n691), .Y(
        n697) );
  AOI222X1 U348 ( .A0(n758), .A1(n546), .B0(a[2]), .B1(n695), .C0(n555), .C1(
        n694), .Y(n696) );
  OAI22X1 U349 ( .A0(n887), .A1(n541), .B0(n549), .B1(n536), .Y(n691) );
  OAI22X1 U350 ( .A0(n582), .A1(n901), .B0(n533), .B1(n581), .Y(d[0]) );
  AOI22X1 U351 ( .A0(n580), .A1(a[0]), .B0(n579), .B1(n578), .Y(n581) );
  AOI31X1 U352 ( .A0(n716), .A1(n847), .A2(n570), .B0(n569), .Y(n582) );
  OAI22X1 U353 ( .A0(n533), .A1(n707), .B0(n706), .B1(n901), .Y(d[4]) );
  AOI211X1 U354 ( .A0(n900), .A1(n687), .B0(n686), .C0(n685), .Y(n707) );
  AOI211X1 U355 ( .A0(n899), .A1(n705), .B0(n704), .C0(n703), .Y(n706) );
  OAI22X1 U356 ( .A0(n533), .A1(n642), .B0(n641), .B1(n901), .Y(d[2]) );
  AOI211X1 U357 ( .A0(n900), .A1(n626), .B0(n625), .C0(n624), .Y(n642) );
  AOI211X1 U358 ( .A0(n900), .A1(n640), .B0(n639), .C0(n910), .Y(n641) );
  OAI21XL U359 ( .A0(n846), .A1(n901), .B0(n845), .Y(d[7]) );
  OAI2BB1X1 U360 ( .A0N(n844), .A1N(n843), .B0(n901), .Y(n845) );
  AOI221X1 U361 ( .A0(n898), .A1(n912), .B0(n897), .B1(n817), .C0(n816), .Y(
        n846) );
  INVX1 U362 ( .A(n610), .Y(d[1]) );
  AOI22X1 U363 ( .A0(n533), .A1(n609), .B0(n608), .B1(n901), .Y(n610) );
  OAI221XL U364 ( .A0(n594), .A1(n766), .B0(n593), .B1(n768), .C0(n592), .Y(
        n609) );
  INVX1 U365 ( .A(n673), .Y(d[3]) );
  AOI22X1 U366 ( .A0(n672), .A1(n901), .B0(n533), .B1(n671), .Y(n673) );
  OAI22X1 U367 ( .A0(a[0]), .A1(n653), .B0(n652), .B1(n847), .Y(n672) );
  INVX1 U368 ( .A(n752), .Y(d[5]) );
  AOI22X1 U369 ( .A0(n751), .A1(n901), .B0(n533), .B1(n750), .Y(n752) );
  OAI221XL U370 ( .A0(n749), .A1(n814), .B0(n748), .B1(n768), .C0(n747), .Y(
        n750) );
  AOI22X1 U371 ( .A0(n532), .A1(n561), .B0(n560), .B1(n896), .Y(n570) );
  OAI221XL U372 ( .A0(n879), .A1(n544), .B0(n542), .B1(n888), .C0(n557), .Y(
        n561) );
  INVX1 U373 ( .A(n662), .Y(n879) );
  OAI21XL U374 ( .A0(n533), .A1(n791), .B0(n790), .Y(d[6]) );
  OAI2BB1X1 U375 ( .A0N(n789), .A1N(n788), .B0(n533), .Y(n790) );
  AOI221X1 U376 ( .A0(n899), .A1(n772), .B0(n900), .B1(n771), .C0(n770), .Y(
        n791) );
  NOR2X1 U377 ( .A(n862), .B(n860), .Y(n803) );
  BUFX3 U378 ( .A(n709), .Y(n536) );
  NAND2X1 U379 ( .A(a[4]), .B(n851), .Y(n709) );
  AOI221X1 U380 ( .A0(n915), .A1(n784), .B0(n850), .B1(n665), .C0(n664), .Y(
        n666) );
  NOR3X1 U381 ( .A(n850), .B(a[7]), .C(n859), .Y(n664) );
  INVX1 U382 ( .A(n761), .Y(n850) );
  OAI221XL U383 ( .A0(n535), .A1(n807), .B0(n801), .B1(n544), .C0(n800), .Y(
        n817) );
  AOI22X1 U384 ( .A0(n538), .A1(n799), .B0(n798), .B1(a[2]), .Y(n800) );
  OAI2BB2X1 U385 ( .B0(n613), .B1(n612), .A0N(n743), .A1N(n613), .Y(n626) );
  NOR2X1 U386 ( .A(n547), .B(n553), .Y(n613) );
  AOI22X1 U387 ( .A0(n881), .A1(n849), .B0(a[2]), .B1(n611), .Y(n612) );
  CLKINVX3 U388 ( .A(a[0]), .Y(n847) );
  AOI211X1 U389 ( .A0(n723), .A1(n577), .B0(n576), .C0(a[0]), .Y(n578) );
  NAND2X1 U390 ( .A(n780), .B(n804), .Y(n577) );
  AOI21X1 U391 ( .A0(n802), .A1(n623), .B0(n896), .Y(n576) );
  BUFX3 U392 ( .A(a[5]), .Y(n532) );
  BUFX3 U393 ( .A(a[6]), .Y(n533) );
endmodule


module aes_key_expand_128 ( clk, kld, key, wo_0, wo_1, wo_2, wo_3 );
  input [127:0] key;
  output [31:0] wo_0;
  output [31:0] wo_1;
  output [31:0] wo_2;
  output [31:0] wo_3;
  input clk, kld;
  wire   N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, n258, n259, n260, n261, n262,
         n263, n264, n265, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474;
  wire   [31:0] subword;
  wire   [31:0] rcon;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23;

  aes_sbox_4 u0 ( .a(wo_3[23:16]), .d(subword[31:24]) );
  aes_sbox_3 u1 ( .a(wo_3[15:8]), .d(subword[23:16]) );
  aes_sbox_2 u2 ( .a(wo_3[7:0]), .d(subword[15:8]) );
  aes_sbox_1 u3 ( .a(wo_3[31:24]), .d(subword[7:0]) );
  aes_rcon r0 ( .clk(clk), .kld(n370), .out({rcon[31:24], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23}) );
  DFFHQX1 \w_reg[2][8]  ( .D(n67), .CK(clk), .Q(wo_2[8]) );
  DFFHQX1 \w_reg[1][8]  ( .D(n66), .CK(clk), .Q(wo_1[8]) );
  DFFHQX1 \w_reg[0][8]  ( .D(n65), .CK(clk), .Q(wo_0[8]) );
  DFFHQX1 \w_reg[2][9]  ( .D(n71), .CK(clk), .Q(wo_2[9]) );
  DFFHQX1 \w_reg[1][9]  ( .D(n70), .CK(clk), .Q(wo_1[9]) );
  DFFHQX1 \w_reg[0][9]  ( .D(n69), .CK(clk), .Q(wo_0[9]) );
  DFFHQX1 \w_reg[2][10]  ( .D(n75), .CK(clk), .Q(wo_2[10]) );
  DFFHQX1 \w_reg[1][10]  ( .D(n74), .CK(clk), .Q(wo_1[10]) );
  DFFHQX1 \w_reg[0][10]  ( .D(n73), .CK(clk), .Q(wo_0[10]) );
  DFFHQX1 \w_reg[2][11]  ( .D(n79), .CK(clk), .Q(wo_2[11]) );
  DFFHQX1 \w_reg[1][11]  ( .D(n78), .CK(clk), .Q(wo_1[11]) );
  DFFHQX1 \w_reg[0][11]  ( .D(n77), .CK(clk), .Q(wo_0[11]) );
  DFFHQX1 \w_reg[2][12]  ( .D(n83), .CK(clk), .Q(wo_2[12]) );
  DFFHQX1 \w_reg[1][12]  ( .D(n82), .CK(clk), .Q(wo_1[12]) );
  DFFHQX1 \w_reg[0][12]  ( .D(n81), .CK(clk), .Q(wo_0[12]) );
  DFFHQX1 \w_reg[2][13]  ( .D(n87), .CK(clk), .Q(wo_2[13]) );
  DFFHQX1 \w_reg[1][13]  ( .D(n86), .CK(clk), .Q(wo_1[13]) );
  DFFHQX1 \w_reg[0][13]  ( .D(n85), .CK(clk), .Q(wo_0[13]) );
  DFFHQX1 \w_reg[2][14]  ( .D(n91), .CK(clk), .Q(wo_2[14]) );
  DFFHQX1 \w_reg[1][14]  ( .D(n90), .CK(clk), .Q(wo_1[14]) );
  DFFHQX1 \w_reg[0][14]  ( .D(n89), .CK(clk), .Q(wo_0[14]) );
  DFFHQX1 \w_reg[2][16]  ( .D(n35), .CK(clk), .Q(wo_2[16]) );
  DFFHQX1 \w_reg[1][16]  ( .D(n34), .CK(clk), .Q(wo_1[16]) );
  DFFHQX1 \w_reg[0][16]  ( .D(n33), .CK(clk), .Q(wo_0[16]) );
  DFFHQX1 \w_reg[2][17]  ( .D(n39), .CK(clk), .Q(wo_2[17]) );
  DFFHQX1 \w_reg[1][17]  ( .D(n38), .CK(clk), .Q(wo_1[17]) );
  DFFHQX1 \w_reg[0][17]  ( .D(n37), .CK(clk), .Q(wo_0[17]) );
  DFFHQX1 \w_reg[2][18]  ( .D(n43), .CK(clk), .Q(wo_2[18]) );
  DFFHQX1 \w_reg[1][18]  ( .D(n42), .CK(clk), .Q(wo_1[18]) );
  DFFHQX1 \w_reg[0][18]  ( .D(n41), .CK(clk), .Q(wo_0[18]) );
  DFFHQX1 \w_reg[2][19]  ( .D(n47), .CK(clk), .Q(wo_2[19]) );
  DFFHQX1 \w_reg[1][19]  ( .D(n46), .CK(clk), .Q(wo_1[19]) );
  DFFHQX1 \w_reg[0][19]  ( .D(n45), .CK(clk), .Q(wo_0[19]) );
  DFFHQX1 \w_reg[2][20]  ( .D(n51), .CK(clk), .Q(wo_2[20]) );
  DFFHQX1 \w_reg[1][20]  ( .D(n50), .CK(clk), .Q(wo_1[20]) );
  DFFHQX1 \w_reg[0][20]  ( .D(n49), .CK(clk), .Q(wo_0[20]) );
  DFFHQX1 \w_reg[2][21]  ( .D(n55), .CK(clk), .Q(wo_2[21]) );
  DFFHQX1 \w_reg[1][21]  ( .D(n54), .CK(clk), .Q(wo_1[21]) );
  DFFHQX1 \w_reg[0][21]  ( .D(n53), .CK(clk), .Q(wo_0[21]) );
  DFFHQX1 \w_reg[2][22]  ( .D(n59), .CK(clk), .Q(wo_2[22]) );
  DFFHQX1 \w_reg[1][22]  ( .D(n58), .CK(clk), .Q(wo_1[22]) );
  DFFHQX1 \w_reg[0][22]  ( .D(n57), .CK(clk), .Q(wo_0[22]) );
  DFFHQX1 \w_reg[2][24]  ( .D(n3), .CK(clk), .Q(wo_2[24]) );
  DFFHQX1 \w_reg[1][24]  ( .D(n2), .CK(clk), .Q(wo_1[24]) );
  DFFHQX1 \w_reg[2][25]  ( .D(n7), .CK(clk), .Q(wo_2[25]) );
  DFFHQX1 \w_reg[1][25]  ( .D(n6), .CK(clk), .Q(wo_1[25]) );
  DFFHQX1 \w_reg[2][26]  ( .D(n11), .CK(clk), .Q(wo_2[26]) );
  DFFHQX1 \w_reg[1][26]  ( .D(n10), .CK(clk), .Q(wo_1[26]) );
  DFFHQX1 \w_reg[2][27]  ( .D(n15), .CK(clk), .Q(wo_2[27]) );
  DFFHQX1 \w_reg[1][27]  ( .D(n14), .CK(clk), .Q(wo_1[27]) );
  DFFHQX1 \w_reg[2][28]  ( .D(n19), .CK(clk), .Q(wo_2[28]) );
  DFFHQX1 \w_reg[1][28]  ( .D(n18), .CK(clk), .Q(wo_1[28]) );
  DFFHQX1 \w_reg[2][29]  ( .D(n23), .CK(clk), .Q(wo_2[29]) );
  DFFHQX1 \w_reg[1][29]  ( .D(n22), .CK(clk), .Q(wo_1[29]) );
  DFFHQX1 \w_reg[2][30]  ( .D(n27), .CK(clk), .Q(wo_2[30]) );
  DFFHQX1 \w_reg[1][30]  ( .D(n26), .CK(clk), .Q(wo_1[30]) );
  DFFHQX1 \w_reg[2][0]  ( .D(n99), .CK(clk), .Q(wo_2[0]) );
  DFFHQX1 \w_reg[1][0]  ( .D(n98), .CK(clk), .Q(wo_1[0]) );
  DFFHQX1 \w_reg[0][0]  ( .D(n97), .CK(clk), .Q(wo_0[0]) );
  DFFHQX1 \w_reg[2][1]  ( .D(n103), .CK(clk), .Q(wo_2[1]) );
  DFFHQX1 \w_reg[1][1]  ( .D(n102), .CK(clk), .Q(wo_1[1]) );
  DFFHQX1 \w_reg[0][1]  ( .D(n101), .CK(clk), .Q(wo_0[1]) );
  DFFHQX1 \w_reg[2][2]  ( .D(n107), .CK(clk), .Q(wo_2[2]) );
  DFFHQX1 \w_reg[1][2]  ( .D(n106), .CK(clk), .Q(wo_1[2]) );
  DFFHQX1 \w_reg[0][2]  ( .D(n105), .CK(clk), .Q(wo_0[2]) );
  DFFHQX1 \w_reg[2][3]  ( .D(n111), .CK(clk), .Q(wo_2[3]) );
  DFFHQX1 \w_reg[1][3]  ( .D(n110), .CK(clk), .Q(wo_1[3]) );
  DFFHQX1 \w_reg[0][3]  ( .D(n109), .CK(clk), .Q(wo_0[3]) );
  DFFHQX1 \w_reg[2][4]  ( .D(n115), .CK(clk), .Q(wo_2[4]) );
  DFFHQX1 \w_reg[1][4]  ( .D(n114), .CK(clk), .Q(wo_1[4]) );
  DFFHQX1 \w_reg[0][4]  ( .D(n113), .CK(clk), .Q(wo_0[4]) );
  DFFHQX1 \w_reg[2][5]  ( .D(n119), .CK(clk), .Q(wo_2[5]) );
  DFFHQX1 \w_reg[1][5]  ( .D(n118), .CK(clk), .Q(wo_1[5]) );
  DFFHQX1 \w_reg[0][5]  ( .D(n117), .CK(clk), .Q(wo_0[5]) );
  DFFHQX1 \w_reg[2][6]  ( .D(n123), .CK(clk), .Q(wo_2[6]) );
  DFFHQX1 \w_reg[1][6]  ( .D(n122), .CK(clk), .Q(wo_1[6]) );
  DFFHQX1 \w_reg[0][6]  ( .D(n121), .CK(clk), .Q(wo_0[6]) );
  DFFHQX1 \w_reg[2][7]  ( .D(n127), .CK(clk), .Q(wo_2[7]) );
  DFFHQX1 \w_reg[1][7]  ( .D(n126), .CK(clk), .Q(wo_1[7]) );
  DFFHQX1 \w_reg[0][7]  ( .D(n125), .CK(clk), .Q(wo_0[7]) );
  DFFHQX1 \w_reg[2][31]  ( .D(n31), .CK(clk), .Q(wo_2[31]) );
  DFFHQX1 \w_reg[1][31]  ( .D(n30), .CK(clk), .Q(wo_1[31]) );
  DFFHQX1 \w_reg[2][23]  ( .D(n63), .CK(clk), .Q(wo_2[23]) );
  DFFHQX1 \w_reg[1][23]  ( .D(n62), .CK(clk), .Q(wo_1[23]) );
  DFFHQX1 \w_reg[0][23]  ( .D(n61), .CK(clk), .Q(wo_0[23]) );
  DFFHQX1 \w_reg[2][15]  ( .D(n95), .CK(clk), .Q(wo_2[15]) );
  DFFHQX1 \w_reg[1][15]  ( .D(n94), .CK(clk), .Q(wo_1[15]) );
  DFFHQX1 \w_reg[0][15]  ( .D(n93), .CK(clk), .Q(wo_0[15]) );
  DFFHQX1 \w_reg[0][24]  ( .D(n1), .CK(clk), .Q(wo_0[24]) );
  DFFHQX1 \w_reg[0][25]  ( .D(n5), .CK(clk), .Q(wo_0[25]) );
  DFFHQX1 \w_reg[0][26]  ( .D(n9), .CK(clk), .Q(wo_0[26]) );
  DFFHQX1 \w_reg[0][27]  ( .D(n13), .CK(clk), .Q(wo_0[27]) );
  DFFHQX1 \w_reg[0][28]  ( .D(n17), .CK(clk), .Q(wo_0[28]) );
  DFFHQX1 \w_reg[0][29]  ( .D(n21), .CK(clk), .Q(wo_0[29]) );
  DFFHQX1 \w_reg[0][30]  ( .D(n25), .CK(clk), .Q(wo_0[30]) );
  DFFHQX1 \w_reg[0][31]  ( .D(n29), .CK(clk), .Q(wo_0[31]) );
  XOR2X1 U260 ( .A(wo_3[0]), .B(N173), .Y(N239) );
  XOR2X1 U285 ( .A(wo_3[5]), .B(N168), .Y(N234) );
  XOR2X1 U270 ( .A(wo_3[2]), .B(N171), .Y(N237) );
  XOR2X1 U295 ( .A(wo_3[7]), .B(N166), .Y(N232) );
  XOR2X1 U290 ( .A(wo_3[6]), .B(N167), .Y(N233) );
  XOR2X1 U265 ( .A(wo_3[1]), .B(N172), .Y(N238) );
  XOR2X1 U280 ( .A(wo_3[4]), .B(N169), .Y(N235) );
  XOR2X1 U300 ( .A(wo_3[8]), .B(N165), .Y(N231) );
  XOR2X1 U340 ( .A(wo_3[16]), .B(N157), .Y(N223) );
  XOR2X1 U325 ( .A(wo_3[13]), .B(N160), .Y(N226) );
  XOR2X1 U365 ( .A(wo_3[21]), .B(N152), .Y(N218) );
  XOR2X1 U310 ( .A(wo_3[10]), .B(N163), .Y(N229) );
  XOR2X1 U350 ( .A(wo_3[18]), .B(N155), .Y(N221) );
  XOR2X1 U335 ( .A(wo_3[15]), .B(N158), .Y(N224) );
  XOR2X1 U375 ( .A(wo_3[23]), .B(N150), .Y(N216) );
  XOR2X1 U330 ( .A(wo_3[14]), .B(N159), .Y(N225) );
  XOR2X1 U370 ( .A(wo_3[22]), .B(N151), .Y(N217) );
  XOR2X1 U305 ( .A(wo_3[9]), .B(N164), .Y(N230) );
  XOR2X1 U320 ( .A(wo_3[12]), .B(N161), .Y(N227) );
  XOR2X1 U360 ( .A(wo_3[20]), .B(N153), .Y(N219) );
  XOR2X1 U345 ( .A(wo_3[17]), .B(N156), .Y(N222) );
  XOR2X1 U405 ( .A(wo_3[29]), .B(N144), .Y(N210) );
  XOR2X1 U415 ( .A(wo_3[31]), .B(N142), .Y(N208) );
  XOR2X1 U410 ( .A(wo_3[30]), .B(N143), .Y(N209) );
  XOR2X1 U385 ( .A(wo_3[25]), .B(N148), .Y(N214) );
  XOR2X1 U400 ( .A(wo_3[28]), .B(N145), .Y(N211) );
  XOR2X1 U315 ( .A(wo_3[11]), .B(N162), .Y(N228) );
  XOR2X1 U355 ( .A(wo_3[19]), .B(N154), .Y(N220) );
  XOR2X1 U275 ( .A(wo_3[3]), .B(N170), .Y(N236) );
  XOR2X1 U333 ( .A(wo_0[14]), .B(subword[14]), .Y(N27) );
  XOR2X1 U373 ( .A(wo_0[22]), .B(subword[22]), .Y(N19) );
  XOR2X1 U293 ( .A(wo_0[6]), .B(subword[6]), .Y(N35) );
  XOR2X1 U388 ( .A(wo_0[25]), .B(subword[25]), .Y(n264) );
  XOR2X1 U389 ( .A(rcon[25]), .B(n264), .Y(N16) );
  XOR2X1 U408 ( .A(wo_0[29]), .B(subword[29]), .Y(n260) );
  XOR2X1 U409 ( .A(rcon[29]), .B(n260), .Y(N12) );
  XOR2X1 U403 ( .A(wo_0[28]), .B(subword[28]), .Y(n261) );
  XOR2X1 U404 ( .A(rcon[28]), .B(n261), .Y(N13) );
  XOR2X1 U418 ( .A(wo_0[31]), .B(subword[31]), .Y(n258) );
  XOR2X1 U419 ( .A(rcon[31]), .B(n258), .Y(N10) );
  XOR2X1 U413 ( .A(wo_0[30]), .B(subword[30]), .Y(n259) );
  XOR2X1 U414 ( .A(rcon[30]), .B(n259), .Y(N11) );
  XOR2X1 U261 ( .A(wo_2[0]), .B(N107), .Y(N173) );
  XOR2X1 U301 ( .A(wo_2[8]), .B(N99), .Y(N165) );
  XOR2X1 U341 ( .A(wo_2[16]), .B(N91), .Y(N157) );
  XOR2X1 U326 ( .A(wo_2[13]), .B(N94), .Y(N160) );
  XOR2X1 U366 ( .A(wo_2[21]), .B(N86), .Y(N152) );
  XOR2X1 U406 ( .A(wo_2[29]), .B(N78), .Y(N144) );
  XOR2X1 U286 ( .A(wo_2[5]), .B(N102), .Y(N168) );
  XOR2X1 U311 ( .A(wo_2[10]), .B(N97), .Y(N163) );
  XOR2X1 U351 ( .A(wo_2[18]), .B(N89), .Y(N155) );
  XOR2X1 U271 ( .A(wo_2[2]), .B(N105), .Y(N171) );
  XOR2X1 U336 ( .A(wo_2[15]), .B(N92), .Y(N158) );
  XOR2X1 U376 ( .A(wo_2[23]), .B(N84), .Y(N150) );
  XOR2X1 U416 ( .A(wo_2[31]), .B(N76), .Y(N142) );
  XOR2X1 U296 ( .A(wo_2[7]), .B(N100), .Y(N166) );
  XOR2X1 U316 ( .A(wo_2[11]), .B(N96), .Y(N162) );
  XOR2X1 U356 ( .A(wo_2[19]), .B(N88), .Y(N154) );
  XOR2X1 U276 ( .A(wo_2[3]), .B(N104), .Y(N170) );
  XOR2X1 U331 ( .A(wo_2[14]), .B(N93), .Y(N159) );
  XOR2X1 U371 ( .A(wo_2[22]), .B(N85), .Y(N151) );
  XOR2X1 U411 ( .A(wo_2[30]), .B(N77), .Y(N143) );
  XOR2X1 U291 ( .A(wo_2[6]), .B(N101), .Y(N167) );
  XOR2X1 U306 ( .A(wo_2[9]), .B(N98), .Y(N164) );
  XOR2X1 U386 ( .A(wo_2[25]), .B(N82), .Y(N148) );
  XOR2X1 U266 ( .A(wo_2[1]), .B(N106), .Y(N172) );
  XOR2X1 U321 ( .A(wo_2[12]), .B(N95), .Y(N161) );
  XOR2X1 U361 ( .A(wo_2[20]), .B(N87), .Y(N153) );
  XOR2X1 U401 ( .A(wo_2[28]), .B(N79), .Y(N145) );
  XOR2X1 U281 ( .A(wo_2[4]), .B(N103), .Y(N169) );
  XOR2X1 U346 ( .A(wo_2[17]), .B(N90), .Y(N156) );
  XOR2X1 U262 ( .A(wo_1[0]), .B(N41), .Y(N107) );
  XOR2X1 U302 ( .A(wo_1[8]), .B(N33), .Y(N99) );
  XOR2X1 U342 ( .A(wo_1[16]), .B(N25), .Y(N91) );
  XOR2X1 U327 ( .A(wo_1[13]), .B(N28), .Y(N94) );
  XOR2X1 U367 ( .A(wo_1[21]), .B(N20), .Y(N86) );
  XOR2X1 U287 ( .A(wo_1[5]), .B(N36), .Y(N102) );
  XOR2X1 U312 ( .A(wo_1[10]), .B(N31), .Y(N97) );
  XOR2X1 U352 ( .A(wo_1[18]), .B(N23), .Y(N89) );
  XOR2X1 U272 ( .A(wo_1[2]), .B(N39), .Y(N105) );
  XOR2X1 U317 ( .A(wo_1[11]), .B(N30), .Y(N96) );
  XOR2X1 U357 ( .A(wo_1[19]), .B(N22), .Y(N88) );
  XOR2X1 U277 ( .A(wo_1[3]), .B(N38), .Y(N104) );
  XOR2X1 U307 ( .A(wo_1[9]), .B(N32), .Y(N98) );
  XOR2X1 U267 ( .A(wo_1[1]), .B(N40), .Y(N106) );
  XOR2X1 U322 ( .A(wo_1[12]), .B(N29), .Y(N95) );
  XOR2X1 U362 ( .A(wo_1[20]), .B(N21), .Y(N87) );
  XOR2X1 U282 ( .A(wo_1[4]), .B(N37), .Y(N103) );
  XOR2X1 U347 ( .A(wo_1[17]), .B(N24), .Y(N90) );
  XOR2X1 U407 ( .A(wo_1[29]), .B(N12), .Y(N78) );
  XOR2X1 U337 ( .A(wo_1[15]), .B(N26), .Y(N92) );
  XOR2X1 U377 ( .A(wo_1[23]), .B(N18), .Y(N84) );
  XOR2X1 U417 ( .A(wo_1[31]), .B(N10), .Y(N76) );
  XOR2X1 U297 ( .A(wo_1[7]), .B(N34), .Y(N100) );
  XOR2X1 U332 ( .A(wo_1[14]), .B(N27), .Y(N93) );
  XOR2X1 U372 ( .A(wo_1[22]), .B(N19), .Y(N85) );
  XOR2X1 U412 ( .A(wo_1[30]), .B(N11), .Y(N77) );
  XOR2X1 U292 ( .A(wo_1[6]), .B(N35), .Y(N101) );
  XOR2X1 U387 ( .A(wo_1[25]), .B(N16), .Y(N82) );
  XOR2X1 U402 ( .A(wo_1[28]), .B(N13), .Y(N79) );
  XOR2X1 U328 ( .A(wo_0[13]), .B(subword[13]), .Y(N28) );
  XOR2X1 U368 ( .A(wo_0[21]), .B(subword[21]), .Y(N20) );
  XOR2X1 U288 ( .A(wo_0[5]), .B(subword[5]), .Y(N36) );
  XOR2X1 U318 ( .A(wo_0[11]), .B(subword[11]), .Y(N30) );
  XOR2X1 U358 ( .A(wo_0[19]), .B(subword[19]), .Y(N22) );
  XOR2X1 U278 ( .A(wo_0[3]), .B(subword[3]), .Y(N38) );
  XOR2X1 U308 ( .A(wo_0[9]), .B(subword[9]), .Y(N32) );
  XOR2X1 U268 ( .A(wo_0[1]), .B(subword[1]), .Y(N40) );
  XOR2X1 U348 ( .A(wo_0[17]), .B(subword[17]), .Y(N24) );
  XOR2X1 U338 ( .A(wo_0[15]), .B(subword[15]), .Y(N26) );
  XOR2X1 U378 ( .A(wo_0[23]), .B(subword[23]), .Y(N18) );
  XOR2X1 U298 ( .A(wo_0[7]), .B(subword[7]), .Y(N34) );
  XOR2X1 U313 ( .A(wo_0[10]), .B(subword[10]), .Y(N31) );
  XOR2X1 U353 ( .A(wo_0[18]), .B(subword[18]), .Y(N23) );
  XOR2X1 U273 ( .A(wo_0[2]), .B(subword[2]), .Y(N39) );
  XOR2X1 U323 ( .A(wo_0[12]), .B(subword[12]), .Y(N29) );
  XOR2X1 U363 ( .A(wo_0[20]), .B(subword[20]), .Y(N21) );
  XOR2X1 U283 ( .A(wo_0[4]), .B(subword[4]), .Y(N37) );
  XOR2X1 U263 ( .A(wo_0[0]), .B(subword[0]), .Y(N41) );
  XOR2X1 U303 ( .A(wo_0[8]), .B(subword[8]), .Y(N33) );
  XOR2X1 U343 ( .A(wo_0[16]), .B(subword[16]), .Y(N25) );
  XOR2X1 U380 ( .A(wo_3[24]), .B(N149), .Y(N215) );
  XOR2X1 U390 ( .A(wo_3[26]), .B(N147), .Y(N213) );
  XOR2X1 U395 ( .A(wo_3[27]), .B(N146), .Y(N212) );
  XOR2X1 U398 ( .A(wo_0[27]), .B(subword[27]), .Y(n262) );
  XOR2X1 U399 ( .A(rcon[27]), .B(n262), .Y(N14) );
  XOR2X1 U383 ( .A(wo_0[24]), .B(subword[24]), .Y(n265) );
  XOR2X1 U384 ( .A(rcon[24]), .B(n265), .Y(N17) );
  XOR2X1 U393 ( .A(wo_0[26]), .B(subword[26]), .Y(n263) );
  XOR2X1 U394 ( .A(rcon[26]), .B(n263), .Y(N15) );
  XOR2X1 U381 ( .A(wo_2[24]), .B(N83), .Y(N149) );
  XOR2X1 U391 ( .A(wo_2[26]), .B(N81), .Y(N147) );
  XOR2X1 U396 ( .A(wo_2[27]), .B(N80), .Y(N146) );
  XOR2X1 U382 ( .A(wo_1[24]), .B(N17), .Y(N83) );
  XOR2X1 U392 ( .A(wo_1[26]), .B(N15), .Y(N81) );
  XOR2X1 U397 ( .A(wo_1[27]), .B(N14), .Y(N80) );
  DFFHQX1 \w_reg[3][14]  ( .D(n92), .CK(clk), .Q(wo_3[14]) );
  DFFHQX1 \w_reg[3][22]  ( .D(n60), .CK(clk), .Q(wo_3[22]) );
  DFFHQX1 \w_reg[3][30]  ( .D(n28), .CK(clk), .Q(wo_3[30]) );
  DFFHQX1 \w_reg[3][6]  ( .D(n124), .CK(clk), .Q(wo_3[6]) );
  DFFHQX1 \w_reg[3][13]  ( .D(n88), .CK(clk), .Q(wo_3[13]) );
  DFFHQX1 \w_reg[3][29]  ( .D(n24), .CK(clk), .Q(wo_3[29]) );
  DFFHQX1 \w_reg[3][5]  ( .D(n120), .CK(clk), .Q(wo_3[5]) );
  DFFHQX1 \w_reg[3][21]  ( .D(n56), .CK(clk), .Q(wo_3[21]) );
  DFFHQX1 \w_reg[3][9]  ( .D(n72), .CK(clk), .Q(wo_3[9]) );
  DFFHQX1 \w_reg[3][25]  ( .D(n8), .CK(clk), .Q(wo_3[25]) );
  DFFHQX1 \w_reg[3][1]  ( .D(n104), .CK(clk), .Q(wo_3[1]) );
  DFFHQX1 \w_reg[3][17]  ( .D(n40), .CK(clk), .Q(wo_3[17]) );
  DFFHQX1 \w_reg[3][15]  ( .D(n96), .CK(clk), .Q(wo_3[15]) );
  DFFHQX1 \w_reg[3][31]  ( .D(n32), .CK(clk), .Q(wo_3[31]) );
  DFFHQX1 \w_reg[3][7]  ( .D(n128), .CK(clk), .Q(wo_3[7]) );
  DFFHQX1 \w_reg[3][23]  ( .D(n64), .CK(clk), .Q(wo_3[23]) );
  DFFHQX1 \w_reg[3][12]  ( .D(n84), .CK(clk), .Q(wo_3[12]) );
  DFFHQX1 \w_reg[3][4]  ( .D(n116), .CK(clk), .Q(wo_3[4]) );
  DFFHQX1 \w_reg[3][20]  ( .D(n52), .CK(clk), .Q(wo_3[20]) );
  DFFHQX1 \w_reg[3][0]  ( .D(n100), .CK(clk), .Q(wo_3[0]) );
  DFFHQX1 \w_reg[3][16]  ( .D(n36), .CK(clk), .Q(wo_3[16]) );
  DFFHQX1 \w_reg[3][8]  ( .D(n68), .CK(clk), .Q(wo_3[8]) );
  DFFHQX1 \w_reg[3][18]  ( .D(n44), .CK(clk), .Q(wo_3[18]) );
  DFFHQX1 \w_reg[3][28]  ( .D(n20), .CK(clk), .Q(wo_3[28]) );
  DFFHQX1 \w_reg[3][24]  ( .D(n4), .CK(clk), .Q(wo_3[24]) );
  DFFHQX1 \w_reg[3][3]  ( .D(n112), .CK(clk), .Q(wo_3[3]) );
  DFFHQX1 \w_reg[3][19]  ( .D(n48), .CK(clk), .Q(wo_3[19]) );
  DFFHQX1 \w_reg[3][11]  ( .D(n80), .CK(clk), .Q(wo_3[11]) );
  DFFHQX1 \w_reg[3][27]  ( .D(n16), .CK(clk), .Q(wo_3[27]) );
  DFFHQX1 \w_reg[3][2]  ( .D(n108), .CK(clk), .Q(wo_3[2]) );
  DFFHQX1 \w_reg[3][10]  ( .D(n76), .CK(clk), .Q(wo_3[10]) );
  DFFHQX1 \w_reg[3][26]  ( .D(n12), .CK(clk), .Q(wo_3[26]) );
  INVX12 U3 ( .A(n438), .Y(n370) );
  INVX12 U4 ( .A(n438), .Y(n371) );
  INVX8 U5 ( .A(n438), .Y(n372) );
  INVX8 U6 ( .A(n438), .Y(n373) );
  CLKINVX3 U7 ( .A(n439), .Y(n438) );
  INVX1 U8 ( .A(n453), .Y(n387) );
  INVX1 U9 ( .A(n454), .Y(n385) );
  INVX1 U10 ( .A(n455), .Y(n383) );
  INVX1 U11 ( .A(n468), .Y(n421) );
  INVX1 U12 ( .A(n441), .Y(n420) );
  INVX1 U13 ( .A(n448), .Y(n405) );
  INVX1 U14 ( .A(n449), .Y(n404) );
  INVX1 U15 ( .A(n469), .Y(n389) );
  INVX1 U16 ( .A(n453), .Y(n388) );
  INVX1 U17 ( .A(n439), .Y(n437) );
  INVX1 U18 ( .A(n440), .Y(n436) );
  INVX1 U19 ( .A(n440), .Y(n435) );
  INVX1 U20 ( .A(n450), .Y(n434) );
  INVX1 U21 ( .A(n451), .Y(n433) );
  INVX1 U22 ( .A(n442), .Y(n432) );
  INVX1 U23 ( .A(n443), .Y(n431) );
  INVX1 U24 ( .A(n467), .Y(n430) );
  INVX1 U25 ( .A(n440), .Y(n429) );
  INVX1 U26 ( .A(n467), .Y(n428) );
  INVX1 U27 ( .A(n470), .Y(n427) );
  INVX1 U28 ( .A(n456), .Y(n426) );
  INVX1 U29 ( .A(n457), .Y(n425) );
  INVX1 U30 ( .A(n472), .Y(n424) );
  INVX1 U31 ( .A(n460), .Y(n423) );
  INVX1 U32 ( .A(n441), .Y(n422) );
  INVX1 U33 ( .A(n454), .Y(n386) );
  INVX1 U34 ( .A(n455), .Y(n384) );
  INVX1 U35 ( .A(n456), .Y(n382) );
  INVX1 U36 ( .A(n456), .Y(n381) );
  INVX1 U37 ( .A(n457), .Y(n380) );
  INVX1 U38 ( .A(n457), .Y(n379) );
  INVX1 U39 ( .A(n449), .Y(n403) );
  INVX1 U40 ( .A(n450), .Y(n402) );
  INVX1 U41 ( .A(n450), .Y(n401) );
  INVX1 U42 ( .A(n451), .Y(n400) );
  INVX1 U43 ( .A(n451), .Y(n399) );
  INVX1 U44 ( .A(n452), .Y(n398) );
  INVX1 U45 ( .A(n452), .Y(n397) );
  INVX1 U46 ( .A(n471), .Y(n396) );
  INVX1 U47 ( .A(n455), .Y(n395) );
  INVX1 U48 ( .A(n470), .Y(n394) );
  INVX1 U49 ( .A(n452), .Y(n393) );
  INVX1 U50 ( .A(n467), .Y(n392) );
  INVX1 U51 ( .A(n468), .Y(n391) );
  INVX1 U52 ( .A(n444), .Y(n390) );
  INVX1 U53 ( .A(n441), .Y(n419) );
  INVX1 U54 ( .A(n442), .Y(n418) );
  INVX1 U55 ( .A(n442), .Y(n417) );
  INVX1 U56 ( .A(n443), .Y(n416) );
  INVX1 U57 ( .A(n443), .Y(n415) );
  INVX1 U58 ( .A(n444), .Y(n414) );
  INVX1 U59 ( .A(n444), .Y(n413) );
  INVX1 U60 ( .A(n445), .Y(n412) );
  INVX1 U61 ( .A(n445), .Y(n411) );
  INVX1 U62 ( .A(n446), .Y(n410) );
  INVX1 U63 ( .A(n446), .Y(n409) );
  INVX1 U64 ( .A(n447), .Y(n408) );
  INVX1 U65 ( .A(n447), .Y(n407) );
  INVX1 U66 ( .A(n448), .Y(n406) );
  INVX1 U67 ( .A(n459), .Y(n375) );
  INVX1 U68 ( .A(n458), .Y(n378) );
  INVX1 U69 ( .A(n458), .Y(n377) );
  INVX1 U70 ( .A(n459), .Y(n376) );
  INVX1 U71 ( .A(n427), .Y(n439) );
  INVX1 U72 ( .A(n392), .Y(n453) );
  INVX1 U73 ( .A(n434), .Y(n440) );
  INVX1 U74 ( .A(n430), .Y(n454) );
  INVX1 U75 ( .A(n462), .Y(n455) );
  INVX1 U76 ( .A(n462), .Y(n456) );
  INVX1 U77 ( .A(n462), .Y(n457) );
  INVX1 U78 ( .A(n464), .Y(n449) );
  INVX1 U79 ( .A(n463), .Y(n450) );
  INVX1 U80 ( .A(n463), .Y(n451) );
  INVX1 U81 ( .A(n463), .Y(n452) );
  INVX1 U82 ( .A(n466), .Y(n441) );
  INVX1 U83 ( .A(n466), .Y(n442) );
  INVX1 U84 ( .A(n466), .Y(n443) );
  INVX1 U85 ( .A(n465), .Y(n444) );
  INVX1 U86 ( .A(n465), .Y(n445) );
  INVX1 U87 ( .A(n465), .Y(n446) );
  INVX1 U88 ( .A(n464), .Y(n447) );
  INVX1 U89 ( .A(n464), .Y(n448) );
  INVX1 U90 ( .A(n460), .Y(n374) );
  INVX1 U91 ( .A(n461), .Y(n460) );
  INVX1 U92 ( .A(n461), .Y(n458) );
  INVX1 U93 ( .A(n461), .Y(n459) );
  INVX1 U94 ( .A(n471), .Y(n462) );
  INVX1 U95 ( .A(n470), .Y(n463) );
  INVX1 U96 ( .A(n468), .Y(n466) );
  INVX1 U97 ( .A(n469), .Y(n465) );
  INVX1 U98 ( .A(n469), .Y(n464) );
  INVX1 U99 ( .A(n474), .Y(n467) );
  INVX1 U100 ( .A(n473), .Y(n470) );
  INVX1 U101 ( .A(n473), .Y(n471) );
  INVX1 U102 ( .A(n474), .Y(n468) );
  INVX1 U103 ( .A(n474), .Y(n469) );
  INVX1 U104 ( .A(n472), .Y(n461) );
  INVX1 U105 ( .A(n473), .Y(n472) );
  INVX1 U106 ( .A(kld), .Y(n474) );
  INVX1 U107 ( .A(kld), .Y(n473) );
  INVX1 U108 ( .A(n143), .Y(n16) );
  AOI22X1 U109 ( .A0(N212), .A1(n380), .B0(key[27]), .B1(n370), .Y(n143) );
  INVX1 U110 ( .A(n139), .Y(n12) );
  AOI22X1 U111 ( .A0(N213), .A1(n378), .B0(key[26]), .B1(n370), .Y(n139) );
  INVX1 U112 ( .A(n132), .Y(n4) );
  AOI22X1 U113 ( .A0(N215), .A1(n375), .B0(key[24]), .B1(n370), .Y(n132) );
  INVX1 U114 ( .A(n161), .Y(n29) );
  AOI22X1 U115 ( .A0(N10), .A1(n389), .B0(key[127]), .B1(n371), .Y(n161) );
  INVX1 U116 ( .A(n177), .Y(n45) );
  AOI22X1 U117 ( .A0(N22), .A1(n397), .B0(key[115]), .B1(n371), .Y(n177) );
  INVX1 U118 ( .A(n209), .Y(n77) );
  AOI22X1 U119 ( .A0(N30), .A1(n413), .B0(key[107]), .B1(n372), .Y(n209) );
  INVX1 U120 ( .A(n130), .Y(n2) );
  AOI22X1 U121 ( .A0(N83), .A1(n374), .B0(n370), .B1(key[88]), .Y(n130) );
  INVX1 U122 ( .A(n238), .Y(n112) );
  AOI22X1 U123 ( .A0(N236), .A1(n428), .B0(key[3]), .B1(n373), .Y(n238) );
  INVX1 U124 ( .A(n175), .Y(n48) );
  AOI22X1 U125 ( .A0(N220), .A1(n396), .B0(key[19]), .B1(n371), .Y(n175) );
  INVX1 U126 ( .A(n207), .Y(n80) );
  AOI22X1 U127 ( .A0(N228), .A1(n412), .B0(key[11]), .B1(n372), .Y(n207) );
  INVX1 U128 ( .A(n148), .Y(n20) );
  AOI22X1 U129 ( .A0(N211), .A1(n383), .B0(key[28]), .B1(n370), .Y(n148) );
  INVX1 U130 ( .A(n135), .Y(n8) );
  AOI22X1 U131 ( .A0(N214), .A1(n376), .B0(key[25]), .B1(n370), .Y(n135) );
  INVX1 U132 ( .A(n156), .Y(n28) );
  AOI22X1 U133 ( .A0(N209), .A1(n387), .B0(key[30]), .B1(n370), .Y(n156) );
  INVX1 U134 ( .A(n159), .Y(n32) );
  AOI22X1 U135 ( .A0(N208), .A1(n388), .B0(key[31]), .B1(n370), .Y(n159) );
  INVX1 U136 ( .A(n152), .Y(n24) );
  AOI22X1 U137 ( .A0(N210), .A1(n385), .B0(key[29]), .B1(n370), .Y(n152) );
  INVX1 U138 ( .A(n157), .Y(n25) );
  AOI22X1 U139 ( .A0(N11), .A1(n387), .B0(key[126]), .B1(n370), .Y(n157) );
  INVX1 U140 ( .A(n153), .Y(n21) );
  AOI22X1 U141 ( .A0(N12), .A1(n385), .B0(key[125]), .B1(n370), .Y(n153) );
  INVX1 U142 ( .A(n149), .Y(n17) );
  AOI22X1 U143 ( .A0(N13), .A1(n383), .B0(key[124]), .B1(n370), .Y(n149) );
  INVX1 U144 ( .A(n145), .Y(n13) );
  AOI22X1 U145 ( .A0(N14), .A1(n381), .B0(key[123]), .B1(n370), .Y(n145) );
  INVX1 U146 ( .A(n141), .Y(n9) );
  AOI22X1 U147 ( .A0(N15), .A1(n379), .B0(key[122]), .B1(n370), .Y(n141) );
  INVX1 U148 ( .A(n137), .Y(n5) );
  AOI22X1 U149 ( .A0(N16), .A1(n377), .B0(key[121]), .B1(n370), .Y(n137) );
  INVX1 U150 ( .A(n133), .Y(n1) );
  AOI22X1 U151 ( .A0(N17), .A1(n375), .B0(key[120]), .B1(n370), .Y(n133) );
  INVX1 U152 ( .A(n158), .Y(n31) );
  AOI22X1 U153 ( .A0(N142), .A1(n388), .B0(key[63]), .B1(n370), .Y(n158) );
  INVX1 U154 ( .A(n154), .Y(n26) );
  AOI22X1 U155 ( .A0(N77), .A1(n386), .B0(key[94]), .B1(n370), .Y(n154) );
  INVX1 U156 ( .A(n155), .Y(n27) );
  AOI22X1 U157 ( .A0(N143), .A1(n386), .B0(key[62]), .B1(n370), .Y(n155) );
  INVX1 U158 ( .A(n150), .Y(n22) );
  AOI22X1 U159 ( .A0(N78), .A1(n384), .B0(key[93]), .B1(n370), .Y(n150) );
  INVX1 U160 ( .A(n151), .Y(n23) );
  AOI22X1 U161 ( .A0(N144), .A1(n384), .B0(key[61]), .B1(n370), .Y(n151) );
  INVX1 U162 ( .A(n146), .Y(n18) );
  AOI22X1 U163 ( .A0(N79), .A1(n382), .B0(key[92]), .B1(n370), .Y(n146) );
  INVX1 U164 ( .A(n147), .Y(n19) );
  AOI22X1 U165 ( .A0(N145), .A1(n382), .B0(key[60]), .B1(n370), .Y(n147) );
  INVX1 U166 ( .A(n144), .Y(n14) );
  AOI22X1 U167 ( .A0(N80), .A1(n381), .B0(key[91]), .B1(n370), .Y(n144) );
  INVX1 U168 ( .A(n142), .Y(n15) );
  AOI22X1 U169 ( .A0(N146), .A1(n380), .B0(key[59]), .B1(n370), .Y(n142) );
  INVX1 U170 ( .A(n140), .Y(n10) );
  AOI22X1 U171 ( .A0(N81), .A1(n379), .B0(key[90]), .B1(n370), .Y(n140) );
  INVX1 U172 ( .A(n138), .Y(n11) );
  AOI22X1 U173 ( .A0(N147), .A1(n378), .B0(key[58]), .B1(n370), .Y(n138) );
  INVX1 U174 ( .A(n136), .Y(n6) );
  AOI22X1 U175 ( .A0(N82), .A1(n377), .B0(key[89]), .B1(n370), .Y(n136) );
  INVX1 U176 ( .A(n134), .Y(n7) );
  AOI22X1 U177 ( .A0(N148), .A1(n376), .B0(key[57]), .B1(n370), .Y(n134) );
  INVX1 U178 ( .A(n131), .Y(n3) );
  AOI22X1 U179 ( .A0(N149), .A1(n374), .B0(key[56]), .B1(n370), .Y(n131) );
  INVX1 U180 ( .A(n166), .Y(n40) );
  AOI22X1 U181 ( .A0(N222), .A1(n392), .B0(key[17]), .B1(n371), .Y(n166) );
  INVX1 U182 ( .A(n179), .Y(n52) );
  AOI22X1 U183 ( .A0(N219), .A1(n398), .B0(key[20]), .B1(n371), .Y(n179) );
  INVX1 U184 ( .A(n211), .Y(n84) );
  AOI22X1 U185 ( .A0(N227), .A1(n414), .B0(key[12]), .B1(n372), .Y(n211) );
  INVX1 U186 ( .A(n198), .Y(n72) );
  AOI22X1 U187 ( .A0(N230), .A1(n408), .B0(key[9]), .B1(n372), .Y(n198) );
  INVX1 U188 ( .A(n187), .Y(n60) );
  AOI22X1 U189 ( .A0(N217), .A1(n402), .B0(key[22]), .B1(n371), .Y(n187) );
  INVX1 U190 ( .A(n219), .Y(n92) );
  AOI22X1 U191 ( .A0(N225), .A1(n418), .B0(key[14]), .B1(n372), .Y(n219) );
  INVX1 U192 ( .A(n190), .Y(n64) );
  AOI22X1 U193 ( .A0(N216), .A1(n404), .B0(key[23]), .B1(n371), .Y(n190) );
  INVX1 U194 ( .A(n222), .Y(n96) );
  AOI22X1 U195 ( .A0(N224), .A1(n420), .B0(key[15]), .B1(n372), .Y(n222) );
  INVX1 U196 ( .A(n171), .Y(n44) );
  AOI22X1 U197 ( .A0(N221), .A1(n394), .B0(key[18]), .B1(n371), .Y(n171) );
  INVX1 U198 ( .A(n203), .Y(n76) );
  AOI22X1 U199 ( .A0(N229), .A1(n410), .B0(key[10]), .B1(n372), .Y(n203) );
  INVX1 U200 ( .A(n183), .Y(n56) );
  AOI22X1 U201 ( .A0(N218), .A1(n400), .B0(key[21]), .B1(n371), .Y(n183) );
  INVX1 U202 ( .A(n215), .Y(n88) );
  AOI22X1 U203 ( .A0(N226), .A1(n416), .B0(key[13]), .B1(n372), .Y(n215) );
  INVX1 U204 ( .A(n163), .Y(n36) );
  AOI22X1 U205 ( .A0(N223), .A1(n390), .B0(key[16]), .B1(n371), .Y(n163) );
  INVX1 U206 ( .A(n195), .Y(n68) );
  AOI22X1 U207 ( .A0(N231), .A1(n406), .B0(key[8]), .B1(n372), .Y(n195) );
  INVX1 U208 ( .A(n224), .Y(n94) );
  AOI22X1 U209 ( .A0(N92), .A1(n421), .B0(key[79]), .B1(n372), .Y(n224) );
  INVX1 U210 ( .A(n223), .Y(n95) );
  AOI22X1 U211 ( .A0(N158), .A1(n420), .B0(key[47]), .B1(n372), .Y(n223) );
  INVX1 U212 ( .A(n192), .Y(n62) );
  AOI22X1 U213 ( .A0(N84), .A1(n405), .B0(key[87]), .B1(n371), .Y(n192) );
  INVX1 U214 ( .A(n191), .Y(n63) );
  AOI22X1 U215 ( .A0(N150), .A1(n404), .B0(key[55]), .B1(n371), .Y(n191) );
  INVX1 U216 ( .A(n160), .Y(n30) );
  AOI22X1 U217 ( .A0(N76), .A1(n389), .B0(key[95]), .B1(n371), .Y(n160) );
  INVX1 U218 ( .A(n188), .Y(n58) );
  AOI22X1 U219 ( .A0(N85), .A1(n403), .B0(key[86]), .B1(n371), .Y(n188) );
  INVX1 U220 ( .A(n186), .Y(n59) );
  AOI22X1 U221 ( .A0(N151), .A1(n402), .B0(key[54]), .B1(n371), .Y(n186) );
  INVX1 U222 ( .A(n184), .Y(n54) );
  AOI22X1 U223 ( .A0(N86), .A1(n401), .B0(key[85]), .B1(n371), .Y(n184) );
  INVX1 U224 ( .A(n182), .Y(n55) );
  AOI22X1 U225 ( .A0(N152), .A1(n400), .B0(key[53]), .B1(n371), .Y(n182) );
  INVX1 U226 ( .A(n180), .Y(n50) );
  AOI22X1 U227 ( .A0(N87), .A1(n399), .B0(key[84]), .B1(n371), .Y(n180) );
  INVX1 U228 ( .A(n178), .Y(n51) );
  AOI22X1 U229 ( .A0(N153), .A1(n398), .B0(key[52]), .B1(n371), .Y(n178) );
  INVX1 U230 ( .A(n176), .Y(n46) );
  AOI22X1 U231 ( .A0(N88), .A1(n397), .B0(key[83]), .B1(n371), .Y(n176) );
  INVX1 U232 ( .A(n174), .Y(n47) );
  AOI22X1 U233 ( .A0(N154), .A1(n396), .B0(key[51]), .B1(n371), .Y(n174) );
  INVX1 U234 ( .A(n172), .Y(n42) );
  AOI22X1 U235 ( .A0(N89), .A1(n395), .B0(key[82]), .B1(n371), .Y(n172) );
  INVX1 U236 ( .A(n170), .Y(n43) );
  AOI22X1 U237 ( .A0(N155), .A1(n394), .B0(key[50]), .B1(n371), .Y(n170) );
  INVX1 U238 ( .A(n168), .Y(n38) );
  AOI22X1 U239 ( .A0(N90), .A1(n393), .B0(key[81]), .B1(n371), .Y(n168) );
  INVX1 U240 ( .A(n167), .Y(n39) );
  AOI22X1 U241 ( .A0(N156), .A1(n392), .B0(key[49]), .B1(n371), .Y(n167) );
  INVX1 U242 ( .A(n164), .Y(n34) );
  AOI22X1 U243 ( .A0(N91), .A1(n391), .B0(key[80]), .B1(n371), .Y(n164) );
  INVX1 U244 ( .A(n162), .Y(n35) );
  AOI22X1 U245 ( .A0(N157), .A1(n390), .B0(key[48]), .B1(n372), .Y(n162) );
  INVX1 U246 ( .A(n220), .Y(n90) );
  AOI22X1 U247 ( .A0(N93), .A1(n419), .B0(key[78]), .B1(n372), .Y(n220) );
  INVX1 U248 ( .A(n218), .Y(n91) );
  AOI22X1 U249 ( .A0(N159), .A1(n418), .B0(key[46]), .B1(n372), .Y(n218) );
  INVX1 U250 ( .A(n216), .Y(n86) );
  AOI22X1 U251 ( .A0(N94), .A1(n417), .B0(key[77]), .B1(n372), .Y(n216) );
  INVX1 U252 ( .A(n214), .Y(n87) );
  AOI22X1 U253 ( .A0(N160), .A1(n416), .B0(key[45]), .B1(n372), .Y(n214) );
  INVX1 U254 ( .A(n212), .Y(n82) );
  AOI22X1 U255 ( .A0(N95), .A1(n415), .B0(key[76]), .B1(n372), .Y(n212) );
  INVX1 U256 ( .A(n210), .Y(n83) );
  AOI22X1 U257 ( .A0(N161), .A1(n414), .B0(key[44]), .B1(n372), .Y(n210) );
  INVX1 U258 ( .A(n208), .Y(n78) );
  AOI22X1 U259 ( .A0(N96), .A1(n413), .B0(key[75]), .B1(n372), .Y(n208) );
  INVX1 U264 ( .A(n206), .Y(n79) );
  AOI22X1 U269 ( .A0(N162), .A1(n412), .B0(key[43]), .B1(n372), .Y(n206) );
  INVX1 U274 ( .A(n204), .Y(n74) );
  AOI22X1 U279 ( .A0(N97), .A1(n411), .B0(key[74]), .B1(n372), .Y(n204) );
  INVX1 U284 ( .A(n202), .Y(n75) );
  AOI22X1 U289 ( .A0(N163), .A1(n410), .B0(key[42]), .B1(n372), .Y(n202) );
  INVX1 U294 ( .A(n200), .Y(n70) );
  AOI22X1 U299 ( .A0(N98), .A1(n409), .B0(key[73]), .B1(n372), .Y(n200) );
  INVX1 U304 ( .A(n199), .Y(n71) );
  AOI22X1 U309 ( .A0(N164), .A1(n408), .B0(key[41]), .B1(n372), .Y(n199) );
  INVX1 U314 ( .A(n196), .Y(n66) );
  AOI22X1 U319 ( .A0(N99), .A1(n407), .B0(key[72]), .B1(n372), .Y(n196) );
  INVX1 U324 ( .A(n194), .Y(n67) );
  AOI22X1 U329 ( .A0(N165), .A1(n406), .B0(key[40]), .B1(n372), .Y(n194) );
  INVX1 U334 ( .A(n243), .Y(n116) );
  AOI22X1 U339 ( .A0(N235), .A1(n430), .B0(key[4]), .B1(n373), .Y(n243) );
  INVX1 U344 ( .A(n230), .Y(n104) );
  AOI22X1 U349 ( .A0(N238), .A1(n424), .B0(key[1]), .B1(n373), .Y(n230) );
  INVX1 U354 ( .A(n251), .Y(n124) );
  AOI22X1 U359 ( .A0(N233), .A1(n434), .B0(key[6]), .B1(n373), .Y(n251) );
  INVX1 U364 ( .A(n254), .Y(n128) );
  AOI22X1 U369 ( .A0(N232), .A1(n436), .B0(key[7]), .B1(n373), .Y(n254) );
  INVX1 U374 ( .A(n234), .Y(n108) );
  AOI22X1 U379 ( .A0(N237), .A1(n426), .B0(key[2]), .B1(n373), .Y(n234) );
  INVX1 U420 ( .A(n247), .Y(n120) );
  AOI22X1 U421 ( .A0(N234), .A1(n432), .B0(key[5]), .B1(n373), .Y(n247) );
  INVX1 U422 ( .A(n226), .Y(n100) );
  AOI22X1 U423 ( .A0(N239), .A1(n422), .B0(key[0]), .B1(n373), .Y(n226) );
  INVX1 U424 ( .A(n256), .Y(n126) );
  AOI22X1 U425 ( .A0(N100), .A1(n437), .B0(key[71]), .B1(n373), .Y(n256) );
  INVX1 U426 ( .A(n255), .Y(n127) );
  AOI22X1 U427 ( .A0(N166), .A1(n436), .B0(key[39]), .B1(n373), .Y(n255) );
  INVX1 U428 ( .A(n252), .Y(n122) );
  AOI22X1 U429 ( .A0(N101), .A1(n435), .B0(key[70]), .B1(n373), .Y(n252) );
  INVX1 U430 ( .A(n250), .Y(n123) );
  AOI22X1 U431 ( .A0(N167), .A1(n434), .B0(key[38]), .B1(n373), .Y(n250) );
  INVX1 U432 ( .A(n248), .Y(n118) );
  AOI22X1 U433 ( .A0(N102), .A1(n433), .B0(key[69]), .B1(n373), .Y(n248) );
  INVX1 U434 ( .A(n246), .Y(n119) );
  AOI22X1 U435 ( .A0(N168), .A1(n432), .B0(key[37]), .B1(n373), .Y(n246) );
  INVX1 U436 ( .A(n244), .Y(n114) );
  AOI22X1 U437 ( .A0(N103), .A1(n431), .B0(key[68]), .B1(n373), .Y(n244) );
  INVX1 U438 ( .A(n242), .Y(n115) );
  AOI22X1 U439 ( .A0(N169), .A1(n430), .B0(key[36]), .B1(n373), .Y(n242) );
  INVX1 U440 ( .A(n241), .Y(n109) );
  AOI22X1 U441 ( .A0(N38), .A1(n429), .B0(key[99]), .B1(n373), .Y(n241) );
  INVX1 U442 ( .A(n240), .Y(n110) );
  AOI22X1 U443 ( .A0(N104), .A1(n429), .B0(key[67]), .B1(n373), .Y(n240) );
  INVX1 U444 ( .A(n239), .Y(n111) );
  AOI22X1 U445 ( .A0(N170), .A1(n428), .B0(key[35]), .B1(n373), .Y(n239) );
  INVX1 U446 ( .A(n236), .Y(n106) );
  AOI22X1 U447 ( .A0(N105), .A1(n427), .B0(key[66]), .B1(n373), .Y(n236) );
  INVX1 U448 ( .A(n235), .Y(n107) );
  AOI22X1 U449 ( .A0(N171), .A1(n426), .B0(key[34]), .B1(n373), .Y(n235) );
  INVX1 U450 ( .A(n232), .Y(n102) );
  AOI22X1 U451 ( .A0(N106), .A1(n425), .B0(key[65]), .B1(n373), .Y(n232) );
  INVX1 U452 ( .A(n231), .Y(n103) );
  AOI22X1 U453 ( .A0(N172), .A1(n424), .B0(key[33]), .B1(n373), .Y(n231) );
  INVX1 U454 ( .A(n228), .Y(n98) );
  AOI22X1 U455 ( .A0(N107), .A1(n423), .B0(key[64]), .B1(n373), .Y(n228) );
  INVX1 U456 ( .A(n227), .Y(n99) );
  AOI22X1 U457 ( .A0(N173), .A1(n422), .B0(key[32]), .B1(n373), .Y(n227) );
  INVX1 U458 ( .A(n225), .Y(n93) );
  AOI22X1 U459 ( .A0(N26), .A1(n421), .B0(key[111]), .B1(n372), .Y(n225) );
  INVX1 U460 ( .A(n193), .Y(n61) );
  AOI22X1 U461 ( .A0(N18), .A1(n405), .B0(key[119]), .B1(n371), .Y(n193) );
  INVX1 U462 ( .A(n189), .Y(n57) );
  AOI22X1 U463 ( .A0(N19), .A1(n403), .B0(key[118]), .B1(n371), .Y(n189) );
  INVX1 U464 ( .A(n181), .Y(n49) );
  AOI22X1 U465 ( .A0(N21), .A1(n399), .B0(key[116]), .B1(n371), .Y(n181) );
  INVX1 U466 ( .A(n173), .Y(n41) );
  AOI22X1 U467 ( .A0(N23), .A1(n395), .B0(key[114]), .B1(n371), .Y(n173) );
  INVX1 U468 ( .A(n221), .Y(n89) );
  AOI22X1 U469 ( .A0(N27), .A1(n419), .B0(key[110]), .B1(n372), .Y(n221) );
  INVX1 U470 ( .A(n213), .Y(n81) );
  AOI22X1 U471 ( .A0(N29), .A1(n415), .B0(key[108]), .B1(n372), .Y(n213) );
  INVX1 U472 ( .A(n205), .Y(n73) );
  AOI22X1 U473 ( .A0(N31), .A1(n411), .B0(key[106]), .B1(n372), .Y(n205) );
  INVX1 U474 ( .A(n257), .Y(n125) );
  AOI22X1 U475 ( .A0(N34), .A1(n437), .B0(key[103]), .B1(n370), .Y(n257) );
  INVX1 U476 ( .A(n185), .Y(n53) );
  AOI22X1 U477 ( .A0(N20), .A1(n401), .B0(key[117]), .B1(n371), .Y(n185) );
  INVX1 U478 ( .A(n169), .Y(n37) );
  AOI22X1 U479 ( .A0(N24), .A1(n393), .B0(key[113]), .B1(n371), .Y(n169) );
  INVX1 U480 ( .A(n165), .Y(n33) );
  AOI22X1 U481 ( .A0(N25), .A1(n391), .B0(key[112]), .B1(n371), .Y(n165) );
  INVX1 U482 ( .A(n217), .Y(n85) );
  AOI22X1 U483 ( .A0(N28), .A1(n417), .B0(key[109]), .B1(n372), .Y(n217) );
  INVX1 U484 ( .A(n201), .Y(n69) );
  AOI22X1 U485 ( .A0(N32), .A1(n409), .B0(key[105]), .B1(n372), .Y(n201) );
  INVX1 U486 ( .A(n197), .Y(n65) );
  AOI22X1 U487 ( .A0(N33), .A1(n407), .B0(key[104]), .B1(n372), .Y(n197) );
  INVX1 U488 ( .A(n253), .Y(n121) );
  AOI22X1 U489 ( .A0(N35), .A1(n435), .B0(key[102]), .B1(n373), .Y(n253) );
  INVX1 U490 ( .A(n249), .Y(n117) );
  AOI22X1 U491 ( .A0(N36), .A1(n433), .B0(key[101]), .B1(n373), .Y(n249) );
  INVX1 U492 ( .A(n245), .Y(n113) );
  AOI22X1 U493 ( .A0(N37), .A1(n431), .B0(key[100]), .B1(n373), .Y(n245) );
  INVX1 U494 ( .A(n237), .Y(n105) );
  AOI22X1 U495 ( .A0(N39), .A1(n427), .B0(key[98]), .B1(n373), .Y(n237) );
  INVX1 U496 ( .A(n233), .Y(n101) );
  AOI22X1 U497 ( .A0(N40), .A1(n425), .B0(key[97]), .B1(n373), .Y(n233) );
  INVX1 U498 ( .A(n229), .Y(n97) );
  AOI22X1 U499 ( .A0(N41), .A1(n423), .B0(key[96]), .B1(n373), .Y(n229) );
endmodule


module aes_sbox_0 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392;

  OAI221X4 U4 ( .A0(n66), .A1(n372), .B0(n61), .B1(n387), .C0(n84), .Y(n81) );
  OAI221X4 U6 ( .A0(n86), .A1(n87), .B0(n88), .B1(n387), .C0(n89), .Y(n80) );
  OAI222X4 U75 ( .A0(n387), .A1(n207), .B0(n181), .B1(n120), .C0(n381), .C1(
        n208), .Y(n204) );
  OAI32X4 U280 ( .A0(n387), .A1(n56), .A2(n53), .B0(n94), .B1(n103), .Y(n366)
         );
  AOI221X1 U1 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n56), .B(n367), .Y(n229) );
  NAND2X2 U5 ( .A(n368), .B(n66), .Y(n181) );
  NAND2X1 U7 ( .A(n39), .B(n367), .Y(n142) );
  NAND2X2 U8 ( .A(n66), .B(n71), .Y(n138) );
  NAND2X1 U9 ( .A(n368), .B(n371), .Y(n103) );
  NAND2X1 U10 ( .A(n367), .B(n181), .Y(n102) );
  NAND2X2 U11 ( .A(n373), .B(n181), .Y(n113) );
  OAI222X1 U12 ( .A0(n94), .A1(n118), .B0(n119), .B1(n381), .C0(a[4]), .C1(
        n120), .Y(n117) );
  NAND2X2 U13 ( .A(n66), .B(n371), .Y(n116) );
  NAND2X2 U14 ( .A(n367), .B(n368), .Y(n115) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n73) );
  NAND2X1 U16 ( .A(n369), .B(n75), .Y(n110) );
  CLKINVX3 U17 ( .A(n369), .Y(n26) );
  NAND2X2 U18 ( .A(n75), .B(n26), .Y(n154) );
  NAND2X2 U19 ( .A(a[0]), .B(n26), .Y(n156) );
  NAND2X1 U20 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U21 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI21XL U22 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  NAND2X1 U23 ( .A(a[4]), .B(n371), .Y(n263) );
  NAND2X1 U24 ( .A(n367), .B(a[4]), .Y(n224) );
  NAND2X2 U25 ( .A(n368), .B(a[4]), .Y(n111) );
  CLKINVX3 U26 ( .A(a[4]), .Y(n66) );
  NAND2X1 U27 ( .A(n53), .B(n392), .Y(n288) );
  CLKINVX3 U28 ( .A(n379), .Y(n376) );
  INVX1 U29 ( .A(n325), .Y(n34) );
  NAND2X1 U30 ( .A(n113), .B(n371), .Y(n214) );
  NAND2X1 U31 ( .A(n46), .B(n371), .Y(n209) );
  NAND2X1 U32 ( .A(n50), .B(n371), .Y(n301) );
  NAND2X1 U33 ( .A(n374), .B(n268), .Y(n212) );
  NAND2X1 U34 ( .A(n147), .B(n214), .Y(n207) );
  NAND2X1 U35 ( .A(n115), .B(n209), .Y(n210) );
  INVX1 U36 ( .A(n374), .Y(n53) );
  INVX1 U37 ( .A(n182), .Y(n57) );
  NOR2X1 U38 ( .A(n371), .B(n39), .Y(n325) );
  CLKINVX3 U39 ( .A(n391), .Y(n386) );
  NAND2X1 U40 ( .A(n371), .B(n71), .Y(n118) );
  NAND2X1 U41 ( .A(n56), .B(n371), .Y(n233) );
  NAND2X1 U42 ( .A(n138), .B(n371), .Y(n223) );
  NAND2X1 U43 ( .A(n39), .B(n371), .Y(n248) );
  NAND2X1 U44 ( .A(n181), .B(n371), .Y(n166) );
  NAND2X1 U45 ( .A(n229), .B(n248), .Y(n87) );
  INVX1 U46 ( .A(n102), .Y(n61) );
  NAND2X1 U47 ( .A(n115), .B(n223), .Y(n306) );
  INVX1 U48 ( .A(n168), .Y(n62) );
  INVX1 U49 ( .A(n230), .Y(n69) );
  INVX1 U50 ( .A(n116), .Y(n64) );
  INVX1 U51 ( .A(n103), .Y(n68) );
  BUFX3 U52 ( .A(n74), .Y(n371) );
  NAND2X1 U53 ( .A(n50), .B(n367), .Y(n147) );
  NAND2X1 U54 ( .A(n367), .B(n375), .Y(n120) );
  NAND2X1 U55 ( .A(n367), .B(n113), .Y(n165) );
  NAND2X1 U56 ( .A(n367), .B(n138), .Y(n182) );
  INVX1 U57 ( .A(n170), .Y(d[5]) );
  INVX1 U58 ( .A(n312), .Y(d[1]) );
  INVX1 U59 ( .A(n373), .Y(n46) );
  NAND2X1 U60 ( .A(n16), .B(n368), .Y(n259) );
  NAND2X1 U61 ( .A(n111), .B(n147), .Y(n96) );
  NOR2X1 U62 ( .A(n373), .B(n371), .Y(n124) );
  NAND2X1 U63 ( .A(n111), .B(n371), .Y(n268) );
  CLKINVX3 U64 ( .A(n111), .Y(n39) );
  NAND2X1 U65 ( .A(n367), .B(n71), .Y(n230) );
  NAND2X1 U66 ( .A(n367), .B(n66), .Y(n337) );
  NAND2BX1 U67 ( .AN(n124), .B(n263), .Y(n196) );
  INVX1 U68 ( .A(n156), .Y(n24) );
  NAND2X1 U69 ( .A(n224), .B(n268), .Y(n141) );
  NAND2BX1 U70 ( .AN(n93), .B(n373), .Y(n299) );
  NAND2X1 U71 ( .A(n224), .B(n233), .Y(n104) );
  NAND2X1 U72 ( .A(n263), .B(n142), .Y(n100) );
  CLKINVX3 U73 ( .A(n370), .Y(n21) );
  CLKINVX3 U74 ( .A(n108), .Y(n22) );
  INVX1 U76 ( .A(n249), .Y(d[3]) );
  BUFX3 U77 ( .A(a[1]), .Y(n367) );
  NAND2X1 U78 ( .A(a[7]), .B(a[2]), .Y(n94) );
  NAND2X1 U79 ( .A(n369), .B(a[0]), .Y(n108) );
  INVX1 U80 ( .A(n238), .Y(n15) );
  NAND2X1 U81 ( .A(n59), .B(n376), .Y(n114) );
  NAND2X1 U82 ( .A(n51), .B(n392), .Y(n238) );
  INVX1 U83 ( .A(n288), .Y(n14) );
  NOR2X1 U84 ( .A(n386), .B(n325), .Y(n199) );
  NOR2X1 U85 ( .A(n49), .B(n62), .Y(n247) );
  NAND2X1 U86 ( .A(n222), .B(n376), .Y(n162) );
  INVX1 U87 ( .A(n301), .Y(n49) );
  INVX1 U88 ( .A(n166), .Y(n60) );
  INVX1 U89 ( .A(n207), .Y(n48) );
  INVX1 U90 ( .A(n228), .Y(n51) );
  INVX4 U91 ( .A(n372), .Y(n392) );
  NOR2BX1 U92 ( .AN(n214), .B(n69), .Y(n88) );
  NOR2X1 U93 ( .A(n53), .B(n70), .Y(n326) );
  NOR2X1 U94 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U95 ( .A(n34), .B(n223), .Y(n183) );
  INVX1 U96 ( .A(n118), .Y(n70) );
  NAND2X1 U97 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U98 ( .A(n233), .Y(n55) );
  INVX1 U99 ( .A(n223), .Y(n59) );
  NOR2X1 U100 ( .A(n57), .B(n55), .Y(n197) );
  INVX1 U101 ( .A(n248), .Y(n37) );
  OAI221XL U102 ( .A0(n58), .A1(n381), .B0(n98), .B1(n94), .C0(n18), .Y(n347)
         );
  INVX1 U103 ( .A(n199), .Y(n18) );
  INVX1 U104 ( .A(n127), .Y(n35) );
  NOR2X1 U105 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U106 ( .A(n212), .Y(n41) );
  NOR2X1 U107 ( .A(n62), .B(n55), .Y(n145) );
  INVX1 U108 ( .A(n306), .Y(n58) );
  INVX1 U109 ( .A(n158), .Y(n42) );
  INVX1 U110 ( .A(n87), .Y(n38) );
  INVX1 U111 ( .A(n210), .Y(n44) );
  NAND2X1 U112 ( .A(n63), .B(n371), .Y(n243) );
  OAI22X1 U113 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U114 ( .A0(n61), .A1(n383), .B0(n392), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U115 ( .A0(n392), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U116 ( .A(n116), .B(n229), .Y(n244) );
  NOR2X1 U117 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U118 ( .A0(n378), .A1(n207), .B0(n381), .B1(n374), .Y(n242) );
  CLKINVX3 U119 ( .A(n113), .Y(n50) );
  NAND2X1 U120 ( .A(n214), .B(n142), .Y(n90) );
  CLKINVX3 U121 ( .A(n181), .Y(n63) );
  AOI22X1 U122 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U123 ( .A0(n98), .A1(n381), .B0(n30), .B1(n378), .C0(n99), .Y(n91)
         );
  OAI221XL U124 ( .A0(n42), .A1(n381), .B0(n51), .B1(n378), .C0(n95), .Y(n92)
         );
  INVX1 U125 ( .A(n104), .Y(n30) );
  NAND2X1 U126 ( .A(n392), .B(n96), .Y(n187) );
  NAND2X1 U127 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U128 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  OAI221XL U129 ( .A0(n46), .A1(n387), .B0(n63), .B1(n381), .C0(n200), .Y(n194) );
  OAI221XL U130 ( .A0(n372), .A1(n196), .B0(n197), .B1(n381), .C0(n198), .Y(
        n195) );
  AOI211X1 U131 ( .A0(n201), .A1(n392), .B0(n202), .C0(n203), .Y(n200) );
  AOI22X1 U132 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U133 ( .A0(n35), .A1(n381), .B0(n44), .B1(n379), .C0(n333), .Y(n332) );
  OAI211X1 U134 ( .A0(n326), .A1(n386), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U135 ( .A0(n35), .A1(n392), .B0(n39), .B1(n390), .Y(n333) );
  AOI22X1 U136 ( .A0(n384), .A1(n63), .B0(n247), .B1(n375), .Y(n334) );
  AOI21X1 U137 ( .A0(n115), .A1(n243), .B0(n386), .Y(n360) );
  INVX1 U138 ( .A(n120), .Y(n4) );
  AND2X2 U139 ( .A(n165), .B(n166), .Y(n129) );
  NAND2X1 U140 ( .A(n374), .B(n214), .Y(n126) );
  OAI21XL U141 ( .A0(n165), .A1(n386), .B0(n187), .Y(n266) );
  INVX1 U142 ( .A(n284), .Y(n10) );
  OAI31X1 U143 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U144 ( .A0(n377), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U145 ( .A(n147), .Y(n47) );
  OAI22X1 U146 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U147 ( .A0(n392), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U148 ( .A0(n11), .A1(n371), .B0(n27), .B1(n392), .C0(n307), .Y(n302) );
  OAI22X1 U149 ( .A0(n64), .A1(n378), .B0(n386), .B1(n306), .Y(n304) );
  AOI222X1 U150 ( .A0(n56), .A1(n376), .B0(n60), .B1(n390), .C0(n384), .C1(n71), .Y(n356) );
  AOI21X1 U151 ( .A0(n50), .A1(n16), .B0(n366), .Y(n365) );
  OAI221XL U152 ( .A0(n387), .A1(n87), .B0(n94), .B1(n104), .C0(n246), .Y(n235) );
  AOI2BB2X1 U153 ( .B0(n11), .B1(n371), .A0N(n372), .A1N(n247), .Y(n246) );
  CLKINVX8 U154 ( .A(n382), .Y(n381) );
  CLKINVX3 U155 ( .A(n377), .Y(n375) );
  NOR2X1 U156 ( .A(n381), .B(n371), .Y(n202) );
  AOI211X1 U157 ( .A0(n45), .A1(n376), .B0(n204), .C0(n205), .Y(n192) );
  INVX1 U158 ( .A(n209), .Y(n45) );
  NAND2BX1 U159 ( .AN(n97), .B(n206), .Y(n205) );
  AOI222X1 U160 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n376), 
        .Y(n198) );
  AOI221X1 U161 ( .A0(n321), .A1(n389), .B0(n376), .B1(n311), .C0(n327), .Y(
        n315) );
  OAI221XL U162 ( .A0(n372), .A1(n209), .B0(n381), .B1(n103), .C0(n288), .Y(
        n327) );
  AOI221X1 U163 ( .A0(n4), .A1(n71), .B0(n389), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI2BB1X1 U164 ( .A0N(n142), .A1N(n383), .B0(n187), .Y(n186) );
  OAI221XL U165 ( .A0(n308), .A1(n387), .B0(n381), .B1(n165), .C0(n162), .Y(
        n307) );
  NOR2X1 U166 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U167 ( .A0(n54), .A1(n381), .B0(n33), .B1(n378), .C0(n232), .Y(n217) );
  INVX1 U168 ( .A(n234), .Y(n54) );
  AOI32X1 U169 ( .A0(n34), .A1(n181), .A2(n392), .B0(n389), .B1(n233), .Y(n232) );
  OAI221XL U170 ( .A0(n67), .A1(n387), .B0(n94), .B1(n374), .C0(n294), .Y(n282) );
  INVX1 U171 ( .A(n115), .Y(n67) );
  AOI211X1 U172 ( .A0(n48), .A1(n392), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U173 ( .A(n114), .Y(n6) );
  AOI211X1 U174 ( .A0(n60), .A1(n376), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U175 ( .A(n381), .B(n39), .C(n61), .Y(n364) );
  INVX1 U176 ( .A(n259), .Y(n13) );
  OAI221XL U177 ( .A0(n372), .A1(n168), .B0(n164), .B1(n387), .C0(n169), .Y(
        n150) );
  AOI22X1 U178 ( .A0(n385), .A1(n34), .B0(n48), .B1(n375), .Y(n169) );
  AOI211X1 U179 ( .A0(n390), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  CLKINVX3 U180 ( .A(n391), .Y(n387) );
  INVX1 U181 ( .A(n125), .Y(n7) );
  AOI221X1 U182 ( .A0(n126), .A1(n388), .B0(n127), .B1(n385), .C0(n128), .Y(
        n125) );
  OAI21XL U183 ( .A0(n372), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U184 ( .A(n372), .Y(n16) );
  NOR2X1 U185 ( .A(n39), .B(n57), .Y(n179) );
  CLKINVX3 U186 ( .A(n110), .Y(n23) );
  NAND3X1 U187 ( .A(n374), .B(n113), .C(n376), .Y(n89) );
  NAND2X1 U188 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U189 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U190 ( .A(n374), .B(n166), .Y(n311) );
  NOR2BX1 U191 ( .AN(n229), .B(n68), .Y(n164) );
  AOI21X1 U192 ( .A0(n181), .A1(n182), .B0(n372), .Y(n180) );
  OAI221XL U193 ( .A0(n36), .A1(n386), .B0(n121), .B1(n379), .C0(n140), .Y(
        n135) );
  INVX1 U194 ( .A(n85), .Y(n36) );
  AOI22X1 U195 ( .A0(n49), .A1(n385), .B0(n392), .B1(n141), .Y(n140) );
  AOI22X1 U196 ( .A0(n57), .A1(n382), .B0(n391), .B1(n113), .Y(n239) );
  AOI22X1 U197 ( .A0(n383), .A1(n311), .B0(n50), .B1(n375), .Y(n350) );
  NOR2X1 U198 ( .A(n138), .B(n372), .Y(n97) );
  NAND2X1 U199 ( .A(n243), .B(n142), .Y(n127) );
  INVX1 U200 ( .A(n154), .Y(n25) );
  NAND2X1 U201 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U202 ( .A(n138), .Y(n56) );
  NAND2X1 U203 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U204 ( .A(n64), .B(n124), .Y(n121) );
  AOI211X1 U205 ( .A0(n392), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  OAI2BB2X1 U206 ( .B0(n381), .B1(n183), .A0N(n188), .A1N(n376), .Y(n335) );
  AOI21X1 U207 ( .A0(n301), .A1(n337), .B0(n386), .Y(n336) );
  NAND2X1 U208 ( .A(n138), .B(n102), .Y(n227) );
  NAND2X1 U209 ( .A(n103), .B(n165), .Y(n188) );
  AOI21X1 U210 ( .A0(n16), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U211 ( .A0(n102), .A1(n103), .B0(n386), .Y(n101) );
  INVX1 U212 ( .A(n337), .Y(n65) );
  AOI22X1 U213 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  OAI221XL U214 ( .A0(n65), .A1(n387), .B0(n31), .B1(n372), .C0(n149), .Y(n143) );
  OAI221XL U215 ( .A0(n145), .A1(n381), .B0(n28), .B1(n387), .C0(n146), .Y(
        n144) );
  AOI2BB2X1 U216 ( .B0(n375), .B1(n87), .A0N(n381), .A1N(n121), .Y(n149) );
  INVX1 U217 ( .A(n208), .Y(n29) );
  INVX1 U218 ( .A(n299), .Y(n11) );
  INVX1 U219 ( .A(n100), .Y(n33) );
  AOI221XL U220 ( .A0(n392), .A1(n52), .B0(n384), .B1(n123), .C0(n324), .Y(
        n316) );
  INVX1 U221 ( .A(n326), .Y(n52) );
  OAI32X1 U222 ( .A0(n94), .A1(n63), .A2(n325), .B0(n37), .B1(n387), .Y(n324)
         );
  INVX1 U223 ( .A(n196), .Y(n31) );
  OAI221XL U224 ( .A0(n56), .A1(n381), .B0(n32), .B1(n379), .C0(n163), .Y(n151) );
  INVX1 U225 ( .A(n167), .Y(n32) );
  AOI22X1 U226 ( .A0(n164), .A1(n16), .B0(n129), .B1(n390), .Y(n163) );
  INVX1 U227 ( .A(n141), .Y(n27) );
  INVX1 U228 ( .A(n148), .Y(n28) );
  OAI221XL U229 ( .A0(n40), .A1(n387), .B0(n58), .B1(n381), .C0(n137), .Y(n136) );
  INVX1 U230 ( .A(n96), .Y(n40) );
  AOI31X1 U231 ( .A0(n102), .A1(n138), .A2(n392), .B0(n8), .Y(n137) );
  INVX1 U232 ( .A(n89), .Y(n8) );
  INVX1 U233 ( .A(n185), .Y(n19) );
  INVX1 U234 ( .A(n380), .Y(n379) );
  INVX1 U235 ( .A(n375), .Y(n378) );
  OAI22X2 U236 ( .A0(n370), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  AOI211X1 U237 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U238 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI2BB2X1 U239 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  OAI22X2 U240 ( .A0(n370), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  AOI211X1 U241 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U242 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U243 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  OAI21X2 U244 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  OAI2BB1X1 U245 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI221X1 U246 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76)
         );
  AOI22X1 U247 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  AOI22X1 U248 ( .A0(n369), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U249 ( .A0(n61), .A1(n387), .B0(n381), .B1(n260), .C0(n261), .Y(
        n254) );
  OAI221XL U250 ( .A0(n41), .A1(n381), .B0(n378), .B1(n181), .C0(n256), .Y(
        n255) );
  AOI21X1 U251 ( .A0(n33), .A1(n392), .B0(n262), .Y(n261) );
  AOI22X1 U252 ( .A0(n348), .A1(n26), .B0(n369), .B1(n349), .Y(n342) );
  OAI221XL U253 ( .A0(n372), .A1(n166), .B0(n286), .B1(n381), .C0(n351), .Y(
        n348) );
  OAI211X1 U254 ( .A0(n88), .A1(n386), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U255 ( .B0(n375), .B1(n196), .A0N(n386), .A1N(n179), .Y(n351) );
  OAI22X1 U256 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U257 ( .A0(n385), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U258 ( .A0(n56), .A1(n4), .B0(n383), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U259 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U260 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U261 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U262 ( .A0(n61), .A1(n388), .B0(n383), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U263 ( .A0(n377), .A1(n71), .B0(n37), .B1(n386), .Y(n157) );
  OAI22X1 U264 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U265 ( .A0(n385), .A1(n111), .B0(n47), .B1(n376), .C0(n112), .Y(
        n109) );
  AOI221X1 U266 ( .A0(n392), .A1(n115), .B0(n388), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U267 ( .A0(n372), .A1(n113), .B0(n44), .B1(n387), .C0(n114), .Y(
        n112) );
  AOI211X1 U268 ( .A0(n55), .A1(n392), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U269 ( .A0(n114), .A1(n206), .A2(n273), .B0(n369), .Y(n272) );
  OAI22X1 U270 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U271 ( .B0(n70), .B1(n388), .A0N(n90), .A1N(n381), .Y(n273) );
  AOI2BB2X1 U272 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  OAI221XL U273 ( .A0(n46), .A1(n387), .B0(n381), .B1(n116), .C0(n267), .Y(
        n264) );
  AOI221XL U274 ( .A0(n384), .A1(n247), .B0(n212), .B1(n376), .C0(n266), .Y(
        n265) );
  AOI22X1 U275 ( .A0(n375), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  AOI22X1 U276 ( .A0(n370), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U277 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  OAI221XL U278 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  AOI22X1 U279 ( .A0(n171), .A1(n21), .B0(n370), .B1(n172), .Y(n170) );
  OAI221XL U281 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  OAI221XL U282 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  AOI22X1 U283 ( .A0(n388), .A1(n368), .B0(n375), .B1(n66), .Y(n292) );
  AOI22X1 U284 ( .A0(n369), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U285 ( .A0(n43), .A1(n381), .B0(n378), .B1(n34), .C0(n365), .Y(n361) );
  OAI221XL U286 ( .A0(n368), .A1(n120), .B0(n201), .B1(n387), .C0(n363), .Y(
        n362) );
  INVX1 U287 ( .A(n260), .Y(n43) );
  AOI22X1 U288 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  OAI21XL U289 ( .A0(n321), .A1(n372), .B0(n322), .Y(n318) );
  OAI221XL U290 ( .A0(n387), .A1(n113), .B0(n88), .B1(n381), .C0(n320), .Y(
        n319) );
  AOI31X1 U291 ( .A0(n374), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  CLKINVX3 U292 ( .A(n368), .Y(n71) );
  OAI21XL U293 ( .A0(n381), .A1(n373), .B0(n120), .Y(n276) );
  NAND2X1 U294 ( .A(n63), .B(n367), .Y(n168) );
  AOI21X1 U295 ( .A0(n224), .A1(n243), .B0(n381), .Y(n295) );
  INVX1 U296 ( .A(n367), .Y(n74) );
  OAI21XL U297 ( .A0(n73), .A1(n301), .B0(n386), .Y(n323) );
  OAI21XL U298 ( .A0(n73), .A1(n243), .B0(n386), .Y(n245) );
  OAI21XL U299 ( .A0(n372), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U300 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U301 ( .A(n162), .Y(n5) );
  AOI211X1 U302 ( .A0(n39), .A1(n376), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U303 ( .A0(n387), .A1(n116), .B0(n73), .B1(n230), .C0(n381), .C1(
        n102), .Y(n275) );
  NAND2X1 U304 ( .A(n62), .B(n390), .Y(n287) );
  OAI21X2 U305 ( .A0(n370), .A1(n131), .B0(n132), .Y(d[6]) );
  OAI2BB1X1 U306 ( .A0N(n133), .A1N(n134), .B0(n370), .Y(n132) );
  AOI221X1 U307 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131) );
  AOI22X1 U308 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  NOR2BX1 U309 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U310 ( .A(n82), .Y(n372) );
  NAND2X1 U311 ( .A(n73), .B(n20), .Y(n82) );
  OAI221XL U312 ( .A0(n367), .A1(n259), .B0(n379), .B1(n214), .C0(n287), .Y(
        n293) );
  BUFX3 U313 ( .A(n139), .Y(n374) );
  NAND2X1 U314 ( .A(n367), .B(n373), .Y(n139) );
  AOI211X1 U315 ( .A0(n376), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  OAI222X1 U316 ( .A0(n387), .A1(n167), .B0(n339), .B1(n372), .C0(n381), .C1(
        n34), .Y(n338) );
  AOI21X1 U317 ( .A0(n373), .A1(n371), .B0(n65), .Y(n339) );
  AOI211X1 U318 ( .A0(n369), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  OAI221XL U319 ( .A0(n381), .A1(n116), .B0(n321), .B1(n377), .C0(n359), .Y(
        n354) );
  AOI21X1 U320 ( .A0(n356), .A1(n357), .B0(n369), .Y(n355) );
  AOI31X1 U321 ( .A0(n392), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  INVX1 U322 ( .A(n93), .Y(n382) );
  INVX1 U323 ( .A(n83), .Y(n390) );
  INVX1 U324 ( .A(n83), .Y(n391) );
  INVX1 U325 ( .A(n380), .Y(n377) );
  INVX1 U326 ( .A(n94), .Y(n380) );
  AOI22X1 U327 ( .A0(n369), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U328 ( .A0(n381), .A1(n141), .B0(n387), .B1(n263), .C0(n29), .C1(
        n377), .Y(n277) );
  OAI221XL U329 ( .A0(n31), .A1(n372), .B0(n387), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U330 ( .B0(n88), .B1(n375), .A0N(n381), .A1N(n197), .Y(n279) );
  NAND2X1 U331 ( .A(n224), .B(n301), .Y(n148) );
  NOR2BX1 U332 ( .AN(n263), .B(n61), .Y(n321) );
  AOI21X1 U333 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI22X1 U334 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U335 ( .A0(n63), .A1(n381), .B0(n378), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U336 ( .A0(n38), .A1(n372), .B0(n381), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U337 ( .A0(n179), .A1(n388), .B0(n180), .Y(n178) );
  AOI22X1 U338 ( .A0(n392), .A1(n66), .B0(n375), .B1(n147), .Y(n146) );
  AOI22X1 U339 ( .A0(n384), .A1(n85), .B0(n41), .B1(n375), .Y(n84) );
  AOI31X1 U340 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U341 ( .A0N(n223), .A1N(n224), .B0(n389), .Y(n220) );
  AOI22X1 U342 ( .A0(n29), .A1(n392), .B0(n222), .B1(n383), .Y(n221) );
  NAND2X1 U343 ( .A(n224), .B(n118), .Y(n208) );
  NAND2X1 U344 ( .A(n263), .B(n337), .Y(n167) );
  AOI21X1 U345 ( .A0(n263), .A1(n182), .B0(n381), .Y(n305) );
  AOI21X1 U346 ( .A0(n111), .A1(n374), .B0(n377), .Y(n203) );
  NAND2X1 U347 ( .A(n16), .B(n367), .Y(n206) );
  XNOR2X1 U348 ( .A(n20), .B(n367), .Y(n185) );
  NAND2X1 U349 ( .A(n375), .B(n373), .Y(n130) );
  XNOR2X1 U350 ( .A(n73), .B(n367), .Y(n161) );
  AOI21X1 U351 ( .A0(n90), .A1(n73), .B0(n392), .Y(n86) );
  AOI221X1 U352 ( .A0(n46), .A1(n376), .B0(n389), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U353 ( .A0(n372), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U354 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  AOI222X1 U355 ( .A0(n385), .A1(n210), .B0(n211), .B1(n212), .C0(n392), .C1(
        n373), .Y(n191) );
  OAI21XL U356 ( .A0(n73), .A1(n214), .B0(n386), .Y(n211) );
  AOI31X1 U357 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U358 ( .A0(n148), .A1(n73), .B0(n29), .B1(n389), .Y(n300) );
  INVX1 U359 ( .A(n93), .Y(n383) );
  INVX1 U360 ( .A(n93), .Y(n385) );
  INVX1 U361 ( .A(n93), .Y(n384) );
  XOR2X1 U362 ( .A(n369), .B(n367), .Y(n358) );
  INVX1 U363 ( .A(n83), .Y(n388) );
  INVX1 U364 ( .A(n83), .Y(n389) );
  NOR2BX1 U365 ( .AN(n93), .B(n390), .Y(n309) );
  OAI22X2 U366 ( .A0(n340), .A1(n21), .B0(n370), .B1(n341), .Y(d[0]) );
  AOI22X1 U367 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U368 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI22X1 U369 ( .A0(n347), .A1(n26), .B0(n392), .B1(n90), .Y(n343) );
  AOI22X1 U370 ( .A0(n250), .A1(n21), .B0(n370), .B1(n251), .Y(n249) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  OAI22X1 U373 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U374 ( .A0(n384), .A1(n230), .B0(n392), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U375 ( .A0(n164), .A1(n383), .B0(a[2]), .B1(n227), .C0(n392), .C1(
        n228), .Y(n226) );
  OAI22X1 U376 ( .A0(n35), .A1(n379), .B0(n386), .B1(n373), .Y(n231) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n373) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI21XL U383 ( .A0(n66), .A1(n386), .B0(n259), .Y(n257) );
  BUFX3 U384 ( .A(a[3]), .Y(n368) );
  AOI22X1 U385 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U386 ( .A(a[0]), .Y(n75) );
  AOI211X1 U387 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U388 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U389 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U390 ( .A(a[5]), .Y(n369) );
  OAI221XL U391 ( .A0(n372), .A1(n115), .B0(n121), .B1(n381), .C0(n122), .Y(
        n105) );
  AOI22X1 U392 ( .A0(n375), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  AOI33X1 U393 ( .A0(n368), .A1(n376), .A2(n19), .B0(n185), .B1(n181), .B2(
        a[2]), .Y(n184) );
  BUFX3 U394 ( .A(a[6]), .Y(n370) );
endmodule


module aes_sbox_19 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556;

  OAI221X4 U4 ( .A0(n66), .A1(n536), .B0(n61), .B1(n551), .C0(n84), .Y(n81) );
  OAI221X4 U6 ( .A0(n86), .A1(n87), .B0(n88), .B1(n551), .C0(n89), .Y(n80) );
  OAI222X4 U75 ( .A0(n551), .A1(n207), .B0(n181), .B1(n120), .C0(n545), .C1(
        n208), .Y(n204) );
  OAI32X4 U280 ( .A0(n551), .A1(n56), .A2(n53), .B0(n94), .B1(n103), .Y(n366)
         );
  AOI221X1 U1 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n56), .B(n531), .Y(n229) );
  NAND2X2 U5 ( .A(n532), .B(n66), .Y(n181) );
  NAND2X1 U7 ( .A(n39), .B(n531), .Y(n142) );
  NAND2X2 U8 ( .A(n66), .B(n71), .Y(n138) );
  NAND2X1 U9 ( .A(n532), .B(n535), .Y(n103) );
  NAND2X1 U10 ( .A(n531), .B(n181), .Y(n102) );
  NAND2X2 U11 ( .A(n537), .B(n181), .Y(n113) );
  OAI222X1 U12 ( .A0(n94), .A1(n118), .B0(n119), .B1(n545), .C0(a[4]), .C1(
        n120), .Y(n117) );
  NAND2X2 U13 ( .A(n66), .B(n535), .Y(n116) );
  NAND2X2 U14 ( .A(n531), .B(n532), .Y(n115) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n73) );
  NAND2X1 U16 ( .A(n533), .B(n75), .Y(n110) );
  CLKINVX3 U17 ( .A(n533), .Y(n26) );
  NAND2X2 U18 ( .A(a[0]), .B(n26), .Y(n156) );
  NAND2X2 U19 ( .A(n75), .B(n26), .Y(n154) );
  NAND2X1 U20 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U21 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI21XL U22 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  NAND2X1 U23 ( .A(a[4]), .B(n535), .Y(n263) );
  NAND2X1 U24 ( .A(n531), .B(a[4]), .Y(n224) );
  NAND2X2 U25 ( .A(n532), .B(a[4]), .Y(n111) );
  CLKINVX3 U26 ( .A(a[4]), .Y(n66) );
  NAND2X1 U27 ( .A(n53), .B(n556), .Y(n288) );
  CLKINVX3 U28 ( .A(n543), .Y(n540) );
  INVX1 U29 ( .A(n325), .Y(n34) );
  NAND2X1 U30 ( .A(n113), .B(n535), .Y(n214) );
  NAND2X1 U31 ( .A(n46), .B(n535), .Y(n209) );
  NAND2X1 U32 ( .A(n50), .B(n535), .Y(n301) );
  NAND2X1 U33 ( .A(n538), .B(n268), .Y(n212) );
  NAND2X1 U34 ( .A(n147), .B(n214), .Y(n207) );
  NAND2X1 U35 ( .A(n115), .B(n209), .Y(n210) );
  INVX1 U36 ( .A(n538), .Y(n53) );
  INVX1 U37 ( .A(n182), .Y(n57) );
  NOR2X1 U38 ( .A(n535), .B(n39), .Y(n325) );
  CLKINVX3 U39 ( .A(n555), .Y(n550) );
  NAND2X1 U40 ( .A(n535), .B(n71), .Y(n118) );
  NAND2X1 U41 ( .A(n56), .B(n535), .Y(n233) );
  NAND2X1 U42 ( .A(n138), .B(n535), .Y(n223) );
  NAND2X1 U43 ( .A(n39), .B(n535), .Y(n248) );
  NAND2X1 U44 ( .A(n181), .B(n535), .Y(n166) );
  NAND2X1 U45 ( .A(n229), .B(n248), .Y(n87) );
  INVX1 U46 ( .A(n102), .Y(n61) );
  NAND2X1 U47 ( .A(n115), .B(n223), .Y(n306) );
  INVX1 U48 ( .A(n168), .Y(n62) );
  INVX1 U49 ( .A(n230), .Y(n69) );
  INVX1 U50 ( .A(n116), .Y(n64) );
  INVX1 U51 ( .A(n103), .Y(n68) );
  BUFX3 U52 ( .A(n74), .Y(n535) );
  NAND2X1 U53 ( .A(n50), .B(n531), .Y(n147) );
  NAND2X1 U54 ( .A(n531), .B(n539), .Y(n120) );
  NAND2X1 U55 ( .A(n531), .B(n113), .Y(n165) );
  NAND2X1 U56 ( .A(n531), .B(n138), .Y(n182) );
  INVX1 U57 ( .A(n170), .Y(d[5]) );
  INVX1 U58 ( .A(n312), .Y(d[1]) );
  INVX1 U59 ( .A(n537), .Y(n46) );
  NAND2X1 U60 ( .A(n16), .B(n532), .Y(n259) );
  NAND2X1 U61 ( .A(n111), .B(n147), .Y(n96) );
  NOR2X1 U62 ( .A(n537), .B(n535), .Y(n124) );
  NAND2X1 U63 ( .A(n111), .B(n535), .Y(n268) );
  CLKINVX3 U64 ( .A(n111), .Y(n39) );
  NAND2X1 U65 ( .A(n531), .B(n71), .Y(n230) );
  NAND2X1 U66 ( .A(n531), .B(n66), .Y(n337) );
  NAND2BX1 U67 ( .AN(n124), .B(n263), .Y(n196) );
  INVX1 U68 ( .A(n156), .Y(n24) );
  NAND2X1 U69 ( .A(n224), .B(n268), .Y(n141) );
  NAND2BX1 U70 ( .AN(n93), .B(n537), .Y(n299) );
  NAND2X1 U71 ( .A(n224), .B(n233), .Y(n104) );
  NAND2X1 U72 ( .A(n263), .B(n142), .Y(n100) );
  CLKINVX3 U73 ( .A(n534), .Y(n21) );
  CLKINVX3 U74 ( .A(n108), .Y(n22) );
  INVX1 U76 ( .A(n249), .Y(d[3]) );
  BUFX3 U77 ( .A(a[1]), .Y(n531) );
  NAND2X1 U78 ( .A(a[7]), .B(a[2]), .Y(n94) );
  NAND2X1 U79 ( .A(n533), .B(a[0]), .Y(n108) );
  INVX1 U80 ( .A(n238), .Y(n15) );
  NAND2X1 U81 ( .A(n59), .B(n540), .Y(n114) );
  NAND2X1 U82 ( .A(n51), .B(n556), .Y(n238) );
  INVX1 U83 ( .A(n288), .Y(n14) );
  NOR2X1 U84 ( .A(n550), .B(n325), .Y(n199) );
  NOR2X1 U85 ( .A(n49), .B(n62), .Y(n247) );
  NAND2X1 U86 ( .A(n222), .B(n540), .Y(n162) );
  INVX1 U87 ( .A(n301), .Y(n49) );
  INVX1 U88 ( .A(n166), .Y(n60) );
  INVX1 U89 ( .A(n207), .Y(n48) );
  INVX1 U90 ( .A(n228), .Y(n51) );
  INVX4 U91 ( .A(n536), .Y(n556) );
  NOR2BX1 U92 ( .AN(n214), .B(n69), .Y(n88) );
  NOR2X1 U93 ( .A(n53), .B(n70), .Y(n326) );
  NOR2X1 U94 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U95 ( .A(n34), .B(n223), .Y(n183) );
  INVX1 U96 ( .A(n118), .Y(n70) );
  NAND2X1 U97 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U98 ( .A(n233), .Y(n55) );
  INVX1 U99 ( .A(n223), .Y(n59) );
  NOR2X1 U100 ( .A(n57), .B(n55), .Y(n197) );
  INVX1 U101 ( .A(n248), .Y(n37) );
  OAI221XL U102 ( .A0(n58), .A1(n545), .B0(n98), .B1(n94), .C0(n18), .Y(n347)
         );
  INVX1 U103 ( .A(n199), .Y(n18) );
  INVX1 U104 ( .A(n127), .Y(n35) );
  NOR2X1 U105 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U106 ( .A(n212), .Y(n41) );
  NOR2X1 U107 ( .A(n62), .B(n55), .Y(n145) );
  INVX1 U108 ( .A(n306), .Y(n58) );
  INVX1 U109 ( .A(n158), .Y(n42) );
  INVX1 U110 ( .A(n87), .Y(n38) );
  INVX1 U111 ( .A(n210), .Y(n44) );
  NAND2X1 U112 ( .A(n63), .B(n535), .Y(n243) );
  OAI22X1 U113 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U114 ( .A0(n61), .A1(n547), .B0(n556), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U115 ( .A0(n556), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U116 ( .A(n116), .B(n229), .Y(n244) );
  NOR2X1 U117 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U118 ( .A0(n542), .A1(n207), .B0(n545), .B1(n538), .Y(n242) );
  CLKINVX3 U119 ( .A(n113), .Y(n50) );
  NAND2X1 U120 ( .A(n214), .B(n142), .Y(n90) );
  CLKINVX3 U121 ( .A(n181), .Y(n63) );
  AOI22X1 U122 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U123 ( .A0(n98), .A1(n545), .B0(n30), .B1(n542), .C0(n99), .Y(n91)
         );
  OAI221XL U124 ( .A0(n42), .A1(n545), .B0(n51), .B1(n542), .C0(n95), .Y(n92)
         );
  INVX1 U125 ( .A(n104), .Y(n30) );
  NAND2X1 U126 ( .A(n556), .B(n96), .Y(n187) );
  NAND2X1 U127 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U128 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  OAI221XL U129 ( .A0(n46), .A1(n551), .B0(n63), .B1(n545), .C0(n200), .Y(n194) );
  OAI221XL U130 ( .A0(n536), .A1(n196), .B0(n197), .B1(n545), .C0(n198), .Y(
        n195) );
  AOI211X1 U131 ( .A0(n201), .A1(n556), .B0(n202), .C0(n203), .Y(n200) );
  AOI22X1 U132 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U133 ( .A0(n35), .A1(n545), .B0(n44), .B1(n543), .C0(n333), .Y(n332) );
  OAI211X1 U134 ( .A0(n326), .A1(n550), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U135 ( .A0(n35), .A1(n556), .B0(n39), .B1(n554), .Y(n333) );
  AOI22X1 U136 ( .A0(n548), .A1(n63), .B0(n247), .B1(n539), .Y(n334) );
  AOI21X1 U137 ( .A0(n115), .A1(n243), .B0(n550), .Y(n360) );
  INVX1 U138 ( .A(n120), .Y(n4) );
  AND2X2 U139 ( .A(n165), .B(n166), .Y(n129) );
  NAND2X1 U140 ( .A(n538), .B(n214), .Y(n126) );
  OAI21XL U141 ( .A0(n165), .A1(n550), .B0(n187), .Y(n266) );
  INVX1 U142 ( .A(n284), .Y(n10) );
  OAI31X1 U143 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U144 ( .A0(n541), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U145 ( .A(n147), .Y(n47) );
  OAI22X1 U146 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U147 ( .A0(n556), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U148 ( .A0(n11), .A1(n535), .B0(n27), .B1(n556), .C0(n307), .Y(n302) );
  OAI22X1 U149 ( .A0(n64), .A1(n542), .B0(n550), .B1(n306), .Y(n304) );
  AOI222X1 U150 ( .A0(n56), .A1(n540), .B0(n60), .B1(n554), .C0(n548), .C1(n71), .Y(n356) );
  AOI21X1 U151 ( .A0(n50), .A1(n16), .B0(n366), .Y(n365) );
  OAI221XL U152 ( .A0(n551), .A1(n87), .B0(n94), .B1(n104), .C0(n246), .Y(n235) );
  AOI2BB2X1 U153 ( .B0(n11), .B1(n535), .A0N(n536), .A1N(n247), .Y(n246) );
  CLKINVX8 U154 ( .A(n546), .Y(n545) );
  CLKINVX3 U155 ( .A(n541), .Y(n539) );
  NOR2X1 U156 ( .A(n545), .B(n535), .Y(n202) );
  AOI211X1 U157 ( .A0(n45), .A1(n540), .B0(n204), .C0(n205), .Y(n192) );
  INVX1 U158 ( .A(n209), .Y(n45) );
  NAND2BX1 U159 ( .AN(n97), .B(n206), .Y(n205) );
  AOI222X1 U160 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n540), 
        .Y(n198) );
  AOI221X1 U161 ( .A0(n321), .A1(n553), .B0(n540), .B1(n311), .C0(n327), .Y(
        n315) );
  OAI221XL U162 ( .A0(n536), .A1(n209), .B0(n545), .B1(n103), .C0(n288), .Y(
        n327) );
  AOI221X1 U163 ( .A0(n4), .A1(n71), .B0(n553), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI2BB1X1 U164 ( .A0N(n142), .A1N(n547), .B0(n187), .Y(n186) );
  OAI221XL U165 ( .A0(n308), .A1(n551), .B0(n545), .B1(n165), .C0(n162), .Y(
        n307) );
  NOR2X1 U166 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U167 ( .A0(n54), .A1(n545), .B0(n33), .B1(n542), .C0(n232), .Y(n217) );
  INVX1 U168 ( .A(n234), .Y(n54) );
  AOI32X1 U169 ( .A0(n34), .A1(n181), .A2(n556), .B0(n553), .B1(n233), .Y(n232) );
  OAI221XL U170 ( .A0(n67), .A1(n551), .B0(n94), .B1(n538), .C0(n294), .Y(n282) );
  INVX1 U171 ( .A(n115), .Y(n67) );
  AOI211X1 U172 ( .A0(n48), .A1(n556), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U173 ( .A(n114), .Y(n6) );
  AOI211X1 U174 ( .A0(n60), .A1(n540), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U175 ( .A(n545), .B(n39), .C(n61), .Y(n364) );
  INVX1 U176 ( .A(n259), .Y(n13) );
  OAI221XL U177 ( .A0(n536), .A1(n168), .B0(n164), .B1(n551), .C0(n169), .Y(
        n150) );
  AOI22X1 U178 ( .A0(n549), .A1(n34), .B0(n48), .B1(n539), .Y(n169) );
  AOI211X1 U179 ( .A0(n554), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  CLKINVX3 U180 ( .A(n555), .Y(n551) );
  INVX1 U181 ( .A(n125), .Y(n7) );
  AOI221X1 U182 ( .A0(n126), .A1(n552), .B0(n127), .B1(n549), .C0(n128), .Y(
        n125) );
  OAI21XL U183 ( .A0(n536), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U184 ( .A(n536), .Y(n16) );
  NOR2X1 U185 ( .A(n39), .B(n57), .Y(n179) );
  CLKINVX3 U186 ( .A(n110), .Y(n23) );
  NAND3X1 U187 ( .A(n538), .B(n113), .C(n540), .Y(n89) );
  NAND2X1 U188 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U189 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U190 ( .A(n538), .B(n166), .Y(n311) );
  NOR2BX1 U191 ( .AN(n229), .B(n68), .Y(n164) );
  AOI21X1 U192 ( .A0(n181), .A1(n182), .B0(n536), .Y(n180) );
  OAI221XL U193 ( .A0(n36), .A1(n550), .B0(n121), .B1(n543), .C0(n140), .Y(
        n135) );
  INVX1 U194 ( .A(n85), .Y(n36) );
  AOI22X1 U195 ( .A0(n49), .A1(n549), .B0(n556), .B1(n141), .Y(n140) );
  AOI22X1 U196 ( .A0(n57), .A1(n546), .B0(n555), .B1(n113), .Y(n239) );
  AOI22X1 U197 ( .A0(n547), .A1(n311), .B0(n50), .B1(n539), .Y(n350) );
  NOR2X1 U198 ( .A(n138), .B(n536), .Y(n97) );
  NAND2X1 U199 ( .A(n243), .B(n142), .Y(n127) );
  INVX1 U200 ( .A(n154), .Y(n25) );
  NAND2X1 U201 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U202 ( .A(n138), .Y(n56) );
  NAND2X1 U203 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U204 ( .A(n64), .B(n124), .Y(n121) );
  AOI211X1 U205 ( .A0(n556), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  OAI2BB2X1 U206 ( .B0(n545), .B1(n183), .A0N(n188), .A1N(n540), .Y(n335) );
  AOI21X1 U207 ( .A0(n301), .A1(n337), .B0(n550), .Y(n336) );
  NAND2X1 U208 ( .A(n138), .B(n102), .Y(n227) );
  NAND2X1 U209 ( .A(n103), .B(n165), .Y(n188) );
  AOI21X1 U210 ( .A0(n16), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U211 ( .A0(n102), .A1(n103), .B0(n550), .Y(n101) );
  INVX1 U212 ( .A(n337), .Y(n65) );
  AOI22X1 U213 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  OAI221XL U214 ( .A0(n65), .A1(n551), .B0(n31), .B1(n536), .C0(n149), .Y(n143) );
  OAI221XL U215 ( .A0(n145), .A1(n545), .B0(n28), .B1(n551), .C0(n146), .Y(
        n144) );
  AOI2BB2X1 U216 ( .B0(n539), .B1(n87), .A0N(n545), .A1N(n121), .Y(n149) );
  INVX1 U217 ( .A(n208), .Y(n29) );
  INVX1 U218 ( .A(n299), .Y(n11) );
  INVX1 U219 ( .A(n100), .Y(n33) );
  AOI221XL U220 ( .A0(n556), .A1(n52), .B0(n548), .B1(n123), .C0(n324), .Y(
        n316) );
  INVX1 U221 ( .A(n326), .Y(n52) );
  OAI32X1 U222 ( .A0(n94), .A1(n63), .A2(n325), .B0(n37), .B1(n551), .Y(n324)
         );
  INVX1 U223 ( .A(n196), .Y(n31) );
  OAI221XL U224 ( .A0(n56), .A1(n545), .B0(n32), .B1(n543), .C0(n163), .Y(n151) );
  INVX1 U225 ( .A(n167), .Y(n32) );
  AOI22X1 U226 ( .A0(n164), .A1(n16), .B0(n129), .B1(n554), .Y(n163) );
  INVX1 U227 ( .A(n141), .Y(n27) );
  INVX1 U228 ( .A(n148), .Y(n28) );
  OAI221XL U229 ( .A0(n40), .A1(n551), .B0(n58), .B1(n545), .C0(n137), .Y(n136) );
  INVX1 U230 ( .A(n96), .Y(n40) );
  AOI31X1 U231 ( .A0(n102), .A1(n138), .A2(n556), .B0(n8), .Y(n137) );
  INVX1 U232 ( .A(n89), .Y(n8) );
  INVX1 U233 ( .A(n185), .Y(n19) );
  INVX1 U234 ( .A(n544), .Y(n543) );
  INVX1 U235 ( .A(n539), .Y(n542) );
  OAI22X2 U236 ( .A0(n534), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  AOI211X1 U237 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U238 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI2BB2X1 U239 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  OAI22X2 U240 ( .A0(n534), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  AOI211X1 U241 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U242 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U243 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  OAI21X2 U244 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  OAI2BB1X1 U245 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI221X1 U246 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76)
         );
  AOI22X1 U247 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  AOI22X1 U248 ( .A0(n533), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U249 ( .A0(n61), .A1(n551), .B0(n545), .B1(n260), .C0(n261), .Y(
        n254) );
  OAI221XL U250 ( .A0(n41), .A1(n545), .B0(n542), .B1(n181), .C0(n256), .Y(
        n255) );
  AOI21X1 U251 ( .A0(n33), .A1(n556), .B0(n262), .Y(n261) );
  AOI22X1 U252 ( .A0(n348), .A1(n26), .B0(n533), .B1(n349), .Y(n342) );
  OAI221XL U253 ( .A0(n536), .A1(n166), .B0(n286), .B1(n545), .C0(n351), .Y(
        n348) );
  OAI211X1 U254 ( .A0(n88), .A1(n550), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U255 ( .B0(n539), .B1(n196), .A0N(n550), .A1N(n179), .Y(n351) );
  OAI22X1 U256 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U257 ( .A0(n549), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U258 ( .A0(n56), .A1(n4), .B0(n547), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U259 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U260 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U261 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U262 ( .A0(n61), .A1(n552), .B0(n547), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U263 ( .A0(n541), .A1(n71), .B0(n37), .B1(n550), .Y(n157) );
  OAI22X1 U264 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U265 ( .A0(n549), .A1(n111), .B0(n47), .B1(n540), .C0(n112), .Y(
        n109) );
  AOI221X1 U266 ( .A0(n556), .A1(n115), .B0(n552), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U267 ( .A0(n536), .A1(n113), .B0(n44), .B1(n551), .C0(n114), .Y(
        n112) );
  AOI211X1 U268 ( .A0(n55), .A1(n556), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U269 ( .A0(n114), .A1(n206), .A2(n273), .B0(n533), .Y(n272) );
  OAI22X1 U270 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U271 ( .B0(n70), .B1(n552), .A0N(n90), .A1N(n545), .Y(n273) );
  AOI2BB2X1 U272 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  OAI221XL U273 ( .A0(n46), .A1(n551), .B0(n545), .B1(n116), .C0(n267), .Y(
        n264) );
  AOI221XL U274 ( .A0(n548), .A1(n247), .B0(n212), .B1(n540), .C0(n266), .Y(
        n265) );
  AOI22X1 U275 ( .A0(n539), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  AOI22X1 U276 ( .A0(n534), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U277 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  OAI221XL U278 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  AOI22X1 U279 ( .A0(n171), .A1(n21), .B0(n534), .B1(n172), .Y(n170) );
  OAI221XL U281 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  OAI221XL U282 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  AOI22X1 U283 ( .A0(n552), .A1(n532), .B0(n539), .B1(n66), .Y(n292) );
  AOI22X1 U284 ( .A0(n533), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U285 ( .A0(n43), .A1(n545), .B0(n542), .B1(n34), .C0(n365), .Y(n361) );
  OAI221XL U286 ( .A0(n532), .A1(n120), .B0(n201), .B1(n551), .C0(n363), .Y(
        n362) );
  INVX1 U287 ( .A(n260), .Y(n43) );
  AOI22X1 U288 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  OAI21XL U289 ( .A0(n321), .A1(n536), .B0(n322), .Y(n318) );
  OAI221XL U290 ( .A0(n551), .A1(n113), .B0(n88), .B1(n545), .C0(n320), .Y(
        n319) );
  AOI31X1 U291 ( .A0(n538), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  CLKINVX3 U292 ( .A(n532), .Y(n71) );
  OAI21XL U293 ( .A0(n545), .A1(n537), .B0(n120), .Y(n276) );
  NAND2X1 U294 ( .A(n63), .B(n531), .Y(n168) );
  AOI21X1 U295 ( .A0(n224), .A1(n243), .B0(n545), .Y(n295) );
  INVX1 U296 ( .A(n531), .Y(n74) );
  OAI21XL U297 ( .A0(n73), .A1(n301), .B0(n550), .Y(n323) );
  OAI21XL U298 ( .A0(n73), .A1(n243), .B0(n550), .Y(n245) );
  OAI21XL U299 ( .A0(n536), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U300 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U301 ( .A(n162), .Y(n5) );
  AOI211X1 U302 ( .A0(n39), .A1(n540), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U303 ( .A0(n551), .A1(n116), .B0(n73), .B1(n230), .C0(n545), .C1(
        n102), .Y(n275) );
  NAND2X1 U304 ( .A(n62), .B(n554), .Y(n287) );
  OAI21X2 U305 ( .A0(n534), .A1(n131), .B0(n132), .Y(d[6]) );
  OAI2BB1X1 U306 ( .A0N(n133), .A1N(n134), .B0(n534), .Y(n132) );
  AOI221X1 U307 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131) );
  AOI22X1 U308 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  NOR2BX1 U309 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U310 ( .A(n82), .Y(n536) );
  NAND2X1 U311 ( .A(n73), .B(n20), .Y(n82) );
  OAI221XL U312 ( .A0(n531), .A1(n259), .B0(n543), .B1(n214), .C0(n287), .Y(
        n293) );
  BUFX3 U313 ( .A(n139), .Y(n538) );
  NAND2X1 U314 ( .A(n531), .B(n537), .Y(n139) );
  AOI211X1 U315 ( .A0(n540), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  OAI222X1 U316 ( .A0(n551), .A1(n167), .B0(n339), .B1(n536), .C0(n545), .C1(
        n34), .Y(n338) );
  AOI21X1 U317 ( .A0(n537), .A1(n535), .B0(n65), .Y(n339) );
  AOI211X1 U318 ( .A0(n533), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  OAI221XL U319 ( .A0(n545), .A1(n116), .B0(n321), .B1(n541), .C0(n359), .Y(
        n354) );
  AOI21X1 U320 ( .A0(n356), .A1(n357), .B0(n533), .Y(n355) );
  AOI31X1 U321 ( .A0(n556), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  INVX1 U322 ( .A(n93), .Y(n546) );
  INVX1 U323 ( .A(n83), .Y(n554) );
  INVX1 U324 ( .A(n83), .Y(n555) );
  INVX1 U325 ( .A(n544), .Y(n541) );
  INVX1 U326 ( .A(n94), .Y(n544) );
  AOI22X1 U327 ( .A0(n533), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U328 ( .A0(n545), .A1(n141), .B0(n551), .B1(n263), .C0(n29), .C1(
        n541), .Y(n277) );
  OAI221XL U329 ( .A0(n31), .A1(n536), .B0(n551), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U330 ( .B0(n88), .B1(n539), .A0N(n545), .A1N(n197), .Y(n279) );
  NAND2X1 U331 ( .A(n224), .B(n301), .Y(n148) );
  NOR2BX1 U332 ( .AN(n263), .B(n61), .Y(n321) );
  AOI21X1 U333 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI22X1 U334 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U335 ( .A0(n63), .A1(n545), .B0(n542), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U336 ( .A0(n38), .A1(n536), .B0(n545), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U337 ( .A0(n179), .A1(n552), .B0(n180), .Y(n178) );
  AOI22X1 U338 ( .A0(n556), .A1(n66), .B0(n539), .B1(n147), .Y(n146) );
  AOI22X1 U339 ( .A0(n548), .A1(n85), .B0(n41), .B1(n539), .Y(n84) );
  AOI31X1 U340 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U341 ( .A0N(n223), .A1N(n224), .B0(n553), .Y(n220) );
  AOI22X1 U342 ( .A0(n29), .A1(n556), .B0(n222), .B1(n547), .Y(n221) );
  NAND2X1 U343 ( .A(n224), .B(n118), .Y(n208) );
  NAND2X1 U344 ( .A(n263), .B(n337), .Y(n167) );
  AOI21X1 U345 ( .A0(n263), .A1(n182), .B0(n545), .Y(n305) );
  AOI21X1 U346 ( .A0(n111), .A1(n538), .B0(n541), .Y(n203) );
  NAND2X1 U347 ( .A(n16), .B(n531), .Y(n206) );
  XNOR2X1 U348 ( .A(n20), .B(n531), .Y(n185) );
  NAND2X1 U349 ( .A(n539), .B(n537), .Y(n130) );
  XNOR2X1 U350 ( .A(n73), .B(n531), .Y(n161) );
  AOI21X1 U351 ( .A0(n90), .A1(n73), .B0(n556), .Y(n86) );
  AOI221X1 U352 ( .A0(n46), .A1(n540), .B0(n553), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U353 ( .A0(n536), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U354 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  AOI222X1 U355 ( .A0(n549), .A1(n210), .B0(n211), .B1(n212), .C0(n556), .C1(
        n537), .Y(n191) );
  OAI21XL U356 ( .A0(n73), .A1(n214), .B0(n550), .Y(n211) );
  AOI31X1 U357 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U358 ( .A0(n148), .A1(n73), .B0(n29), .B1(n553), .Y(n300) );
  INVX1 U359 ( .A(n93), .Y(n547) );
  INVX1 U360 ( .A(n93), .Y(n549) );
  INVX1 U361 ( .A(n93), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n358) );
  INVX1 U363 ( .A(n83), .Y(n552) );
  INVX1 U364 ( .A(n83), .Y(n553) );
  NOR2BX1 U365 ( .AN(n93), .B(n554), .Y(n309) );
  OAI22X2 U366 ( .A0(n340), .A1(n21), .B0(n534), .B1(n341), .Y(d[0]) );
  AOI22X1 U367 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U368 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI22X1 U369 ( .A0(n347), .A1(n26), .B0(n556), .B1(n90), .Y(n343) );
  AOI22X1 U370 ( .A0(n250), .A1(n21), .B0(n534), .B1(n251), .Y(n249) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  OAI22X1 U373 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U374 ( .A0(n548), .A1(n230), .B0(n556), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U375 ( .A0(n164), .A1(n547), .B0(a[2]), .B1(n227), .C0(n556), .C1(
        n228), .Y(n226) );
  OAI22X1 U376 ( .A0(n35), .A1(n543), .B0(n550), .B1(n537), .Y(n231) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI21XL U383 ( .A0(n66), .A1(n550), .B0(n259), .Y(n257) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI22X1 U385 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U386 ( .A(a[0]), .Y(n75) );
  AOI211X1 U387 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U388 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U389 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U390 ( .A(a[5]), .Y(n533) );
  OAI221XL U391 ( .A0(n536), .A1(n115), .B0(n121), .B1(n545), .C0(n122), .Y(
        n105) );
  AOI22X1 U392 ( .A0(n539), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  AOI33X1 U393 ( .A0(n532), .A1(n540), .A2(n19), .B0(n185), .B1(n181), .B2(
        a[2]), .Y(n184) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_18 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556;

  OAI221X4 U4 ( .A0(n66), .A1(n536), .B0(n61), .B1(n551), .C0(n84), .Y(n81) );
  OAI221X4 U6 ( .A0(n86), .A1(n87), .B0(n88), .B1(n551), .C0(n89), .Y(n80) );
  OAI222X4 U75 ( .A0(n551), .A1(n207), .B0(n181), .B1(n120), .C0(n545), .C1(
        n208), .Y(n204) );
  OAI32X4 U280 ( .A0(n551), .A1(n56), .A2(n53), .B0(n94), .B1(n103), .Y(n366)
         );
  AOI221X1 U1 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n56), .B(n531), .Y(n229) );
  NAND2X2 U5 ( .A(n532), .B(n66), .Y(n181) );
  NAND2X1 U7 ( .A(n39), .B(n531), .Y(n142) );
  NAND2X2 U8 ( .A(n66), .B(n71), .Y(n138) );
  NAND2X1 U9 ( .A(n532), .B(n535), .Y(n103) );
  NAND2X1 U10 ( .A(n531), .B(n181), .Y(n102) );
  NAND2X2 U11 ( .A(n537), .B(n181), .Y(n113) );
  OAI222X1 U12 ( .A0(n94), .A1(n118), .B0(n119), .B1(n545), .C0(a[4]), .C1(
        n120), .Y(n117) );
  NAND2X2 U13 ( .A(n66), .B(n535), .Y(n116) );
  NAND2X2 U14 ( .A(n531), .B(n532), .Y(n115) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n73) );
  NAND2X1 U16 ( .A(n533), .B(n75), .Y(n110) );
  CLKINVX3 U17 ( .A(n533), .Y(n26) );
  NAND2X2 U18 ( .A(a[0]), .B(n26), .Y(n156) );
  NAND2X2 U19 ( .A(n75), .B(n26), .Y(n154) );
  NAND2X1 U20 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U21 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI21XL U22 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  NAND2X1 U23 ( .A(a[4]), .B(n535), .Y(n263) );
  NAND2X1 U24 ( .A(n531), .B(a[4]), .Y(n224) );
  NAND2X2 U25 ( .A(n532), .B(a[4]), .Y(n111) );
  CLKINVX3 U26 ( .A(a[4]), .Y(n66) );
  NAND2X1 U27 ( .A(n53), .B(n556), .Y(n288) );
  CLKINVX3 U28 ( .A(n543), .Y(n540) );
  INVX1 U29 ( .A(n325), .Y(n34) );
  NAND2X1 U30 ( .A(n113), .B(n535), .Y(n214) );
  NAND2X1 U31 ( .A(n46), .B(n535), .Y(n209) );
  NAND2X1 U32 ( .A(n50), .B(n535), .Y(n301) );
  NAND2X1 U33 ( .A(n538), .B(n268), .Y(n212) );
  NAND2X1 U34 ( .A(n147), .B(n214), .Y(n207) );
  NAND2X1 U35 ( .A(n115), .B(n209), .Y(n210) );
  INVX1 U36 ( .A(n538), .Y(n53) );
  INVX1 U37 ( .A(n182), .Y(n57) );
  NOR2X1 U38 ( .A(n535), .B(n39), .Y(n325) );
  CLKINVX3 U39 ( .A(n555), .Y(n550) );
  NAND2X1 U40 ( .A(n535), .B(n71), .Y(n118) );
  NAND2X1 U41 ( .A(n56), .B(n535), .Y(n233) );
  NAND2X1 U42 ( .A(n138), .B(n535), .Y(n223) );
  NAND2X1 U43 ( .A(n39), .B(n535), .Y(n248) );
  NAND2X1 U44 ( .A(n181), .B(n535), .Y(n166) );
  NAND2X1 U45 ( .A(n229), .B(n248), .Y(n87) );
  INVX1 U46 ( .A(n102), .Y(n61) );
  NAND2X1 U47 ( .A(n115), .B(n223), .Y(n306) );
  INVX1 U48 ( .A(n168), .Y(n62) );
  INVX1 U49 ( .A(n230), .Y(n69) );
  INVX1 U50 ( .A(n116), .Y(n64) );
  INVX1 U51 ( .A(n103), .Y(n68) );
  BUFX3 U52 ( .A(n74), .Y(n535) );
  NAND2X1 U53 ( .A(n50), .B(n531), .Y(n147) );
  NAND2X1 U54 ( .A(n531), .B(n539), .Y(n120) );
  NAND2X1 U55 ( .A(n531), .B(n113), .Y(n165) );
  NAND2X1 U56 ( .A(n531), .B(n138), .Y(n182) );
  INVX1 U57 ( .A(n170), .Y(d[5]) );
  INVX1 U58 ( .A(n312), .Y(d[1]) );
  INVX1 U59 ( .A(n537), .Y(n46) );
  NAND2X1 U60 ( .A(n16), .B(n532), .Y(n259) );
  NAND2X1 U61 ( .A(n111), .B(n147), .Y(n96) );
  NOR2X1 U62 ( .A(n537), .B(n535), .Y(n124) );
  NAND2X1 U63 ( .A(n111), .B(n535), .Y(n268) );
  CLKINVX3 U64 ( .A(n111), .Y(n39) );
  NAND2X1 U65 ( .A(n531), .B(n71), .Y(n230) );
  NAND2X1 U66 ( .A(n531), .B(n66), .Y(n337) );
  NAND2BX1 U67 ( .AN(n124), .B(n263), .Y(n196) );
  INVX1 U68 ( .A(n156), .Y(n24) );
  NAND2X1 U69 ( .A(n224), .B(n268), .Y(n141) );
  NAND2BX1 U70 ( .AN(n93), .B(n537), .Y(n299) );
  NAND2X1 U71 ( .A(n224), .B(n233), .Y(n104) );
  NAND2X1 U72 ( .A(n263), .B(n142), .Y(n100) );
  CLKINVX3 U73 ( .A(n534), .Y(n21) );
  CLKINVX3 U74 ( .A(n108), .Y(n22) );
  INVX1 U76 ( .A(n249), .Y(d[3]) );
  BUFX3 U77 ( .A(a[1]), .Y(n531) );
  NAND2X1 U78 ( .A(a[7]), .B(a[2]), .Y(n94) );
  NAND2X1 U79 ( .A(n533), .B(a[0]), .Y(n108) );
  INVX1 U80 ( .A(n238), .Y(n15) );
  NAND2X1 U81 ( .A(n59), .B(n540), .Y(n114) );
  NAND2X1 U82 ( .A(n51), .B(n556), .Y(n238) );
  INVX1 U83 ( .A(n288), .Y(n14) );
  NOR2X1 U84 ( .A(n550), .B(n325), .Y(n199) );
  NOR2X1 U85 ( .A(n49), .B(n62), .Y(n247) );
  NAND2X1 U86 ( .A(n222), .B(n540), .Y(n162) );
  INVX1 U87 ( .A(n301), .Y(n49) );
  INVX1 U88 ( .A(n166), .Y(n60) );
  INVX1 U89 ( .A(n207), .Y(n48) );
  INVX1 U90 ( .A(n228), .Y(n51) );
  INVX4 U91 ( .A(n536), .Y(n556) );
  NOR2BX1 U92 ( .AN(n214), .B(n69), .Y(n88) );
  NOR2X1 U93 ( .A(n53), .B(n70), .Y(n326) );
  NOR2X1 U94 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U95 ( .A(n34), .B(n223), .Y(n183) );
  INVX1 U96 ( .A(n118), .Y(n70) );
  NAND2X1 U97 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U98 ( .A(n233), .Y(n55) );
  INVX1 U99 ( .A(n223), .Y(n59) );
  NOR2X1 U100 ( .A(n57), .B(n55), .Y(n197) );
  INVX1 U101 ( .A(n248), .Y(n37) );
  OAI221XL U102 ( .A0(n58), .A1(n545), .B0(n98), .B1(n94), .C0(n18), .Y(n347)
         );
  INVX1 U103 ( .A(n199), .Y(n18) );
  INVX1 U104 ( .A(n127), .Y(n35) );
  NOR2X1 U105 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U106 ( .A(n212), .Y(n41) );
  NOR2X1 U107 ( .A(n62), .B(n55), .Y(n145) );
  INVX1 U108 ( .A(n306), .Y(n58) );
  INVX1 U109 ( .A(n158), .Y(n42) );
  INVX1 U110 ( .A(n87), .Y(n38) );
  INVX1 U111 ( .A(n210), .Y(n44) );
  NAND2X1 U112 ( .A(n63), .B(n535), .Y(n243) );
  OAI22X1 U113 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U114 ( .A0(n61), .A1(n547), .B0(n556), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U115 ( .A0(n556), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U116 ( .A(n116), .B(n229), .Y(n244) );
  NOR2X1 U117 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U118 ( .A0(n542), .A1(n207), .B0(n545), .B1(n538), .Y(n242) );
  CLKINVX3 U119 ( .A(n113), .Y(n50) );
  NAND2X1 U120 ( .A(n214), .B(n142), .Y(n90) );
  CLKINVX3 U121 ( .A(n181), .Y(n63) );
  AOI22X1 U122 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U123 ( .A0(n98), .A1(n545), .B0(n30), .B1(n542), .C0(n99), .Y(n91)
         );
  OAI221XL U124 ( .A0(n42), .A1(n545), .B0(n51), .B1(n542), .C0(n95), .Y(n92)
         );
  INVX1 U125 ( .A(n104), .Y(n30) );
  NAND2X1 U126 ( .A(n556), .B(n96), .Y(n187) );
  NAND2X1 U127 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U128 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  OAI221XL U129 ( .A0(n46), .A1(n551), .B0(n63), .B1(n545), .C0(n200), .Y(n194) );
  OAI221XL U130 ( .A0(n536), .A1(n196), .B0(n197), .B1(n545), .C0(n198), .Y(
        n195) );
  AOI211X1 U131 ( .A0(n201), .A1(n556), .B0(n202), .C0(n203), .Y(n200) );
  AOI22X1 U132 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U133 ( .A0(n35), .A1(n545), .B0(n44), .B1(n543), .C0(n333), .Y(n332) );
  OAI211X1 U134 ( .A0(n326), .A1(n550), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U135 ( .A0(n35), .A1(n556), .B0(n39), .B1(n554), .Y(n333) );
  AOI22X1 U136 ( .A0(n548), .A1(n63), .B0(n247), .B1(n539), .Y(n334) );
  AOI21X1 U137 ( .A0(n115), .A1(n243), .B0(n550), .Y(n360) );
  INVX1 U138 ( .A(n120), .Y(n4) );
  AND2X2 U139 ( .A(n165), .B(n166), .Y(n129) );
  NAND2X1 U140 ( .A(n538), .B(n214), .Y(n126) );
  OAI21XL U141 ( .A0(n165), .A1(n550), .B0(n187), .Y(n266) );
  INVX1 U142 ( .A(n284), .Y(n10) );
  OAI31X1 U143 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U144 ( .A0(n541), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U145 ( .A(n147), .Y(n47) );
  OAI22X1 U146 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U147 ( .A0(n556), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U148 ( .A0(n11), .A1(n535), .B0(n27), .B1(n556), .C0(n307), .Y(n302) );
  OAI22X1 U149 ( .A0(n64), .A1(n542), .B0(n550), .B1(n306), .Y(n304) );
  AOI222X1 U150 ( .A0(n56), .A1(n540), .B0(n60), .B1(n554), .C0(n548), .C1(n71), .Y(n356) );
  AOI21X1 U151 ( .A0(n50), .A1(n16), .B0(n366), .Y(n365) );
  OAI221XL U152 ( .A0(n551), .A1(n87), .B0(n94), .B1(n104), .C0(n246), .Y(n235) );
  AOI2BB2X1 U153 ( .B0(n11), .B1(n535), .A0N(n536), .A1N(n247), .Y(n246) );
  CLKINVX8 U154 ( .A(n546), .Y(n545) );
  CLKINVX3 U155 ( .A(n541), .Y(n539) );
  NOR2X1 U156 ( .A(n545), .B(n535), .Y(n202) );
  AOI211X1 U157 ( .A0(n45), .A1(n540), .B0(n204), .C0(n205), .Y(n192) );
  INVX1 U158 ( .A(n209), .Y(n45) );
  NAND2BX1 U159 ( .AN(n97), .B(n206), .Y(n205) );
  AOI222X1 U160 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n540), 
        .Y(n198) );
  AOI221X1 U161 ( .A0(n321), .A1(n553), .B0(n540), .B1(n311), .C0(n327), .Y(
        n315) );
  OAI221XL U162 ( .A0(n536), .A1(n209), .B0(n545), .B1(n103), .C0(n288), .Y(
        n327) );
  AOI221X1 U163 ( .A0(n4), .A1(n71), .B0(n553), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI2BB1X1 U164 ( .A0N(n142), .A1N(n547), .B0(n187), .Y(n186) );
  OAI221XL U165 ( .A0(n308), .A1(n551), .B0(n545), .B1(n165), .C0(n162), .Y(
        n307) );
  NOR2X1 U166 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U167 ( .A0(n54), .A1(n545), .B0(n33), .B1(n542), .C0(n232), .Y(n217) );
  INVX1 U168 ( .A(n234), .Y(n54) );
  AOI32X1 U169 ( .A0(n34), .A1(n181), .A2(n556), .B0(n553), .B1(n233), .Y(n232) );
  OAI221XL U170 ( .A0(n67), .A1(n551), .B0(n94), .B1(n538), .C0(n294), .Y(n282) );
  INVX1 U171 ( .A(n115), .Y(n67) );
  AOI211X1 U172 ( .A0(n48), .A1(n556), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U173 ( .A(n114), .Y(n6) );
  AOI211X1 U174 ( .A0(n60), .A1(n540), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U175 ( .A(n545), .B(n39), .C(n61), .Y(n364) );
  INVX1 U176 ( .A(n259), .Y(n13) );
  OAI221XL U177 ( .A0(n536), .A1(n168), .B0(n164), .B1(n551), .C0(n169), .Y(
        n150) );
  AOI22X1 U178 ( .A0(n549), .A1(n34), .B0(n48), .B1(n539), .Y(n169) );
  AOI211X1 U179 ( .A0(n554), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  CLKINVX3 U180 ( .A(n555), .Y(n551) );
  INVX1 U181 ( .A(n125), .Y(n7) );
  AOI221X1 U182 ( .A0(n126), .A1(n552), .B0(n127), .B1(n549), .C0(n128), .Y(
        n125) );
  OAI21XL U183 ( .A0(n536), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U184 ( .A(n536), .Y(n16) );
  NOR2X1 U185 ( .A(n39), .B(n57), .Y(n179) );
  CLKINVX3 U186 ( .A(n110), .Y(n23) );
  NAND3X1 U187 ( .A(n538), .B(n113), .C(n540), .Y(n89) );
  NAND2X1 U188 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U189 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U190 ( .A(n538), .B(n166), .Y(n311) );
  NOR2BX1 U191 ( .AN(n229), .B(n68), .Y(n164) );
  AOI21X1 U192 ( .A0(n181), .A1(n182), .B0(n536), .Y(n180) );
  OAI221XL U193 ( .A0(n36), .A1(n550), .B0(n121), .B1(n543), .C0(n140), .Y(
        n135) );
  INVX1 U194 ( .A(n85), .Y(n36) );
  AOI22X1 U195 ( .A0(n49), .A1(n549), .B0(n556), .B1(n141), .Y(n140) );
  AOI22X1 U196 ( .A0(n57), .A1(n546), .B0(n555), .B1(n113), .Y(n239) );
  AOI22X1 U197 ( .A0(n547), .A1(n311), .B0(n50), .B1(n539), .Y(n350) );
  NOR2X1 U198 ( .A(n138), .B(n536), .Y(n97) );
  NAND2X1 U199 ( .A(n243), .B(n142), .Y(n127) );
  INVX1 U200 ( .A(n154), .Y(n25) );
  NAND2X1 U201 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U202 ( .A(n138), .Y(n56) );
  NAND2X1 U203 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U204 ( .A(n64), .B(n124), .Y(n121) );
  AOI211X1 U205 ( .A0(n556), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  OAI2BB2X1 U206 ( .B0(n545), .B1(n183), .A0N(n188), .A1N(n540), .Y(n335) );
  AOI21X1 U207 ( .A0(n301), .A1(n337), .B0(n550), .Y(n336) );
  NAND2X1 U208 ( .A(n138), .B(n102), .Y(n227) );
  NAND2X1 U209 ( .A(n103), .B(n165), .Y(n188) );
  AOI21X1 U210 ( .A0(n16), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U211 ( .A0(n102), .A1(n103), .B0(n550), .Y(n101) );
  INVX1 U212 ( .A(n337), .Y(n65) );
  AOI22X1 U213 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  OAI221XL U214 ( .A0(n65), .A1(n551), .B0(n31), .B1(n536), .C0(n149), .Y(n143) );
  OAI221XL U215 ( .A0(n145), .A1(n545), .B0(n28), .B1(n551), .C0(n146), .Y(
        n144) );
  AOI2BB2X1 U216 ( .B0(n539), .B1(n87), .A0N(n545), .A1N(n121), .Y(n149) );
  INVX1 U217 ( .A(n208), .Y(n29) );
  INVX1 U218 ( .A(n299), .Y(n11) );
  INVX1 U219 ( .A(n100), .Y(n33) );
  AOI221XL U220 ( .A0(n556), .A1(n52), .B0(n548), .B1(n123), .C0(n324), .Y(
        n316) );
  INVX1 U221 ( .A(n326), .Y(n52) );
  OAI32X1 U222 ( .A0(n94), .A1(n63), .A2(n325), .B0(n37), .B1(n551), .Y(n324)
         );
  INVX1 U223 ( .A(n196), .Y(n31) );
  OAI221XL U224 ( .A0(n56), .A1(n545), .B0(n32), .B1(n543), .C0(n163), .Y(n151) );
  INVX1 U225 ( .A(n167), .Y(n32) );
  AOI22X1 U226 ( .A0(n164), .A1(n16), .B0(n129), .B1(n554), .Y(n163) );
  INVX1 U227 ( .A(n141), .Y(n27) );
  INVX1 U228 ( .A(n148), .Y(n28) );
  OAI221XL U229 ( .A0(n40), .A1(n551), .B0(n58), .B1(n545), .C0(n137), .Y(n136) );
  INVX1 U230 ( .A(n96), .Y(n40) );
  AOI31X1 U231 ( .A0(n102), .A1(n138), .A2(n556), .B0(n8), .Y(n137) );
  INVX1 U232 ( .A(n89), .Y(n8) );
  INVX1 U233 ( .A(n185), .Y(n19) );
  INVX1 U234 ( .A(n544), .Y(n543) );
  INVX1 U235 ( .A(n539), .Y(n542) );
  OAI22X2 U236 ( .A0(n534), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  AOI211X1 U237 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U238 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI2BB2X1 U239 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  OAI22X2 U240 ( .A0(n534), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  AOI211X1 U241 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U242 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U243 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  OAI21X2 U244 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  OAI2BB1X1 U245 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI221X1 U246 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76)
         );
  AOI22X1 U247 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  AOI22X1 U248 ( .A0(n533), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U249 ( .A0(n61), .A1(n551), .B0(n545), .B1(n260), .C0(n261), .Y(
        n254) );
  OAI221XL U250 ( .A0(n41), .A1(n545), .B0(n542), .B1(n181), .C0(n256), .Y(
        n255) );
  AOI21X1 U251 ( .A0(n33), .A1(n556), .B0(n262), .Y(n261) );
  AOI22X1 U252 ( .A0(n348), .A1(n26), .B0(n533), .B1(n349), .Y(n342) );
  OAI221XL U253 ( .A0(n536), .A1(n166), .B0(n286), .B1(n545), .C0(n351), .Y(
        n348) );
  OAI211X1 U254 ( .A0(n88), .A1(n550), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U255 ( .B0(n539), .B1(n196), .A0N(n550), .A1N(n179), .Y(n351) );
  OAI22X1 U256 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U257 ( .A0(n549), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U258 ( .A0(n56), .A1(n4), .B0(n547), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U259 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U260 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U261 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U262 ( .A0(n61), .A1(n552), .B0(n547), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U263 ( .A0(n541), .A1(n71), .B0(n37), .B1(n550), .Y(n157) );
  OAI22X1 U264 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U265 ( .A0(n549), .A1(n111), .B0(n47), .B1(n540), .C0(n112), .Y(
        n109) );
  AOI221X1 U266 ( .A0(n556), .A1(n115), .B0(n552), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U267 ( .A0(n536), .A1(n113), .B0(n44), .B1(n551), .C0(n114), .Y(
        n112) );
  AOI211X1 U268 ( .A0(n55), .A1(n556), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U269 ( .A0(n114), .A1(n206), .A2(n273), .B0(n533), .Y(n272) );
  OAI22X1 U270 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U271 ( .B0(n70), .B1(n552), .A0N(n90), .A1N(n545), .Y(n273) );
  AOI2BB2X1 U272 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  OAI221XL U273 ( .A0(n46), .A1(n551), .B0(n545), .B1(n116), .C0(n267), .Y(
        n264) );
  AOI221XL U274 ( .A0(n548), .A1(n247), .B0(n212), .B1(n540), .C0(n266), .Y(
        n265) );
  AOI22X1 U275 ( .A0(n539), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  AOI22X1 U276 ( .A0(n534), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U277 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  OAI221XL U278 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  AOI22X1 U279 ( .A0(n171), .A1(n21), .B0(n534), .B1(n172), .Y(n170) );
  OAI221XL U281 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  OAI221XL U282 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  AOI22X1 U283 ( .A0(n552), .A1(n532), .B0(n539), .B1(n66), .Y(n292) );
  AOI22X1 U284 ( .A0(n533), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U285 ( .A0(n43), .A1(n545), .B0(n542), .B1(n34), .C0(n365), .Y(n361) );
  OAI221XL U286 ( .A0(n532), .A1(n120), .B0(n201), .B1(n551), .C0(n363), .Y(
        n362) );
  INVX1 U287 ( .A(n260), .Y(n43) );
  AOI22X1 U288 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  OAI21XL U289 ( .A0(n321), .A1(n536), .B0(n322), .Y(n318) );
  OAI221XL U290 ( .A0(n551), .A1(n113), .B0(n88), .B1(n545), .C0(n320), .Y(
        n319) );
  AOI31X1 U291 ( .A0(n538), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  CLKINVX3 U292 ( .A(n532), .Y(n71) );
  OAI21XL U293 ( .A0(n545), .A1(n537), .B0(n120), .Y(n276) );
  NAND2X1 U294 ( .A(n63), .B(n531), .Y(n168) );
  AOI21X1 U295 ( .A0(n224), .A1(n243), .B0(n545), .Y(n295) );
  INVX1 U296 ( .A(n531), .Y(n74) );
  OAI21XL U297 ( .A0(n73), .A1(n301), .B0(n550), .Y(n323) );
  OAI21XL U298 ( .A0(n73), .A1(n243), .B0(n550), .Y(n245) );
  OAI21XL U299 ( .A0(n536), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U300 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U301 ( .A(n162), .Y(n5) );
  AOI211X1 U302 ( .A0(n39), .A1(n540), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U303 ( .A0(n551), .A1(n116), .B0(n73), .B1(n230), .C0(n545), .C1(
        n102), .Y(n275) );
  NAND2X1 U304 ( .A(n62), .B(n554), .Y(n287) );
  OAI21X2 U305 ( .A0(n534), .A1(n131), .B0(n132), .Y(d[6]) );
  OAI2BB1X1 U306 ( .A0N(n133), .A1N(n134), .B0(n534), .Y(n132) );
  AOI221X1 U307 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131) );
  AOI22X1 U308 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  NOR2BX1 U309 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U310 ( .A(n82), .Y(n536) );
  NAND2X1 U311 ( .A(n73), .B(n20), .Y(n82) );
  OAI221XL U312 ( .A0(n531), .A1(n259), .B0(n543), .B1(n214), .C0(n287), .Y(
        n293) );
  BUFX3 U313 ( .A(n139), .Y(n538) );
  NAND2X1 U314 ( .A(n531), .B(n537), .Y(n139) );
  AOI211X1 U315 ( .A0(n540), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  OAI222X1 U316 ( .A0(n551), .A1(n167), .B0(n339), .B1(n536), .C0(n545), .C1(
        n34), .Y(n338) );
  AOI21X1 U317 ( .A0(n537), .A1(n535), .B0(n65), .Y(n339) );
  AOI211X1 U318 ( .A0(n533), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  OAI221XL U319 ( .A0(n545), .A1(n116), .B0(n321), .B1(n541), .C0(n359), .Y(
        n354) );
  AOI21X1 U320 ( .A0(n356), .A1(n357), .B0(n533), .Y(n355) );
  AOI31X1 U321 ( .A0(n556), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  INVX1 U322 ( .A(n93), .Y(n546) );
  INVX1 U323 ( .A(n83), .Y(n554) );
  INVX1 U324 ( .A(n83), .Y(n555) );
  INVX1 U325 ( .A(n544), .Y(n541) );
  INVX1 U326 ( .A(n94), .Y(n544) );
  AOI22X1 U327 ( .A0(n533), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U328 ( .A0(n545), .A1(n141), .B0(n551), .B1(n263), .C0(n29), .C1(
        n541), .Y(n277) );
  OAI221XL U329 ( .A0(n31), .A1(n536), .B0(n551), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U330 ( .B0(n88), .B1(n539), .A0N(n545), .A1N(n197), .Y(n279) );
  NAND2X1 U331 ( .A(n224), .B(n301), .Y(n148) );
  NOR2BX1 U332 ( .AN(n263), .B(n61), .Y(n321) );
  AOI21X1 U333 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI22X1 U334 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U335 ( .A0(n63), .A1(n545), .B0(n542), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U336 ( .A0(n38), .A1(n536), .B0(n545), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U337 ( .A0(n179), .A1(n552), .B0(n180), .Y(n178) );
  AOI22X1 U338 ( .A0(n556), .A1(n66), .B0(n539), .B1(n147), .Y(n146) );
  AOI22X1 U339 ( .A0(n548), .A1(n85), .B0(n41), .B1(n539), .Y(n84) );
  AOI31X1 U340 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U341 ( .A0N(n223), .A1N(n224), .B0(n553), .Y(n220) );
  AOI22X1 U342 ( .A0(n29), .A1(n556), .B0(n222), .B1(n547), .Y(n221) );
  NAND2X1 U343 ( .A(n224), .B(n118), .Y(n208) );
  NAND2X1 U344 ( .A(n263), .B(n337), .Y(n167) );
  AOI21X1 U345 ( .A0(n263), .A1(n182), .B0(n545), .Y(n305) );
  AOI21X1 U346 ( .A0(n111), .A1(n538), .B0(n541), .Y(n203) );
  NAND2X1 U347 ( .A(n16), .B(n531), .Y(n206) );
  XNOR2X1 U348 ( .A(n20), .B(n531), .Y(n185) );
  NAND2X1 U349 ( .A(n539), .B(n537), .Y(n130) );
  XNOR2X1 U350 ( .A(n73), .B(n531), .Y(n161) );
  AOI21X1 U351 ( .A0(n90), .A1(n73), .B0(n556), .Y(n86) );
  AOI221X1 U352 ( .A0(n46), .A1(n540), .B0(n553), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U353 ( .A0(n536), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U354 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  AOI222X1 U355 ( .A0(n549), .A1(n210), .B0(n211), .B1(n212), .C0(n556), .C1(
        n537), .Y(n191) );
  OAI21XL U356 ( .A0(n73), .A1(n214), .B0(n550), .Y(n211) );
  AOI31X1 U357 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U358 ( .A0(n148), .A1(n73), .B0(n29), .B1(n553), .Y(n300) );
  INVX1 U359 ( .A(n93), .Y(n547) );
  INVX1 U360 ( .A(n93), .Y(n549) );
  INVX1 U361 ( .A(n93), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n358) );
  INVX1 U363 ( .A(n83), .Y(n552) );
  INVX1 U364 ( .A(n83), .Y(n553) );
  NOR2BX1 U365 ( .AN(n93), .B(n554), .Y(n309) );
  OAI22X2 U366 ( .A0(n340), .A1(n21), .B0(n534), .B1(n341), .Y(d[0]) );
  AOI22X1 U367 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U368 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI22X1 U369 ( .A0(n347), .A1(n26), .B0(n556), .B1(n90), .Y(n343) );
  AOI22X1 U370 ( .A0(n250), .A1(n21), .B0(n534), .B1(n251), .Y(n249) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  OAI22X1 U373 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U374 ( .A0(n548), .A1(n230), .B0(n556), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U375 ( .A0(n164), .A1(n547), .B0(a[2]), .B1(n227), .C0(n556), .C1(
        n228), .Y(n226) );
  OAI22X1 U376 ( .A0(n35), .A1(n543), .B0(n550), .B1(n537), .Y(n231) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI21XL U383 ( .A0(n66), .A1(n550), .B0(n259), .Y(n257) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI22X1 U385 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U386 ( .A(a[0]), .Y(n75) );
  AOI211X1 U387 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U388 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U389 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U390 ( .A(a[5]), .Y(n533) );
  OAI221XL U391 ( .A0(n536), .A1(n115), .B0(n121), .B1(n545), .C0(n122), .Y(
        n105) );
  AOI22X1 U392 ( .A0(n539), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  AOI33X1 U393 ( .A0(n532), .A1(n540), .A2(n19), .B0(n185), .B1(n181), .B2(
        a[2]), .Y(n184) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_16 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556;

  OAI221X4 U4 ( .A0(n66), .A1(n536), .B0(n61), .B1(n551), .C0(n84), .Y(n81) );
  OAI221X4 U6 ( .A0(n86), .A1(n87), .B0(n88), .B1(n551), .C0(n89), .Y(n80) );
  OAI222X4 U75 ( .A0(n551), .A1(n207), .B0(n181), .B1(n120), .C0(n545), .C1(
        n208), .Y(n204) );
  OAI32X4 U280 ( .A0(n551), .A1(n56), .A2(n53), .B0(n94), .B1(n103), .Y(n366)
         );
  AOI221X1 U1 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n103) );
  OAI222X1 U5 ( .A0(n94), .A1(n118), .B0(n119), .B1(n545), .C0(a[4]), .C1(n120), .Y(n117) );
  NAND2X2 U7 ( .A(n531), .B(n532), .Y(n115) );
  NAND2X1 U8 ( .A(n56), .B(n531), .Y(n229) );
  NAND2X2 U9 ( .A(n532), .B(n66), .Y(n181) );
  NAND2X1 U10 ( .A(n39), .B(n531), .Y(n142) );
  NAND2X2 U11 ( .A(n537), .B(n181), .Y(n113) );
  NAND2X2 U12 ( .A(n66), .B(n535), .Y(n116) );
  NAND2X2 U13 ( .A(n66), .B(n71), .Y(n138) );
  NAND2X1 U14 ( .A(n531), .B(n181), .Y(n102) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n73) );
  NAND2X1 U16 ( .A(n533), .B(n75), .Y(n110) );
  CLKINVX3 U17 ( .A(n533), .Y(n26) );
  NAND2X2 U18 ( .A(n75), .B(n26), .Y(n154) );
  NAND2X2 U19 ( .A(a[0]), .B(n26), .Y(n156) );
  CLKINVX3 U20 ( .A(n534), .Y(n21) );
  OAI22X2 U21 ( .A0(n340), .A1(n21), .B0(n534), .B1(n341), .Y(d[0]) );
  OAI22X2 U22 ( .A0(n534), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  INVX1 U23 ( .A(n249), .Y(d[3]) );
  OAI21X2 U24 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  AOI221X1 U25 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76) );
  OAI22X2 U26 ( .A0(n534), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  OAI21X2 U27 ( .A0(n534), .A1(n131), .B0(n132), .Y(d[6]) );
  AOI221X1 U28 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131)
         );
  NAND2X1 U29 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U30 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI21XL U31 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  NAND2X1 U32 ( .A(a[4]), .B(n535), .Y(n263) );
  NAND2X1 U33 ( .A(n531), .B(a[4]), .Y(n224) );
  NAND2X2 U34 ( .A(n532), .B(a[4]), .Y(n111) );
  CLKINVX3 U35 ( .A(a[4]), .Y(n66) );
  NAND2X1 U36 ( .A(n53), .B(n16), .Y(n288) );
  CLKINVX3 U37 ( .A(n542), .Y(n540) );
  INVX1 U38 ( .A(n325), .Y(n34) );
  NAND2X1 U39 ( .A(n113), .B(n535), .Y(n214) );
  NAND2X1 U40 ( .A(n56), .B(n535), .Y(n233) );
  NAND2X1 U41 ( .A(n46), .B(n535), .Y(n209) );
  NAND2X1 U42 ( .A(n50), .B(n535), .Y(n301) );
  NAND2X1 U43 ( .A(n538), .B(n268), .Y(n212) );
  NAND2X1 U44 ( .A(n147), .B(n214), .Y(n207) );
  NAND2X1 U45 ( .A(n115), .B(n209), .Y(n210) );
  INVX1 U46 ( .A(n168), .Y(n62) );
  INVX1 U47 ( .A(n538), .Y(n53) );
  INVX1 U48 ( .A(n182), .Y(n57) );
  NOR2X1 U49 ( .A(n535), .B(n39), .Y(n325) );
  CLKINVX3 U50 ( .A(n555), .Y(n550) );
  NAND2X1 U51 ( .A(n535), .B(n71), .Y(n118) );
  NAND2X1 U52 ( .A(n138), .B(n535), .Y(n223) );
  NAND2X1 U53 ( .A(n39), .B(n535), .Y(n248) );
  NAND2X1 U54 ( .A(n181), .B(n535), .Y(n166) );
  NAND2X1 U55 ( .A(n229), .B(n248), .Y(n87) );
  INVX1 U56 ( .A(n102), .Y(n61) );
  NAND2X1 U57 ( .A(n115), .B(n223), .Y(n306) );
  INVX1 U58 ( .A(n230), .Y(n69) );
  INVX1 U59 ( .A(n116), .Y(n64) );
  INVX1 U60 ( .A(n103), .Y(n68) );
  BUFX3 U61 ( .A(n74), .Y(n535) );
  NAND2X1 U62 ( .A(n50), .B(n531), .Y(n147) );
  NAND2X1 U63 ( .A(n531), .B(n539), .Y(n120) );
  NAND2X1 U64 ( .A(n111), .B(n535), .Y(n268) );
  NAND2X1 U65 ( .A(n531), .B(n113), .Y(n165) );
  NAND2X1 U66 ( .A(n531), .B(n138), .Y(n182) );
  INVX1 U67 ( .A(n312), .Y(d[1]) );
  INVX1 U68 ( .A(n170), .Y(d[5]) );
  INVX1 U69 ( .A(n537), .Y(n46) );
  NAND2X1 U70 ( .A(n16), .B(n532), .Y(n259) );
  NAND2X1 U71 ( .A(n111), .B(n147), .Y(n96) );
  NOR2X1 U72 ( .A(n537), .B(n535), .Y(n124) );
  CLKINVX3 U73 ( .A(n111), .Y(n39) );
  NAND2X1 U74 ( .A(n531), .B(n71), .Y(n230) );
  NAND2X1 U76 ( .A(n531), .B(n66), .Y(n337) );
  NAND2BX1 U77 ( .AN(n124), .B(n263), .Y(n196) );
  INVX1 U78 ( .A(n156), .Y(n24) );
  NAND2X1 U79 ( .A(n224), .B(n268), .Y(n141) );
  NAND2BX1 U80 ( .AN(n93), .B(n537), .Y(n299) );
  NAND2X1 U81 ( .A(n224), .B(n233), .Y(n104) );
  NAND2X1 U82 ( .A(n263), .B(n142), .Y(n100) );
  CLKINVX3 U83 ( .A(n108), .Y(n22) );
  BUFX3 U84 ( .A(a[1]), .Y(n531) );
  NAND2X1 U85 ( .A(a[7]), .B(a[2]), .Y(n94) );
  NAND2X1 U86 ( .A(n533), .B(a[0]), .Y(n108) );
  INVX1 U87 ( .A(n238), .Y(n15) );
  NAND2X1 U88 ( .A(n59), .B(n540), .Y(n114) );
  NAND2X1 U89 ( .A(n51), .B(n556), .Y(n238) );
  INVX1 U90 ( .A(n288), .Y(n14) );
  NOR2X1 U91 ( .A(n550), .B(n325), .Y(n199) );
  NOR2X1 U92 ( .A(n49), .B(n62), .Y(n247) );
  NAND2X1 U93 ( .A(n222), .B(n540), .Y(n162) );
  INVX1 U94 ( .A(n301), .Y(n49) );
  INVX1 U95 ( .A(n166), .Y(n60) );
  INVX1 U96 ( .A(n207), .Y(n48) );
  INVX1 U97 ( .A(n228), .Y(n51) );
  INVX4 U98 ( .A(n536), .Y(n556) );
  NOR2BX1 U99 ( .AN(n214), .B(n69), .Y(n88) );
  NOR2X1 U100 ( .A(n53), .B(n70), .Y(n326) );
  NOR2X1 U101 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U102 ( .A(n34), .B(n223), .Y(n183) );
  INVX1 U103 ( .A(n118), .Y(n70) );
  NAND2X1 U104 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U105 ( .A(n233), .Y(n55) );
  INVX1 U106 ( .A(n223), .Y(n59) );
  NOR2X1 U107 ( .A(n57), .B(n55), .Y(n197) );
  INVX1 U108 ( .A(n248), .Y(n37) );
  OAI221XL U109 ( .A0(n58), .A1(n545), .B0(n98), .B1(n542), .C0(n18), .Y(n347)
         );
  INVX1 U110 ( .A(n199), .Y(n18) );
  INVX1 U111 ( .A(n127), .Y(n35) );
  NOR2X1 U112 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U113 ( .A(n212), .Y(n41) );
  NOR2X1 U114 ( .A(n62), .B(n55), .Y(n145) );
  INVX1 U115 ( .A(n306), .Y(n58) );
  INVX1 U116 ( .A(n158), .Y(n42) );
  INVX1 U117 ( .A(n87), .Y(n38) );
  INVX1 U118 ( .A(n210), .Y(n44) );
  NAND2X1 U119 ( .A(n63), .B(n535), .Y(n243) );
  OAI22X1 U120 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U121 ( .A0(n61), .A1(n547), .B0(n556), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U122 ( .A0(n556), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U123 ( .A(n116), .B(n229), .Y(n244) );
  NOR2X1 U124 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U125 ( .A0(n542), .A1(n207), .B0(n545), .B1(n538), .Y(n242) );
  CLKINVX3 U126 ( .A(n113), .Y(n50) );
  CLKINVX3 U127 ( .A(n181), .Y(n63) );
  AOI22X1 U128 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U129 ( .A0(n98), .A1(n545), .B0(n30), .B1(n543), .C0(n99), .Y(n91)
         );
  OAI221XL U130 ( .A0(n42), .A1(n545), .B0(n51), .B1(n543), .C0(n95), .Y(n92)
         );
  INVX1 U131 ( .A(n104), .Y(n30) );
  NAND2X1 U132 ( .A(n556), .B(n96), .Y(n187) );
  NAND2X1 U133 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U134 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  OAI221XL U135 ( .A0(n46), .A1(n551), .B0(n63), .B1(n545), .C0(n200), .Y(n194) );
  OAI221XL U136 ( .A0(n536), .A1(n196), .B0(n197), .B1(n545), .C0(n198), .Y(
        n195) );
  AOI211X1 U137 ( .A0(n201), .A1(n556), .B0(n202), .C0(n203), .Y(n200) );
  AOI22X1 U138 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U139 ( .A0(n35), .A1(n545), .B0(n44), .B1(n543), .C0(n333), .Y(n332) );
  OAI211X1 U140 ( .A0(n326), .A1(n550), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U141 ( .A0(n35), .A1(n556), .B0(n39), .B1(n554), .Y(n333) );
  AOI22X1 U142 ( .A0(n548), .A1(n63), .B0(n247), .B1(n539), .Y(n334) );
  AOI21X1 U143 ( .A0(n115), .A1(n243), .B0(n550), .Y(n360) );
  INVX1 U144 ( .A(n120), .Y(n4) );
  AND2X2 U145 ( .A(n165), .B(n166), .Y(n129) );
  OAI21XL U146 ( .A0(n165), .A1(n550), .B0(n187), .Y(n266) );
  INVX1 U147 ( .A(n284), .Y(n10) );
  OAI31X1 U148 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U149 ( .A0(n541), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U150 ( .A(n147), .Y(n47) );
  OAI22X1 U151 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U152 ( .A0(n556), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U153 ( .A0(n11), .A1(n535), .B0(n27), .B1(n556), .C0(n307), .Y(n302) );
  OAI22X1 U154 ( .A0(n64), .A1(n543), .B0(n550), .B1(n306), .Y(n304) );
  AOI222X1 U155 ( .A0(n56), .A1(n540), .B0(n60), .B1(n554), .C0(n549), .C1(n71), .Y(n356) );
  AOI21X1 U156 ( .A0(n50), .A1(n556), .B0(n366), .Y(n365) );
  OAI221XL U157 ( .A0(n551), .A1(n87), .B0(n94), .B1(n104), .C0(n246), .Y(n235) );
  AOI2BB2X1 U158 ( .B0(n11), .B1(n535), .A0N(n536), .A1N(n247), .Y(n246) );
  CLKINVX8 U159 ( .A(n546), .Y(n545) );
  CLKINVX3 U160 ( .A(n541), .Y(n539) );
  NOR2X1 U161 ( .A(n545), .B(n535), .Y(n202) );
  AOI211X1 U162 ( .A0(n45), .A1(n540), .B0(n204), .C0(n205), .Y(n192) );
  INVX1 U163 ( .A(n209), .Y(n45) );
  NAND2BX1 U164 ( .AN(n97), .B(n206), .Y(n205) );
  AOI222X1 U165 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n540), 
        .Y(n198) );
  AOI221X1 U166 ( .A0(n321), .A1(n553), .B0(n540), .B1(n311), .C0(n327), .Y(
        n315) );
  OAI221XL U167 ( .A0(n536), .A1(n209), .B0(n545), .B1(n103), .C0(n288), .Y(
        n327) );
  AOI221X1 U168 ( .A0(n4), .A1(n71), .B0(n553), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI2BB1X1 U169 ( .A0N(n142), .A1N(n547), .B0(n187), .Y(n186) );
  OAI221XL U170 ( .A0(n308), .A1(n551), .B0(n545), .B1(n165), .C0(n162), .Y(
        n307) );
  NOR2X1 U171 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U172 ( .A0(n54), .A1(n545), .B0(n33), .B1(n543), .C0(n232), .Y(n217) );
  INVX1 U173 ( .A(n234), .Y(n54) );
  AOI32X1 U174 ( .A0(n34), .A1(n181), .A2(n556), .B0(n553), .B1(n233), .Y(n232) );
  OAI221XL U175 ( .A0(n67), .A1(n551), .B0(n94), .B1(n538), .C0(n294), .Y(n282) );
  INVX1 U176 ( .A(n115), .Y(n67) );
  AOI211X1 U177 ( .A0(n48), .A1(n556), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U178 ( .A(n114), .Y(n6) );
  AOI211X1 U179 ( .A0(n60), .A1(n540), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U180 ( .A(n545), .B(n39), .C(n61), .Y(n364) );
  INVX1 U181 ( .A(n259), .Y(n13) );
  OAI221XL U182 ( .A0(n536), .A1(n168), .B0(n164), .B1(n551), .C0(n169), .Y(
        n150) );
  AOI22X1 U183 ( .A0(n549), .A1(n34), .B0(n48), .B1(n539), .Y(n169) );
  AOI211X1 U184 ( .A0(n554), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  CLKINVX3 U185 ( .A(n555), .Y(n551) );
  INVX1 U186 ( .A(n544), .Y(n542) );
  INVX1 U187 ( .A(n125), .Y(n7) );
  AOI221X1 U188 ( .A0(n126), .A1(n552), .B0(n127), .B1(n548), .C0(n128), .Y(
        n125) );
  OAI21XL U189 ( .A0(n536), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U190 ( .A(n536), .Y(n16) );
  NOR2X1 U191 ( .A(n39), .B(n57), .Y(n179) );
  CLKINVX3 U192 ( .A(n110), .Y(n23) );
  NAND3X1 U193 ( .A(n538), .B(n113), .C(n540), .Y(n89) );
  NAND2X1 U194 ( .A(n214), .B(n142), .Y(n90) );
  NAND2X1 U195 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U196 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U197 ( .A(n538), .B(n166), .Y(n311) );
  NOR2BX1 U198 ( .AN(n229), .B(n68), .Y(n164) );
  AOI21X1 U199 ( .A0(n181), .A1(n182), .B0(n536), .Y(n180) );
  OAI221XL U200 ( .A0(n36), .A1(n550), .B0(n121), .B1(n541), .C0(n140), .Y(
        n135) );
  INVX1 U201 ( .A(n85), .Y(n36) );
  AOI22X1 U202 ( .A0(n49), .A1(n548), .B0(n556), .B1(n141), .Y(n140) );
  AOI22X1 U203 ( .A0(n57), .A1(n546), .B0(n555), .B1(n113), .Y(n239) );
  AOI22X1 U204 ( .A0(n547), .A1(n311), .B0(n50), .B1(n539), .Y(n350) );
  NOR2X1 U205 ( .A(n138), .B(n536), .Y(n97) );
  NAND2X1 U206 ( .A(n243), .B(n142), .Y(n127) );
  INVX1 U207 ( .A(n154), .Y(n25) );
  NAND2X1 U208 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U209 ( .A(n138), .Y(n56) );
  NAND2X1 U210 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U211 ( .A(n64), .B(n124), .Y(n121) );
  AOI211X1 U212 ( .A0(n556), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  OAI2BB2X1 U213 ( .B0(n545), .B1(n183), .A0N(n188), .A1N(n540), .Y(n335) );
  AOI21X1 U214 ( .A0(n301), .A1(n337), .B0(n550), .Y(n336) );
  NAND2X1 U215 ( .A(n538), .B(n214), .Y(n126) );
  NAND2X1 U216 ( .A(n138), .B(n102), .Y(n227) );
  NAND2X1 U217 ( .A(n103), .B(n165), .Y(n188) );
  AOI21X1 U218 ( .A0(n556), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U219 ( .A0(n102), .A1(n103), .B0(n550), .Y(n101) );
  INVX1 U220 ( .A(n337), .Y(n65) );
  AOI22X1 U221 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  OAI221XL U222 ( .A0(n65), .A1(n551), .B0(n31), .B1(n536), .C0(n149), .Y(n143) );
  OAI221XL U223 ( .A0(n145), .A1(n545), .B0(n28), .B1(n551), .C0(n146), .Y(
        n144) );
  AOI2BB2X1 U224 ( .B0(n539), .B1(n87), .A0N(n545), .A1N(n121), .Y(n149) );
  INVX1 U225 ( .A(n208), .Y(n29) );
  INVX1 U226 ( .A(n299), .Y(n11) );
  INVX1 U227 ( .A(n100), .Y(n33) );
  AOI221XL U228 ( .A0(n556), .A1(n52), .B0(n548), .B1(n123), .C0(n324), .Y(
        n316) );
  INVX1 U229 ( .A(n326), .Y(n52) );
  OAI32X1 U230 ( .A0(n94), .A1(n63), .A2(n325), .B0(n37), .B1(n551), .Y(n324)
         );
  INVX1 U231 ( .A(n196), .Y(n31) );
  OAI221XL U232 ( .A0(n56), .A1(n545), .B0(n32), .B1(n543), .C0(n163), .Y(n151) );
  INVX1 U233 ( .A(n167), .Y(n32) );
  AOI22X1 U234 ( .A0(n164), .A1(n16), .B0(n129), .B1(n552), .Y(n163) );
  INVX1 U235 ( .A(n141), .Y(n27) );
  INVX1 U236 ( .A(n148), .Y(n28) );
  OAI221XL U237 ( .A0(n40), .A1(n551), .B0(n58), .B1(n545), .C0(n137), .Y(n136) );
  INVX1 U238 ( .A(n96), .Y(n40) );
  AOI31X1 U239 ( .A0(n102), .A1(n138), .A2(n556), .B0(n8), .Y(n137) );
  INVX1 U240 ( .A(n89), .Y(n8) );
  INVX1 U241 ( .A(n185), .Y(n19) );
  INVX1 U242 ( .A(n539), .Y(n543) );
  AOI211X1 U243 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U244 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI2BB2X1 U245 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  AOI211X1 U246 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U247 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U248 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  AOI22X1 U249 ( .A0(n533), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U250 ( .A0(n61), .A1(n551), .B0(n545), .B1(n260), .C0(n261), .Y(
        n254) );
  OAI221XL U251 ( .A0(n41), .A1(n545), .B0(n541), .B1(n181), .C0(n256), .Y(
        n255) );
  AOI21X1 U252 ( .A0(n33), .A1(n16), .B0(n262), .Y(n261) );
  AOI22X1 U253 ( .A0(n348), .A1(n26), .B0(n533), .B1(n349), .Y(n342) );
  OAI221XL U254 ( .A0(n536), .A1(n166), .B0(n286), .B1(n545), .C0(n351), .Y(
        n348) );
  OAI211X1 U255 ( .A0(n88), .A1(n550), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U256 ( .B0(n539), .B1(n196), .A0N(n550), .A1N(n179), .Y(n351) );
  OAI22X1 U257 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U258 ( .A0(n549), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U259 ( .A0(n56), .A1(n4), .B0(n547), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U260 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U261 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U262 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U263 ( .A0(n61), .A1(n554), .B0(n547), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U264 ( .A0(n541), .A1(n71), .B0(n37), .B1(n550), .Y(n157) );
  OAI22X1 U265 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U266 ( .A0(n549), .A1(n111), .B0(n47), .B1(n540), .C0(n112), .Y(
        n109) );
  AOI221X1 U267 ( .A0(n556), .A1(n115), .B0(n552), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U268 ( .A0(n536), .A1(n113), .B0(n44), .B1(n551), .C0(n114), .Y(
        n112) );
  AOI211X1 U269 ( .A0(n55), .A1(n556), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U270 ( .A0(n114), .A1(n206), .A2(n273), .B0(n533), .Y(n272) );
  OAI22X1 U271 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U272 ( .B0(n70), .B1(n552), .A0N(n90), .A1N(n545), .Y(n273) );
  AOI2BB2X1 U273 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  OAI221XL U274 ( .A0(n46), .A1(n551), .B0(n545), .B1(n116), .C0(n267), .Y(
        n264) );
  AOI221XL U275 ( .A0(n548), .A1(n247), .B0(n212), .B1(n540), .C0(n266), .Y(
        n265) );
  AOI22X1 U276 ( .A0(n539), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  AOI22X1 U277 ( .A0(n534), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U278 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  OAI221XL U279 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  AOI22X1 U281 ( .A0(n171), .A1(n21), .B0(n534), .B1(n172), .Y(n170) );
  OAI221XL U282 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  OAI221XL U283 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  AOI22X1 U284 ( .A0(n554), .A1(n532), .B0(n539), .B1(n66), .Y(n292) );
  AOI22X1 U285 ( .A0(n533), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U286 ( .A0(n43), .A1(n545), .B0(n94), .B1(n34), .C0(n365), .Y(n361)
         );
  OAI221XL U287 ( .A0(n532), .A1(n120), .B0(n201), .B1(n551), .C0(n363), .Y(
        n362) );
  INVX1 U288 ( .A(n260), .Y(n43) );
  AOI22X1 U289 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  OAI21XL U290 ( .A0(n321), .A1(n536), .B0(n322), .Y(n318) );
  OAI221XL U291 ( .A0(n551), .A1(n113), .B0(n88), .B1(n545), .C0(n320), .Y(
        n319) );
  AOI31X1 U292 ( .A0(n538), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  CLKINVX3 U293 ( .A(n532), .Y(n71) );
  OAI21XL U294 ( .A0(n545), .A1(n537), .B0(n120), .Y(n276) );
  NAND2X1 U295 ( .A(n63), .B(n531), .Y(n168) );
  AOI21X1 U296 ( .A0(n224), .A1(n243), .B0(n545), .Y(n295) );
  INVX1 U297 ( .A(n531), .Y(n74) );
  OAI21XL U298 ( .A0(n73), .A1(n301), .B0(n550), .Y(n323) );
  OAI21XL U299 ( .A0(n536), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U300 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U301 ( .A(n162), .Y(n5) );
  OAI2BB1X1 U302 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI22X1 U303 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  AOI211X1 U304 ( .A0(n39), .A1(n540), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U305 ( .A0(n551), .A1(n116), .B0(n73), .B1(n230), .C0(n545), .C1(
        n102), .Y(n275) );
  NAND2X1 U306 ( .A(n62), .B(n552), .Y(n287) );
  OAI2BB1X1 U307 ( .A0N(n133), .A1N(n134), .B0(n534), .Y(n132) );
  AOI22X1 U308 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  NOR2BX1 U309 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U310 ( .A(n82), .Y(n536) );
  NAND2X1 U311 ( .A(n73), .B(n20), .Y(n82) );
  OAI221XL U312 ( .A0(n531), .A1(n259), .B0(n542), .B1(n214), .C0(n287), .Y(
        n293) );
  BUFX3 U313 ( .A(n139), .Y(n538) );
  NAND2X1 U314 ( .A(n531), .B(n537), .Y(n139) );
  AOI211X1 U315 ( .A0(n540), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  OAI222X1 U316 ( .A0(n551), .A1(n167), .B0(n339), .B1(n536), .C0(n545), .C1(
        n34), .Y(n338) );
  AOI21X1 U317 ( .A0(n537), .A1(n535), .B0(n65), .Y(n339) );
  AOI211X1 U318 ( .A0(n533), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  OAI221XL U319 ( .A0(n545), .A1(n116), .B0(n321), .B1(n542), .C0(n359), .Y(
        n354) );
  AOI21X1 U320 ( .A0(n356), .A1(n357), .B0(n533), .Y(n355) );
  AOI31X1 U321 ( .A0(n556), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  INVX1 U322 ( .A(n93), .Y(n546) );
  INVX1 U323 ( .A(n83), .Y(n554) );
  INVX1 U324 ( .A(n83), .Y(n555) );
  INVX1 U325 ( .A(n544), .Y(n541) );
  INVX1 U326 ( .A(n94), .Y(n544) );
  AOI22X1 U327 ( .A0(n533), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U328 ( .A0(n545), .A1(n141), .B0(n551), .B1(n263), .C0(n29), .C1(
        n541), .Y(n277) );
  OAI221XL U329 ( .A0(n31), .A1(n536), .B0(n551), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U330 ( .B0(n88), .B1(n539), .A0N(n545), .A1N(n197), .Y(n279) );
  NAND2X1 U331 ( .A(n224), .B(n301), .Y(n148) );
  NOR2BX1 U332 ( .AN(n263), .B(n61), .Y(n321) );
  AOI21X1 U333 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI22X1 U334 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U335 ( .A0(n63), .A1(n545), .B0(n543), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U336 ( .A0(n38), .A1(n536), .B0(n545), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U337 ( .A0(n179), .A1(n552), .B0(n180), .Y(n178) );
  AOI22X1 U338 ( .A0(n556), .A1(n66), .B0(n539), .B1(n147), .Y(n146) );
  AOI22X1 U339 ( .A0(n549), .A1(n85), .B0(n41), .B1(n539), .Y(n84) );
  AOI31X1 U340 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U341 ( .A0N(n223), .A1N(n224), .B0(n553), .Y(n220) );
  AOI22X1 U342 ( .A0(n29), .A1(n556), .B0(n222), .B1(n547), .Y(n221) );
  NAND2X1 U343 ( .A(n224), .B(n118), .Y(n208) );
  NAND2X1 U344 ( .A(n263), .B(n337), .Y(n167) );
  AOI21X1 U345 ( .A0(n263), .A1(n182), .B0(n545), .Y(n305) );
  AOI21X1 U346 ( .A0(n111), .A1(n538), .B0(n542), .Y(n203) );
  NAND2X1 U347 ( .A(n16), .B(n531), .Y(n206) );
  OAI21XL U348 ( .A0(n73), .A1(n243), .B0(n550), .Y(n245) );
  XNOR2X1 U349 ( .A(n20), .B(n531), .Y(n185) );
  NAND2X1 U350 ( .A(n539), .B(n537), .Y(n130) );
  XNOR2X1 U351 ( .A(n73), .B(n531), .Y(n161) );
  AOI21X1 U352 ( .A0(n90), .A1(n73), .B0(n556), .Y(n86) );
  AOI221X1 U353 ( .A0(n46), .A1(n540), .B0(n553), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U354 ( .A0(n536), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U355 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  AOI222X1 U356 ( .A0(n549), .A1(n210), .B0(n211), .B1(n212), .C0(n556), .C1(
        n537), .Y(n191) );
  OAI21XL U357 ( .A0(n73), .A1(n214), .B0(n550), .Y(n211) );
  AOI31X1 U358 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U359 ( .A0(n148), .A1(n73), .B0(n29), .B1(n553), .Y(n300) );
  INVX1 U360 ( .A(n93), .Y(n547) );
  INVX1 U361 ( .A(n93), .Y(n549) );
  INVX1 U362 ( .A(n93), .Y(n548) );
  XOR2X1 U363 ( .A(n533), .B(n531), .Y(n358) );
  INVX1 U364 ( .A(n83), .Y(n552) );
  INVX1 U365 ( .A(n83), .Y(n553) );
  NOR2BX1 U366 ( .AN(n93), .B(n554), .Y(n309) );
  AOI22X1 U367 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U368 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI22X1 U369 ( .A0(n347), .A1(n26), .B0(n556), .B1(n90), .Y(n343) );
  AOI22X1 U370 ( .A0(n250), .A1(n21), .B0(n534), .B1(n251), .Y(n249) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  OAI22X1 U373 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U374 ( .A0(n548), .A1(n230), .B0(n556), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U375 ( .A0(n164), .A1(n547), .B0(a[2]), .B1(n227), .C0(n556), .C1(
        n228), .Y(n226) );
  OAI22X1 U376 ( .A0(n35), .A1(n543), .B0(n550), .B1(n537), .Y(n231) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI21XL U383 ( .A0(n66), .A1(n550), .B0(n259), .Y(n257) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI22X1 U385 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U386 ( .A(a[0]), .Y(n75) );
  AOI211X1 U387 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U388 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U389 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U390 ( .A(a[5]), .Y(n533) );
  OAI221XL U391 ( .A0(n536), .A1(n115), .B0(n121), .B1(n545), .C0(n122), .Y(
        n105) );
  AOI22X1 U392 ( .A0(n539), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  AOI33X1 U393 ( .A0(n532), .A1(n540), .A2(n19), .B0(n185), .B1(n181), .B2(
        a[2]), .Y(n184) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_15 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556;

  OAI221X4 U4 ( .A0(n66), .A1(n536), .B0(n61), .B1(n551), .C0(n84), .Y(n81) );
  OAI221X4 U6 ( .A0(n86), .A1(n87), .B0(n88), .B1(n551), .C0(n89), .Y(n80) );
  OAI222X4 U75 ( .A0(n551), .A1(n207), .B0(n181), .B1(n120), .C0(n545), .C1(
        n208), .Y(n204) );
  OAI32X4 U280 ( .A0(n551), .A1(n56), .A2(n53), .B0(n94), .B1(n103), .Y(n366)
         );
  AOI221X1 U1 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n103) );
  OAI222X1 U5 ( .A0(n94), .A1(n118), .B0(n119), .B1(n545), .C0(a[4]), .C1(n120), .Y(n117) );
  NAND2X2 U7 ( .A(n531), .B(n532), .Y(n115) );
  NAND2X1 U8 ( .A(n56), .B(n531), .Y(n229) );
  NAND2X2 U9 ( .A(n532), .B(n66), .Y(n181) );
  NAND2X1 U10 ( .A(n39), .B(n531), .Y(n142) );
  NAND2X2 U11 ( .A(n537), .B(n181), .Y(n113) );
  NAND2X2 U12 ( .A(n66), .B(n535), .Y(n116) );
  NAND2X2 U13 ( .A(n66), .B(n71), .Y(n138) );
  NAND2X1 U14 ( .A(n531), .B(n181), .Y(n102) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n73) );
  NAND2X1 U16 ( .A(n533), .B(n75), .Y(n110) );
  CLKINVX3 U17 ( .A(n533), .Y(n26) );
  NAND2X2 U18 ( .A(n75), .B(n26), .Y(n154) );
  NAND2X2 U19 ( .A(a[0]), .B(n26), .Y(n156) );
  CLKINVX3 U20 ( .A(n534), .Y(n21) );
  OAI22X2 U21 ( .A0(n340), .A1(n21), .B0(n534), .B1(n341), .Y(d[0]) );
  OAI22X2 U22 ( .A0(n534), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  INVX1 U23 ( .A(n249), .Y(d[3]) );
  OAI21X2 U24 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  AOI221X1 U25 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76) );
  OAI22X2 U26 ( .A0(n534), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  OAI21X2 U27 ( .A0(n534), .A1(n131), .B0(n132), .Y(d[6]) );
  AOI221X1 U28 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131)
         );
  NAND2X1 U29 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U30 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI21XL U31 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  NAND2X1 U32 ( .A(a[4]), .B(n535), .Y(n263) );
  NAND2X1 U33 ( .A(n531), .B(a[4]), .Y(n224) );
  NAND2X2 U34 ( .A(n532), .B(a[4]), .Y(n111) );
  CLKINVX3 U35 ( .A(a[4]), .Y(n66) );
  NAND2X1 U36 ( .A(n53), .B(n16), .Y(n288) );
  CLKINVX3 U37 ( .A(n542), .Y(n540) );
  INVX1 U38 ( .A(n325), .Y(n34) );
  NAND2X1 U39 ( .A(n113), .B(n535), .Y(n214) );
  NAND2X1 U40 ( .A(n56), .B(n535), .Y(n233) );
  NAND2X1 U41 ( .A(n46), .B(n535), .Y(n209) );
  NAND2X1 U42 ( .A(n50), .B(n535), .Y(n301) );
  NAND2X1 U43 ( .A(n538), .B(n268), .Y(n212) );
  NAND2X1 U44 ( .A(n147), .B(n214), .Y(n207) );
  NAND2X1 U45 ( .A(n115), .B(n209), .Y(n210) );
  INVX1 U46 ( .A(n168), .Y(n62) );
  INVX1 U47 ( .A(n538), .Y(n53) );
  INVX1 U48 ( .A(n182), .Y(n57) );
  NOR2X1 U49 ( .A(n535), .B(n39), .Y(n325) );
  CLKINVX3 U50 ( .A(n555), .Y(n550) );
  NAND2X1 U51 ( .A(n535), .B(n71), .Y(n118) );
  NAND2X1 U52 ( .A(n138), .B(n535), .Y(n223) );
  NAND2X1 U53 ( .A(n39), .B(n535), .Y(n248) );
  NAND2X1 U54 ( .A(n181), .B(n535), .Y(n166) );
  NAND2X1 U55 ( .A(n229), .B(n248), .Y(n87) );
  INVX1 U56 ( .A(n102), .Y(n61) );
  NAND2X1 U57 ( .A(n115), .B(n223), .Y(n306) );
  INVX1 U58 ( .A(n230), .Y(n69) );
  INVX1 U59 ( .A(n116), .Y(n64) );
  INVX1 U60 ( .A(n103), .Y(n68) );
  BUFX3 U61 ( .A(n74), .Y(n535) );
  NAND2X1 U62 ( .A(n50), .B(n531), .Y(n147) );
  NAND2X1 U63 ( .A(n531), .B(n539), .Y(n120) );
  NAND2X1 U64 ( .A(n111), .B(n535), .Y(n268) );
  NAND2X1 U65 ( .A(n531), .B(n113), .Y(n165) );
  NAND2X1 U66 ( .A(n531), .B(n138), .Y(n182) );
  INVX1 U67 ( .A(n312), .Y(d[1]) );
  INVX1 U68 ( .A(n170), .Y(d[5]) );
  INVX1 U69 ( .A(n537), .Y(n46) );
  NAND2X1 U70 ( .A(n16), .B(n532), .Y(n259) );
  NAND2X1 U71 ( .A(n111), .B(n147), .Y(n96) );
  NOR2X1 U72 ( .A(n537), .B(n535), .Y(n124) );
  CLKINVX3 U73 ( .A(n111), .Y(n39) );
  NAND2X1 U74 ( .A(n531), .B(n71), .Y(n230) );
  NAND2X1 U76 ( .A(n531), .B(n66), .Y(n337) );
  NAND2BX1 U77 ( .AN(n124), .B(n263), .Y(n196) );
  INVX1 U78 ( .A(n156), .Y(n24) );
  NAND2X1 U79 ( .A(n224), .B(n268), .Y(n141) );
  NAND2BX1 U80 ( .AN(n93), .B(n537), .Y(n299) );
  NAND2X1 U81 ( .A(n224), .B(n233), .Y(n104) );
  NAND2X1 U82 ( .A(n263), .B(n142), .Y(n100) );
  CLKINVX3 U83 ( .A(n108), .Y(n22) );
  BUFX3 U84 ( .A(a[1]), .Y(n531) );
  NAND2X1 U85 ( .A(a[7]), .B(a[2]), .Y(n94) );
  NAND2X1 U86 ( .A(n533), .B(a[0]), .Y(n108) );
  INVX1 U87 ( .A(n238), .Y(n15) );
  NAND2X1 U88 ( .A(n59), .B(n540), .Y(n114) );
  NAND2X1 U89 ( .A(n51), .B(n556), .Y(n238) );
  INVX1 U90 ( .A(n288), .Y(n14) );
  NOR2X1 U91 ( .A(n550), .B(n325), .Y(n199) );
  NOR2X1 U92 ( .A(n49), .B(n62), .Y(n247) );
  NAND2X1 U93 ( .A(n222), .B(n540), .Y(n162) );
  INVX1 U94 ( .A(n301), .Y(n49) );
  INVX1 U95 ( .A(n166), .Y(n60) );
  INVX1 U96 ( .A(n207), .Y(n48) );
  INVX1 U97 ( .A(n228), .Y(n51) );
  INVX4 U98 ( .A(n536), .Y(n556) );
  NOR2BX1 U99 ( .AN(n214), .B(n69), .Y(n88) );
  NOR2X1 U100 ( .A(n53), .B(n70), .Y(n326) );
  NOR2X1 U101 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U102 ( .A(n34), .B(n223), .Y(n183) );
  INVX1 U103 ( .A(n118), .Y(n70) );
  NAND2X1 U104 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U105 ( .A(n233), .Y(n55) );
  INVX1 U106 ( .A(n223), .Y(n59) );
  NOR2X1 U107 ( .A(n57), .B(n55), .Y(n197) );
  INVX1 U108 ( .A(n248), .Y(n37) );
  OAI221XL U109 ( .A0(n58), .A1(n545), .B0(n98), .B1(n542), .C0(n18), .Y(n347)
         );
  INVX1 U110 ( .A(n199), .Y(n18) );
  INVX1 U111 ( .A(n127), .Y(n35) );
  NOR2X1 U112 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U113 ( .A(n212), .Y(n41) );
  NOR2X1 U114 ( .A(n62), .B(n55), .Y(n145) );
  INVX1 U115 ( .A(n306), .Y(n58) );
  INVX1 U116 ( .A(n158), .Y(n42) );
  INVX1 U117 ( .A(n87), .Y(n38) );
  INVX1 U118 ( .A(n210), .Y(n44) );
  NAND2X1 U119 ( .A(n63), .B(n535), .Y(n243) );
  OAI22X1 U120 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U121 ( .A0(n61), .A1(n547), .B0(n556), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U122 ( .A0(n556), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U123 ( .A(n116), .B(n229), .Y(n244) );
  NOR2X1 U124 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U125 ( .A0(n542), .A1(n207), .B0(n545), .B1(n538), .Y(n242) );
  CLKINVX3 U126 ( .A(n113), .Y(n50) );
  CLKINVX3 U127 ( .A(n181), .Y(n63) );
  AOI22X1 U128 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U129 ( .A0(n98), .A1(n545), .B0(n30), .B1(n543), .C0(n99), .Y(n91)
         );
  OAI221XL U130 ( .A0(n42), .A1(n545), .B0(n51), .B1(n543), .C0(n95), .Y(n92)
         );
  INVX1 U131 ( .A(n104), .Y(n30) );
  NAND2X1 U132 ( .A(n556), .B(n96), .Y(n187) );
  NAND2X1 U133 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U134 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  OAI221XL U135 ( .A0(n46), .A1(n551), .B0(n63), .B1(n545), .C0(n200), .Y(n194) );
  OAI221XL U136 ( .A0(n536), .A1(n196), .B0(n197), .B1(n545), .C0(n198), .Y(
        n195) );
  AOI211X1 U137 ( .A0(n201), .A1(n556), .B0(n202), .C0(n203), .Y(n200) );
  AOI22X1 U138 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U139 ( .A0(n35), .A1(n545), .B0(n44), .B1(n543), .C0(n333), .Y(n332) );
  OAI211X1 U140 ( .A0(n326), .A1(n550), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U141 ( .A0(n35), .A1(n556), .B0(n39), .B1(n554), .Y(n333) );
  AOI22X1 U142 ( .A0(n548), .A1(n63), .B0(n247), .B1(n539), .Y(n334) );
  AOI21X1 U143 ( .A0(n115), .A1(n243), .B0(n550), .Y(n360) );
  INVX1 U144 ( .A(n120), .Y(n4) );
  AND2X2 U145 ( .A(n165), .B(n166), .Y(n129) );
  OAI21XL U146 ( .A0(n165), .A1(n550), .B0(n187), .Y(n266) );
  INVX1 U147 ( .A(n284), .Y(n10) );
  OAI31X1 U148 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U149 ( .A0(n541), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U150 ( .A(n147), .Y(n47) );
  OAI22X1 U151 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U152 ( .A0(n556), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U153 ( .A0(n11), .A1(n535), .B0(n27), .B1(n556), .C0(n307), .Y(n302) );
  OAI22X1 U154 ( .A0(n64), .A1(n543), .B0(n550), .B1(n306), .Y(n304) );
  AOI222X1 U155 ( .A0(n56), .A1(n540), .B0(n60), .B1(n554), .C0(n549), .C1(n71), .Y(n356) );
  AOI21X1 U156 ( .A0(n50), .A1(n556), .B0(n366), .Y(n365) );
  OAI221XL U157 ( .A0(n551), .A1(n87), .B0(n94), .B1(n104), .C0(n246), .Y(n235) );
  AOI2BB2X1 U158 ( .B0(n11), .B1(n535), .A0N(n536), .A1N(n247), .Y(n246) );
  CLKINVX8 U159 ( .A(n546), .Y(n545) );
  CLKINVX3 U160 ( .A(n541), .Y(n539) );
  NOR2X1 U161 ( .A(n545), .B(n535), .Y(n202) );
  AOI211X1 U162 ( .A0(n45), .A1(n540), .B0(n204), .C0(n205), .Y(n192) );
  INVX1 U163 ( .A(n209), .Y(n45) );
  NAND2BX1 U164 ( .AN(n97), .B(n206), .Y(n205) );
  AOI222X1 U165 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n540), 
        .Y(n198) );
  AOI221X1 U166 ( .A0(n321), .A1(n553), .B0(n540), .B1(n311), .C0(n327), .Y(
        n315) );
  OAI221XL U167 ( .A0(n536), .A1(n209), .B0(n545), .B1(n103), .C0(n288), .Y(
        n327) );
  AOI221X1 U168 ( .A0(n4), .A1(n71), .B0(n553), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI2BB1X1 U169 ( .A0N(n142), .A1N(n547), .B0(n187), .Y(n186) );
  OAI221XL U170 ( .A0(n308), .A1(n551), .B0(n545), .B1(n165), .C0(n162), .Y(
        n307) );
  NOR2X1 U171 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U172 ( .A0(n54), .A1(n545), .B0(n33), .B1(n543), .C0(n232), .Y(n217) );
  INVX1 U173 ( .A(n234), .Y(n54) );
  AOI32X1 U174 ( .A0(n34), .A1(n181), .A2(n556), .B0(n553), .B1(n233), .Y(n232) );
  OAI221XL U175 ( .A0(n67), .A1(n551), .B0(n94), .B1(n538), .C0(n294), .Y(n282) );
  INVX1 U176 ( .A(n115), .Y(n67) );
  AOI211X1 U177 ( .A0(n48), .A1(n556), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U178 ( .A(n114), .Y(n6) );
  AOI211X1 U179 ( .A0(n60), .A1(n540), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U180 ( .A(n545), .B(n39), .C(n61), .Y(n364) );
  INVX1 U181 ( .A(n259), .Y(n13) );
  OAI221XL U182 ( .A0(n536), .A1(n168), .B0(n164), .B1(n551), .C0(n169), .Y(
        n150) );
  AOI22X1 U183 ( .A0(n549), .A1(n34), .B0(n48), .B1(n539), .Y(n169) );
  AOI211X1 U184 ( .A0(n554), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  CLKINVX3 U185 ( .A(n555), .Y(n551) );
  INVX1 U186 ( .A(n544), .Y(n542) );
  INVX1 U187 ( .A(n125), .Y(n7) );
  AOI221X1 U188 ( .A0(n126), .A1(n552), .B0(n127), .B1(n548), .C0(n128), .Y(
        n125) );
  OAI21XL U189 ( .A0(n536), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U190 ( .A(n536), .Y(n16) );
  NOR2X1 U191 ( .A(n39), .B(n57), .Y(n179) );
  CLKINVX3 U192 ( .A(n110), .Y(n23) );
  NAND3X1 U193 ( .A(n538), .B(n113), .C(n540), .Y(n89) );
  NAND2X1 U194 ( .A(n214), .B(n142), .Y(n90) );
  NAND2X1 U195 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U196 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U197 ( .A(n538), .B(n166), .Y(n311) );
  NOR2BX1 U198 ( .AN(n229), .B(n68), .Y(n164) );
  AOI21X1 U199 ( .A0(n181), .A1(n182), .B0(n536), .Y(n180) );
  OAI221XL U200 ( .A0(n36), .A1(n550), .B0(n121), .B1(n541), .C0(n140), .Y(
        n135) );
  INVX1 U201 ( .A(n85), .Y(n36) );
  AOI22X1 U202 ( .A0(n49), .A1(n548), .B0(n556), .B1(n141), .Y(n140) );
  AOI22X1 U203 ( .A0(n57), .A1(n546), .B0(n555), .B1(n113), .Y(n239) );
  AOI22X1 U204 ( .A0(n547), .A1(n311), .B0(n50), .B1(n539), .Y(n350) );
  NOR2X1 U205 ( .A(n138), .B(n536), .Y(n97) );
  NAND2X1 U206 ( .A(n243), .B(n142), .Y(n127) );
  INVX1 U207 ( .A(n154), .Y(n25) );
  NAND2X1 U208 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U209 ( .A(n138), .Y(n56) );
  NAND2X1 U210 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U211 ( .A(n64), .B(n124), .Y(n121) );
  AOI211X1 U212 ( .A0(n556), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  OAI2BB2X1 U213 ( .B0(n545), .B1(n183), .A0N(n188), .A1N(n540), .Y(n335) );
  AOI21X1 U214 ( .A0(n301), .A1(n337), .B0(n550), .Y(n336) );
  NAND2X1 U215 ( .A(n538), .B(n214), .Y(n126) );
  NAND2X1 U216 ( .A(n138), .B(n102), .Y(n227) );
  NAND2X1 U217 ( .A(n103), .B(n165), .Y(n188) );
  AOI21X1 U218 ( .A0(n556), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U219 ( .A0(n102), .A1(n103), .B0(n550), .Y(n101) );
  INVX1 U220 ( .A(n337), .Y(n65) );
  AOI22X1 U221 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  OAI221XL U222 ( .A0(n65), .A1(n551), .B0(n31), .B1(n536), .C0(n149), .Y(n143) );
  OAI221XL U223 ( .A0(n145), .A1(n545), .B0(n28), .B1(n551), .C0(n146), .Y(
        n144) );
  AOI2BB2X1 U224 ( .B0(n539), .B1(n87), .A0N(n545), .A1N(n121), .Y(n149) );
  INVX1 U225 ( .A(n208), .Y(n29) );
  INVX1 U226 ( .A(n299), .Y(n11) );
  INVX1 U227 ( .A(n100), .Y(n33) );
  AOI221XL U228 ( .A0(n556), .A1(n52), .B0(n548), .B1(n123), .C0(n324), .Y(
        n316) );
  INVX1 U229 ( .A(n326), .Y(n52) );
  OAI32X1 U230 ( .A0(n94), .A1(n63), .A2(n325), .B0(n37), .B1(n551), .Y(n324)
         );
  INVX1 U231 ( .A(n196), .Y(n31) );
  OAI221XL U232 ( .A0(n56), .A1(n545), .B0(n32), .B1(n543), .C0(n163), .Y(n151) );
  INVX1 U233 ( .A(n167), .Y(n32) );
  AOI22X1 U234 ( .A0(n164), .A1(n16), .B0(n129), .B1(n552), .Y(n163) );
  INVX1 U235 ( .A(n141), .Y(n27) );
  INVX1 U236 ( .A(n148), .Y(n28) );
  OAI221XL U237 ( .A0(n40), .A1(n551), .B0(n58), .B1(n545), .C0(n137), .Y(n136) );
  INVX1 U238 ( .A(n96), .Y(n40) );
  AOI31X1 U239 ( .A0(n102), .A1(n138), .A2(n556), .B0(n8), .Y(n137) );
  INVX1 U240 ( .A(n89), .Y(n8) );
  INVX1 U241 ( .A(n185), .Y(n19) );
  INVX1 U242 ( .A(n539), .Y(n543) );
  AOI211X1 U243 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U244 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI2BB2X1 U245 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  AOI211X1 U246 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U247 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U248 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  AOI22X1 U249 ( .A0(n533), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U250 ( .A0(n61), .A1(n551), .B0(n545), .B1(n260), .C0(n261), .Y(
        n254) );
  OAI221XL U251 ( .A0(n41), .A1(n545), .B0(n541), .B1(n181), .C0(n256), .Y(
        n255) );
  AOI21X1 U252 ( .A0(n33), .A1(n16), .B0(n262), .Y(n261) );
  AOI22X1 U253 ( .A0(n348), .A1(n26), .B0(n533), .B1(n349), .Y(n342) );
  OAI221XL U254 ( .A0(n536), .A1(n166), .B0(n286), .B1(n545), .C0(n351), .Y(
        n348) );
  OAI211X1 U255 ( .A0(n88), .A1(n550), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U256 ( .B0(n539), .B1(n196), .A0N(n550), .A1N(n179), .Y(n351) );
  OAI22X1 U257 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U258 ( .A0(n549), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U259 ( .A0(n56), .A1(n4), .B0(n547), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U260 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U261 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U262 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U263 ( .A0(n61), .A1(n554), .B0(n547), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U264 ( .A0(n541), .A1(n71), .B0(n37), .B1(n550), .Y(n157) );
  OAI22X1 U265 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U266 ( .A0(n549), .A1(n111), .B0(n47), .B1(n540), .C0(n112), .Y(
        n109) );
  AOI221X1 U267 ( .A0(n556), .A1(n115), .B0(n552), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U268 ( .A0(n536), .A1(n113), .B0(n44), .B1(n551), .C0(n114), .Y(
        n112) );
  AOI211X1 U269 ( .A0(n55), .A1(n556), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U270 ( .A0(n114), .A1(n206), .A2(n273), .B0(n533), .Y(n272) );
  OAI22X1 U271 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U272 ( .B0(n70), .B1(n552), .A0N(n90), .A1N(n545), .Y(n273) );
  AOI2BB2X1 U273 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  OAI221XL U274 ( .A0(n46), .A1(n551), .B0(n545), .B1(n116), .C0(n267), .Y(
        n264) );
  AOI221XL U275 ( .A0(n548), .A1(n247), .B0(n212), .B1(n540), .C0(n266), .Y(
        n265) );
  AOI22X1 U276 ( .A0(n539), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  AOI22X1 U277 ( .A0(n534), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U278 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  OAI221XL U279 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  AOI22X1 U281 ( .A0(n171), .A1(n21), .B0(n534), .B1(n172), .Y(n170) );
  OAI221XL U282 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  OAI221XL U283 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  AOI22X1 U284 ( .A0(n554), .A1(n532), .B0(n539), .B1(n66), .Y(n292) );
  AOI22X1 U285 ( .A0(n533), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U286 ( .A0(n43), .A1(n545), .B0(n94), .B1(n34), .C0(n365), .Y(n361)
         );
  OAI221XL U287 ( .A0(n532), .A1(n120), .B0(n201), .B1(n551), .C0(n363), .Y(
        n362) );
  INVX1 U288 ( .A(n260), .Y(n43) );
  AOI22X1 U289 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  OAI21XL U290 ( .A0(n321), .A1(n536), .B0(n322), .Y(n318) );
  OAI221XL U291 ( .A0(n551), .A1(n113), .B0(n88), .B1(n545), .C0(n320), .Y(
        n319) );
  AOI31X1 U292 ( .A0(n538), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  CLKINVX3 U293 ( .A(n532), .Y(n71) );
  OAI21XL U294 ( .A0(n545), .A1(n537), .B0(n120), .Y(n276) );
  NAND2X1 U295 ( .A(n63), .B(n531), .Y(n168) );
  AOI21X1 U296 ( .A0(n224), .A1(n243), .B0(n545), .Y(n295) );
  INVX1 U297 ( .A(n531), .Y(n74) );
  OAI21XL U298 ( .A0(n73), .A1(n301), .B0(n550), .Y(n323) );
  OAI21XL U299 ( .A0(n536), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U300 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U301 ( .A(n162), .Y(n5) );
  OAI2BB1X1 U302 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI22X1 U303 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  AOI211X1 U304 ( .A0(n39), .A1(n540), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U305 ( .A0(n551), .A1(n116), .B0(n73), .B1(n230), .C0(n545), .C1(
        n102), .Y(n275) );
  NAND2X1 U306 ( .A(n62), .B(n552), .Y(n287) );
  OAI2BB1X1 U307 ( .A0N(n133), .A1N(n134), .B0(n534), .Y(n132) );
  AOI22X1 U308 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  NOR2BX1 U309 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U310 ( .A(n82), .Y(n536) );
  NAND2X1 U311 ( .A(n73), .B(n20), .Y(n82) );
  OAI221XL U312 ( .A0(n531), .A1(n259), .B0(n542), .B1(n214), .C0(n287), .Y(
        n293) );
  BUFX3 U313 ( .A(n139), .Y(n538) );
  NAND2X1 U314 ( .A(n531), .B(n537), .Y(n139) );
  AOI211X1 U315 ( .A0(n540), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  OAI222X1 U316 ( .A0(n551), .A1(n167), .B0(n339), .B1(n536), .C0(n545), .C1(
        n34), .Y(n338) );
  AOI21X1 U317 ( .A0(n537), .A1(n535), .B0(n65), .Y(n339) );
  AOI211X1 U318 ( .A0(n533), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  OAI221XL U319 ( .A0(n545), .A1(n116), .B0(n321), .B1(n542), .C0(n359), .Y(
        n354) );
  AOI21X1 U320 ( .A0(n356), .A1(n357), .B0(n533), .Y(n355) );
  AOI31X1 U321 ( .A0(n556), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  INVX1 U322 ( .A(n93), .Y(n546) );
  INVX1 U323 ( .A(n83), .Y(n554) );
  INVX1 U324 ( .A(n83), .Y(n555) );
  INVX1 U325 ( .A(n544), .Y(n541) );
  INVX1 U326 ( .A(n94), .Y(n544) );
  AOI22X1 U327 ( .A0(n533), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U328 ( .A0(n545), .A1(n141), .B0(n551), .B1(n263), .C0(n29), .C1(
        n541), .Y(n277) );
  OAI221XL U329 ( .A0(n31), .A1(n536), .B0(n551), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U330 ( .B0(n88), .B1(n539), .A0N(n545), .A1N(n197), .Y(n279) );
  NAND2X1 U331 ( .A(n224), .B(n301), .Y(n148) );
  NOR2BX1 U332 ( .AN(n263), .B(n61), .Y(n321) );
  AOI21X1 U333 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI22X1 U334 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U335 ( .A0(n63), .A1(n545), .B0(n543), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U336 ( .A0(n38), .A1(n536), .B0(n545), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U337 ( .A0(n179), .A1(n552), .B0(n180), .Y(n178) );
  AOI22X1 U338 ( .A0(n556), .A1(n66), .B0(n539), .B1(n147), .Y(n146) );
  AOI22X1 U339 ( .A0(n549), .A1(n85), .B0(n41), .B1(n539), .Y(n84) );
  AOI31X1 U340 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U341 ( .A0N(n223), .A1N(n224), .B0(n553), .Y(n220) );
  AOI22X1 U342 ( .A0(n29), .A1(n556), .B0(n222), .B1(n547), .Y(n221) );
  NAND2X1 U343 ( .A(n224), .B(n118), .Y(n208) );
  NAND2X1 U344 ( .A(n263), .B(n337), .Y(n167) );
  AOI21X1 U345 ( .A0(n263), .A1(n182), .B0(n545), .Y(n305) );
  AOI21X1 U346 ( .A0(n111), .A1(n538), .B0(n542), .Y(n203) );
  NAND2X1 U347 ( .A(n16), .B(n531), .Y(n206) );
  OAI21XL U348 ( .A0(n73), .A1(n243), .B0(n550), .Y(n245) );
  XNOR2X1 U349 ( .A(n20), .B(n531), .Y(n185) );
  NAND2X1 U350 ( .A(n539), .B(n537), .Y(n130) );
  XNOR2X1 U351 ( .A(n73), .B(n531), .Y(n161) );
  AOI21X1 U352 ( .A0(n90), .A1(n73), .B0(n556), .Y(n86) );
  AOI221X1 U353 ( .A0(n46), .A1(n540), .B0(n553), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U354 ( .A0(n536), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U355 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  AOI222X1 U356 ( .A0(n549), .A1(n210), .B0(n211), .B1(n212), .C0(n556), .C1(
        n537), .Y(n191) );
  OAI21XL U357 ( .A0(n73), .A1(n214), .B0(n550), .Y(n211) );
  AOI31X1 U358 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U359 ( .A0(n148), .A1(n73), .B0(n29), .B1(n553), .Y(n300) );
  INVX1 U360 ( .A(n93), .Y(n547) );
  INVX1 U361 ( .A(n93), .Y(n549) );
  INVX1 U362 ( .A(n93), .Y(n548) );
  XOR2X1 U363 ( .A(n533), .B(n531), .Y(n358) );
  INVX1 U364 ( .A(n83), .Y(n552) );
  INVX1 U365 ( .A(n83), .Y(n553) );
  NOR2BX1 U366 ( .AN(n93), .B(n554), .Y(n309) );
  AOI22X1 U367 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U368 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI22X1 U369 ( .A0(n347), .A1(n26), .B0(n556), .B1(n90), .Y(n343) );
  AOI22X1 U370 ( .A0(n250), .A1(n21), .B0(n534), .B1(n251), .Y(n249) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  OAI22X1 U373 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U374 ( .A0(n548), .A1(n230), .B0(n556), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U375 ( .A0(n164), .A1(n547), .B0(a[2]), .B1(n227), .C0(n556), .C1(
        n228), .Y(n226) );
  OAI22X1 U376 ( .A0(n35), .A1(n543), .B0(n550), .B1(n537), .Y(n231) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI21XL U383 ( .A0(n66), .A1(n550), .B0(n259), .Y(n257) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI22X1 U385 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U386 ( .A(a[0]), .Y(n75) );
  AOI211X1 U387 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U388 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U389 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U390 ( .A(a[5]), .Y(n533) );
  OAI221XL U391 ( .A0(n536), .A1(n115), .B0(n121), .B1(n545), .C0(n122), .Y(
        n105) );
  AOI22X1 U392 ( .A0(n539), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  AOI33X1 U393 ( .A0(n532), .A1(n540), .A2(n19), .B0(n185), .B1(n181), .B2(
        a[2]), .Y(n184) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_13 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556;

  OAI221X4 U4 ( .A0(n66), .A1(n536), .B0(n61), .B1(n551), .C0(n84), .Y(n81) );
  OAI221X4 U6 ( .A0(n86), .A1(n87), .B0(n88), .B1(n551), .C0(n89), .Y(n80) );
  OAI222X4 U75 ( .A0(n551), .A1(n207), .B0(n181), .B1(n120), .C0(n545), .C1(
        n208), .Y(n204) );
  OAI32X4 U280 ( .A0(n551), .A1(n56), .A2(n53), .B0(n94), .B1(n103), .Y(n366)
         );
  AOI221X1 U1 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n103) );
  OAI222X1 U5 ( .A0(n94), .A1(n118), .B0(n119), .B1(n545), .C0(a[4]), .C1(n120), .Y(n117) );
  NAND2X2 U7 ( .A(n531), .B(n532), .Y(n115) );
  NAND2X1 U8 ( .A(n56), .B(n531), .Y(n229) );
  NAND2X2 U9 ( .A(n532), .B(n66), .Y(n181) );
  NAND2X1 U10 ( .A(n39), .B(n531), .Y(n142) );
  NAND2X2 U11 ( .A(n537), .B(n181), .Y(n113) );
  NAND2X2 U12 ( .A(n66), .B(n535), .Y(n116) );
  NAND2X2 U13 ( .A(n66), .B(n71), .Y(n138) );
  NAND2X1 U14 ( .A(n531), .B(n181), .Y(n102) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n73) );
  NAND2X1 U16 ( .A(n533), .B(n75), .Y(n110) );
  CLKINVX3 U17 ( .A(n533), .Y(n26) );
  NAND2X2 U18 ( .A(n75), .B(n26), .Y(n154) );
  NAND2X2 U19 ( .A(a[0]), .B(n26), .Y(n156) );
  CLKINVX3 U20 ( .A(n534), .Y(n21) );
  OAI22X2 U21 ( .A0(n340), .A1(n21), .B0(n534), .B1(n341), .Y(d[0]) );
  OAI22X2 U22 ( .A0(n534), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  INVX1 U23 ( .A(n249), .Y(d[3]) );
  OAI21X2 U24 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  AOI221X1 U25 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76) );
  OAI22X2 U26 ( .A0(n534), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  OAI21X2 U27 ( .A0(n534), .A1(n131), .B0(n132), .Y(d[6]) );
  AOI221X1 U28 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131)
         );
  NAND2X1 U29 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U30 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI21XL U31 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  NAND2X1 U32 ( .A(a[4]), .B(n535), .Y(n263) );
  NAND2X1 U33 ( .A(n531), .B(a[4]), .Y(n224) );
  NAND2X2 U34 ( .A(n532), .B(a[4]), .Y(n111) );
  CLKINVX3 U35 ( .A(a[4]), .Y(n66) );
  NAND2X1 U36 ( .A(n53), .B(n16), .Y(n288) );
  CLKINVX3 U37 ( .A(n542), .Y(n540) );
  INVX1 U38 ( .A(n325), .Y(n34) );
  NAND2X1 U39 ( .A(n113), .B(n535), .Y(n214) );
  NAND2X1 U40 ( .A(n56), .B(n535), .Y(n233) );
  NAND2X1 U41 ( .A(n46), .B(n535), .Y(n209) );
  NAND2X1 U42 ( .A(n50), .B(n535), .Y(n301) );
  NAND2X1 U43 ( .A(n538), .B(n268), .Y(n212) );
  NAND2X1 U44 ( .A(n147), .B(n214), .Y(n207) );
  NAND2X1 U45 ( .A(n115), .B(n209), .Y(n210) );
  INVX1 U46 ( .A(n168), .Y(n62) );
  INVX1 U47 ( .A(n538), .Y(n53) );
  INVX1 U48 ( .A(n182), .Y(n57) );
  NOR2X1 U49 ( .A(n535), .B(n39), .Y(n325) );
  CLKINVX3 U50 ( .A(n555), .Y(n550) );
  NAND2X1 U51 ( .A(n535), .B(n71), .Y(n118) );
  NAND2X1 U52 ( .A(n138), .B(n535), .Y(n223) );
  NAND2X1 U53 ( .A(n39), .B(n535), .Y(n248) );
  NAND2X1 U54 ( .A(n181), .B(n535), .Y(n166) );
  NAND2X1 U55 ( .A(n229), .B(n248), .Y(n87) );
  INVX1 U56 ( .A(n102), .Y(n61) );
  NAND2X1 U57 ( .A(n115), .B(n223), .Y(n306) );
  INVX1 U58 ( .A(n230), .Y(n69) );
  INVX1 U59 ( .A(n116), .Y(n64) );
  INVX1 U60 ( .A(n103), .Y(n68) );
  BUFX3 U61 ( .A(n74), .Y(n535) );
  NAND2X1 U62 ( .A(n50), .B(n531), .Y(n147) );
  NAND2X1 U63 ( .A(n531), .B(n539), .Y(n120) );
  NAND2X1 U64 ( .A(n111), .B(n535), .Y(n268) );
  NAND2X1 U65 ( .A(n531), .B(n113), .Y(n165) );
  NAND2X1 U66 ( .A(n531), .B(n138), .Y(n182) );
  INVX1 U67 ( .A(n312), .Y(d[1]) );
  INVX1 U68 ( .A(n170), .Y(d[5]) );
  INVX1 U69 ( .A(n537), .Y(n46) );
  NAND2X1 U70 ( .A(n16), .B(n532), .Y(n259) );
  NAND2X1 U71 ( .A(n111), .B(n147), .Y(n96) );
  NOR2X1 U72 ( .A(n537), .B(n535), .Y(n124) );
  CLKINVX3 U73 ( .A(n111), .Y(n39) );
  NAND2X1 U74 ( .A(n531), .B(n71), .Y(n230) );
  NAND2X1 U76 ( .A(n531), .B(n66), .Y(n337) );
  NAND2BX1 U77 ( .AN(n124), .B(n263), .Y(n196) );
  INVX1 U78 ( .A(n156), .Y(n24) );
  NAND2X1 U79 ( .A(n224), .B(n268), .Y(n141) );
  NAND2BX1 U80 ( .AN(n93), .B(n537), .Y(n299) );
  NAND2X1 U81 ( .A(n224), .B(n233), .Y(n104) );
  NAND2X1 U82 ( .A(n263), .B(n142), .Y(n100) );
  CLKINVX3 U83 ( .A(n108), .Y(n22) );
  BUFX3 U84 ( .A(a[1]), .Y(n531) );
  NAND2X1 U85 ( .A(a[7]), .B(a[2]), .Y(n94) );
  NAND2X1 U86 ( .A(n533), .B(a[0]), .Y(n108) );
  INVX1 U87 ( .A(n238), .Y(n15) );
  NAND2X1 U88 ( .A(n59), .B(n540), .Y(n114) );
  NAND2X1 U89 ( .A(n51), .B(n556), .Y(n238) );
  INVX1 U90 ( .A(n288), .Y(n14) );
  NOR2X1 U91 ( .A(n550), .B(n325), .Y(n199) );
  NOR2X1 U92 ( .A(n49), .B(n62), .Y(n247) );
  NAND2X1 U93 ( .A(n222), .B(n540), .Y(n162) );
  INVX1 U94 ( .A(n301), .Y(n49) );
  INVX1 U95 ( .A(n166), .Y(n60) );
  INVX1 U96 ( .A(n207), .Y(n48) );
  INVX1 U97 ( .A(n228), .Y(n51) );
  INVX4 U98 ( .A(n536), .Y(n556) );
  NOR2BX1 U99 ( .AN(n214), .B(n69), .Y(n88) );
  NOR2X1 U100 ( .A(n53), .B(n70), .Y(n326) );
  NOR2X1 U101 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U102 ( .A(n34), .B(n223), .Y(n183) );
  INVX1 U103 ( .A(n118), .Y(n70) );
  NAND2X1 U104 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U105 ( .A(n233), .Y(n55) );
  INVX1 U106 ( .A(n223), .Y(n59) );
  NOR2X1 U107 ( .A(n57), .B(n55), .Y(n197) );
  INVX1 U108 ( .A(n248), .Y(n37) );
  OAI221XL U109 ( .A0(n58), .A1(n545), .B0(n98), .B1(n542), .C0(n18), .Y(n347)
         );
  INVX1 U110 ( .A(n199), .Y(n18) );
  INVX1 U111 ( .A(n127), .Y(n35) );
  NOR2X1 U112 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U113 ( .A(n212), .Y(n41) );
  NOR2X1 U114 ( .A(n62), .B(n55), .Y(n145) );
  INVX1 U115 ( .A(n306), .Y(n58) );
  INVX1 U116 ( .A(n158), .Y(n42) );
  INVX1 U117 ( .A(n87), .Y(n38) );
  INVX1 U118 ( .A(n210), .Y(n44) );
  NAND2X1 U119 ( .A(n63), .B(n535), .Y(n243) );
  OAI22X1 U120 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U121 ( .A0(n61), .A1(n547), .B0(n556), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U122 ( .A0(n556), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U123 ( .A(n116), .B(n229), .Y(n244) );
  NOR2X1 U124 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U125 ( .A0(n542), .A1(n207), .B0(n545), .B1(n538), .Y(n242) );
  CLKINVX3 U126 ( .A(n113), .Y(n50) );
  CLKINVX3 U127 ( .A(n181), .Y(n63) );
  AOI22X1 U128 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U129 ( .A0(n98), .A1(n545), .B0(n30), .B1(n543), .C0(n99), .Y(n91)
         );
  OAI221XL U130 ( .A0(n42), .A1(n545), .B0(n51), .B1(n543), .C0(n95), .Y(n92)
         );
  INVX1 U131 ( .A(n104), .Y(n30) );
  NAND2X1 U132 ( .A(n556), .B(n96), .Y(n187) );
  NAND2X1 U133 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U134 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  OAI221XL U135 ( .A0(n46), .A1(n551), .B0(n63), .B1(n545), .C0(n200), .Y(n194) );
  OAI221XL U136 ( .A0(n536), .A1(n196), .B0(n197), .B1(n545), .C0(n198), .Y(
        n195) );
  AOI211X1 U137 ( .A0(n201), .A1(n556), .B0(n202), .C0(n203), .Y(n200) );
  AOI22X1 U138 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U139 ( .A0(n35), .A1(n545), .B0(n44), .B1(n543), .C0(n333), .Y(n332) );
  OAI211X1 U140 ( .A0(n326), .A1(n550), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U141 ( .A0(n35), .A1(n556), .B0(n39), .B1(n554), .Y(n333) );
  AOI22X1 U142 ( .A0(n548), .A1(n63), .B0(n247), .B1(n539), .Y(n334) );
  AOI21X1 U143 ( .A0(n115), .A1(n243), .B0(n550), .Y(n360) );
  INVX1 U144 ( .A(n120), .Y(n4) );
  AND2X2 U145 ( .A(n165), .B(n166), .Y(n129) );
  OAI21XL U146 ( .A0(n165), .A1(n550), .B0(n187), .Y(n266) );
  INVX1 U147 ( .A(n284), .Y(n10) );
  OAI31X1 U148 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U149 ( .A0(n541), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U150 ( .A(n147), .Y(n47) );
  OAI22X1 U151 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U152 ( .A0(n556), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U153 ( .A0(n11), .A1(n535), .B0(n27), .B1(n556), .C0(n307), .Y(n302) );
  OAI22X1 U154 ( .A0(n64), .A1(n543), .B0(n550), .B1(n306), .Y(n304) );
  AOI222X1 U155 ( .A0(n56), .A1(n540), .B0(n60), .B1(n554), .C0(n549), .C1(n71), .Y(n356) );
  AOI21X1 U156 ( .A0(n50), .A1(n556), .B0(n366), .Y(n365) );
  OAI221XL U157 ( .A0(n551), .A1(n87), .B0(n94), .B1(n104), .C0(n246), .Y(n235) );
  AOI2BB2X1 U158 ( .B0(n11), .B1(n535), .A0N(n536), .A1N(n247), .Y(n246) );
  CLKINVX8 U159 ( .A(n546), .Y(n545) );
  CLKINVX3 U160 ( .A(n541), .Y(n539) );
  NOR2X1 U161 ( .A(n545), .B(n535), .Y(n202) );
  AOI211X1 U162 ( .A0(n45), .A1(n540), .B0(n204), .C0(n205), .Y(n192) );
  INVX1 U163 ( .A(n209), .Y(n45) );
  NAND2BX1 U164 ( .AN(n97), .B(n206), .Y(n205) );
  AOI222X1 U165 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n540), 
        .Y(n198) );
  AOI221X1 U166 ( .A0(n321), .A1(n553), .B0(n540), .B1(n311), .C0(n327), .Y(
        n315) );
  OAI221XL U167 ( .A0(n536), .A1(n209), .B0(n545), .B1(n103), .C0(n288), .Y(
        n327) );
  AOI221X1 U168 ( .A0(n4), .A1(n71), .B0(n553), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI2BB1X1 U169 ( .A0N(n142), .A1N(n547), .B0(n187), .Y(n186) );
  OAI221XL U170 ( .A0(n308), .A1(n551), .B0(n545), .B1(n165), .C0(n162), .Y(
        n307) );
  NOR2X1 U171 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U172 ( .A0(n54), .A1(n545), .B0(n33), .B1(n543), .C0(n232), .Y(n217) );
  INVX1 U173 ( .A(n234), .Y(n54) );
  AOI32X1 U174 ( .A0(n34), .A1(n181), .A2(n556), .B0(n553), .B1(n233), .Y(n232) );
  OAI221XL U175 ( .A0(n67), .A1(n551), .B0(n94), .B1(n538), .C0(n294), .Y(n282) );
  INVX1 U176 ( .A(n115), .Y(n67) );
  AOI211X1 U177 ( .A0(n48), .A1(n556), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U178 ( .A(n114), .Y(n6) );
  AOI211X1 U179 ( .A0(n60), .A1(n540), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U180 ( .A(n545), .B(n39), .C(n61), .Y(n364) );
  INVX1 U181 ( .A(n259), .Y(n13) );
  OAI221XL U182 ( .A0(n536), .A1(n168), .B0(n164), .B1(n551), .C0(n169), .Y(
        n150) );
  AOI22X1 U183 ( .A0(n549), .A1(n34), .B0(n48), .B1(n539), .Y(n169) );
  AOI211X1 U184 ( .A0(n554), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  CLKINVX3 U185 ( .A(n555), .Y(n551) );
  INVX1 U186 ( .A(n544), .Y(n542) );
  INVX1 U187 ( .A(n125), .Y(n7) );
  AOI221X1 U188 ( .A0(n126), .A1(n552), .B0(n127), .B1(n548), .C0(n128), .Y(
        n125) );
  OAI21XL U189 ( .A0(n536), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U190 ( .A(n536), .Y(n16) );
  NOR2X1 U191 ( .A(n39), .B(n57), .Y(n179) );
  CLKINVX3 U192 ( .A(n110), .Y(n23) );
  NAND3X1 U193 ( .A(n538), .B(n113), .C(n540), .Y(n89) );
  NAND2X1 U194 ( .A(n214), .B(n142), .Y(n90) );
  NAND2X1 U195 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U196 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U197 ( .A(n538), .B(n166), .Y(n311) );
  NOR2BX1 U198 ( .AN(n229), .B(n68), .Y(n164) );
  AOI21X1 U199 ( .A0(n181), .A1(n182), .B0(n536), .Y(n180) );
  OAI221XL U200 ( .A0(n36), .A1(n550), .B0(n121), .B1(n541), .C0(n140), .Y(
        n135) );
  INVX1 U201 ( .A(n85), .Y(n36) );
  AOI22X1 U202 ( .A0(n49), .A1(n548), .B0(n556), .B1(n141), .Y(n140) );
  AOI22X1 U203 ( .A0(n57), .A1(n546), .B0(n555), .B1(n113), .Y(n239) );
  AOI22X1 U204 ( .A0(n547), .A1(n311), .B0(n50), .B1(n539), .Y(n350) );
  NOR2X1 U205 ( .A(n138), .B(n536), .Y(n97) );
  NAND2X1 U206 ( .A(n243), .B(n142), .Y(n127) );
  INVX1 U207 ( .A(n154), .Y(n25) );
  NAND2X1 U208 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U209 ( .A(n138), .Y(n56) );
  NAND2X1 U210 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U211 ( .A(n64), .B(n124), .Y(n121) );
  AOI211X1 U212 ( .A0(n556), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  OAI2BB2X1 U213 ( .B0(n545), .B1(n183), .A0N(n188), .A1N(n540), .Y(n335) );
  AOI21X1 U214 ( .A0(n301), .A1(n337), .B0(n550), .Y(n336) );
  NAND2X1 U215 ( .A(n538), .B(n214), .Y(n126) );
  NAND2X1 U216 ( .A(n138), .B(n102), .Y(n227) );
  NAND2X1 U217 ( .A(n103), .B(n165), .Y(n188) );
  AOI21X1 U218 ( .A0(n556), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U219 ( .A0(n102), .A1(n103), .B0(n550), .Y(n101) );
  INVX1 U220 ( .A(n337), .Y(n65) );
  AOI22X1 U221 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  OAI221XL U222 ( .A0(n65), .A1(n551), .B0(n31), .B1(n536), .C0(n149), .Y(n143) );
  OAI221XL U223 ( .A0(n145), .A1(n545), .B0(n28), .B1(n551), .C0(n146), .Y(
        n144) );
  AOI2BB2X1 U224 ( .B0(n539), .B1(n87), .A0N(n545), .A1N(n121), .Y(n149) );
  INVX1 U225 ( .A(n208), .Y(n29) );
  INVX1 U226 ( .A(n299), .Y(n11) );
  INVX1 U227 ( .A(n100), .Y(n33) );
  AOI221XL U228 ( .A0(n556), .A1(n52), .B0(n548), .B1(n123), .C0(n324), .Y(
        n316) );
  INVX1 U229 ( .A(n326), .Y(n52) );
  OAI32X1 U230 ( .A0(n94), .A1(n63), .A2(n325), .B0(n37), .B1(n551), .Y(n324)
         );
  INVX1 U231 ( .A(n196), .Y(n31) );
  OAI221XL U232 ( .A0(n56), .A1(n545), .B0(n32), .B1(n543), .C0(n163), .Y(n151) );
  INVX1 U233 ( .A(n167), .Y(n32) );
  AOI22X1 U234 ( .A0(n164), .A1(n16), .B0(n129), .B1(n552), .Y(n163) );
  INVX1 U235 ( .A(n141), .Y(n27) );
  INVX1 U236 ( .A(n148), .Y(n28) );
  OAI221XL U237 ( .A0(n40), .A1(n551), .B0(n58), .B1(n545), .C0(n137), .Y(n136) );
  INVX1 U238 ( .A(n96), .Y(n40) );
  AOI31X1 U239 ( .A0(n102), .A1(n138), .A2(n556), .B0(n8), .Y(n137) );
  INVX1 U240 ( .A(n89), .Y(n8) );
  INVX1 U241 ( .A(n185), .Y(n19) );
  INVX1 U242 ( .A(n539), .Y(n543) );
  AOI211X1 U243 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U244 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI2BB2X1 U245 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  AOI211X1 U246 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U247 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U248 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  AOI22X1 U249 ( .A0(n533), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U250 ( .A0(n61), .A1(n551), .B0(n545), .B1(n260), .C0(n261), .Y(
        n254) );
  OAI221XL U251 ( .A0(n41), .A1(n545), .B0(n541), .B1(n181), .C0(n256), .Y(
        n255) );
  AOI21X1 U252 ( .A0(n33), .A1(n16), .B0(n262), .Y(n261) );
  AOI22X1 U253 ( .A0(n348), .A1(n26), .B0(n533), .B1(n349), .Y(n342) );
  OAI221XL U254 ( .A0(n536), .A1(n166), .B0(n286), .B1(n545), .C0(n351), .Y(
        n348) );
  OAI211X1 U255 ( .A0(n88), .A1(n550), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U256 ( .B0(n539), .B1(n196), .A0N(n550), .A1N(n179), .Y(n351) );
  OAI22X1 U257 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U258 ( .A0(n549), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U259 ( .A0(n56), .A1(n4), .B0(n547), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U260 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U261 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U262 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U263 ( .A0(n61), .A1(n554), .B0(n547), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U264 ( .A0(n541), .A1(n71), .B0(n37), .B1(n550), .Y(n157) );
  OAI22X1 U265 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U266 ( .A0(n549), .A1(n111), .B0(n47), .B1(n540), .C0(n112), .Y(
        n109) );
  AOI221X1 U267 ( .A0(n556), .A1(n115), .B0(n552), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U268 ( .A0(n536), .A1(n113), .B0(n44), .B1(n551), .C0(n114), .Y(
        n112) );
  AOI211X1 U269 ( .A0(n55), .A1(n556), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U270 ( .A0(n114), .A1(n206), .A2(n273), .B0(n533), .Y(n272) );
  OAI22X1 U271 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U272 ( .B0(n70), .B1(n552), .A0N(n90), .A1N(n545), .Y(n273) );
  AOI2BB2X1 U273 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  OAI221XL U274 ( .A0(n46), .A1(n551), .B0(n545), .B1(n116), .C0(n267), .Y(
        n264) );
  AOI221XL U275 ( .A0(n548), .A1(n247), .B0(n212), .B1(n540), .C0(n266), .Y(
        n265) );
  AOI22X1 U276 ( .A0(n539), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  AOI22X1 U277 ( .A0(n534), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U278 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  OAI221XL U279 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  AOI22X1 U281 ( .A0(n171), .A1(n21), .B0(n534), .B1(n172), .Y(n170) );
  OAI221XL U282 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  OAI221XL U283 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  AOI22X1 U284 ( .A0(n554), .A1(n532), .B0(n539), .B1(n66), .Y(n292) );
  AOI22X1 U285 ( .A0(n533), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U286 ( .A0(n43), .A1(n545), .B0(n94), .B1(n34), .C0(n365), .Y(n361)
         );
  OAI221XL U287 ( .A0(n532), .A1(n120), .B0(n201), .B1(n551), .C0(n363), .Y(
        n362) );
  INVX1 U288 ( .A(n260), .Y(n43) );
  AOI22X1 U289 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  OAI21XL U290 ( .A0(n321), .A1(n536), .B0(n322), .Y(n318) );
  OAI221XL U291 ( .A0(n551), .A1(n113), .B0(n88), .B1(n545), .C0(n320), .Y(
        n319) );
  AOI31X1 U292 ( .A0(n538), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  CLKINVX3 U293 ( .A(n532), .Y(n71) );
  OAI21XL U294 ( .A0(n545), .A1(n537), .B0(n120), .Y(n276) );
  NAND2X1 U295 ( .A(n63), .B(n531), .Y(n168) );
  AOI21X1 U296 ( .A0(n224), .A1(n243), .B0(n545), .Y(n295) );
  INVX1 U297 ( .A(n531), .Y(n74) );
  OAI21XL U298 ( .A0(n73), .A1(n301), .B0(n550), .Y(n323) );
  OAI21XL U299 ( .A0(n536), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U300 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U301 ( .A(n162), .Y(n5) );
  OAI2BB1X1 U302 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI22X1 U303 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  AOI211X1 U304 ( .A0(n39), .A1(n540), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U305 ( .A0(n551), .A1(n116), .B0(n73), .B1(n230), .C0(n545), .C1(
        n102), .Y(n275) );
  NAND2X1 U306 ( .A(n62), .B(n552), .Y(n287) );
  OAI2BB1X1 U307 ( .A0N(n133), .A1N(n134), .B0(n534), .Y(n132) );
  AOI22X1 U308 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  NOR2BX1 U309 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U310 ( .A(n82), .Y(n536) );
  NAND2X1 U311 ( .A(n73), .B(n20), .Y(n82) );
  OAI221XL U312 ( .A0(n531), .A1(n259), .B0(n542), .B1(n214), .C0(n287), .Y(
        n293) );
  BUFX3 U313 ( .A(n139), .Y(n538) );
  NAND2X1 U314 ( .A(n531), .B(n537), .Y(n139) );
  AOI211X1 U315 ( .A0(n540), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  OAI222X1 U316 ( .A0(n551), .A1(n167), .B0(n339), .B1(n536), .C0(n545), .C1(
        n34), .Y(n338) );
  AOI21X1 U317 ( .A0(n537), .A1(n535), .B0(n65), .Y(n339) );
  AOI211X1 U318 ( .A0(n533), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  OAI221XL U319 ( .A0(n545), .A1(n116), .B0(n321), .B1(n542), .C0(n359), .Y(
        n354) );
  AOI21X1 U320 ( .A0(n356), .A1(n357), .B0(n533), .Y(n355) );
  AOI31X1 U321 ( .A0(n556), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  INVX1 U322 ( .A(n93), .Y(n546) );
  INVX1 U323 ( .A(n83), .Y(n554) );
  INVX1 U324 ( .A(n83), .Y(n555) );
  INVX1 U325 ( .A(n544), .Y(n541) );
  INVX1 U326 ( .A(n94), .Y(n544) );
  AOI22X1 U327 ( .A0(n533), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U328 ( .A0(n545), .A1(n141), .B0(n551), .B1(n263), .C0(n29), .C1(
        n541), .Y(n277) );
  OAI221XL U329 ( .A0(n31), .A1(n536), .B0(n551), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U330 ( .B0(n88), .B1(n539), .A0N(n545), .A1N(n197), .Y(n279) );
  NAND2X1 U331 ( .A(n224), .B(n301), .Y(n148) );
  NOR2BX1 U332 ( .AN(n263), .B(n61), .Y(n321) );
  AOI21X1 U333 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI22X1 U334 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U335 ( .A0(n63), .A1(n545), .B0(n543), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U336 ( .A0(n38), .A1(n536), .B0(n545), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U337 ( .A0(n179), .A1(n552), .B0(n180), .Y(n178) );
  AOI22X1 U338 ( .A0(n556), .A1(n66), .B0(n539), .B1(n147), .Y(n146) );
  AOI22X1 U339 ( .A0(n549), .A1(n85), .B0(n41), .B1(n539), .Y(n84) );
  AOI31X1 U340 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U341 ( .A0N(n223), .A1N(n224), .B0(n553), .Y(n220) );
  AOI22X1 U342 ( .A0(n29), .A1(n556), .B0(n222), .B1(n547), .Y(n221) );
  NAND2X1 U343 ( .A(n224), .B(n118), .Y(n208) );
  NAND2X1 U344 ( .A(n263), .B(n337), .Y(n167) );
  AOI21X1 U345 ( .A0(n263), .A1(n182), .B0(n545), .Y(n305) );
  AOI21X1 U346 ( .A0(n111), .A1(n538), .B0(n542), .Y(n203) );
  NAND2X1 U347 ( .A(n16), .B(n531), .Y(n206) );
  OAI21XL U348 ( .A0(n73), .A1(n243), .B0(n550), .Y(n245) );
  XNOR2X1 U349 ( .A(n20), .B(n531), .Y(n185) );
  NAND2X1 U350 ( .A(n539), .B(n537), .Y(n130) );
  XNOR2X1 U351 ( .A(n73), .B(n531), .Y(n161) );
  AOI21X1 U352 ( .A0(n90), .A1(n73), .B0(n556), .Y(n86) );
  AOI221X1 U353 ( .A0(n46), .A1(n540), .B0(n553), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U354 ( .A0(n536), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U355 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  AOI222X1 U356 ( .A0(n549), .A1(n210), .B0(n211), .B1(n212), .C0(n556), .C1(
        n537), .Y(n191) );
  OAI21XL U357 ( .A0(n73), .A1(n214), .B0(n550), .Y(n211) );
  AOI31X1 U358 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U359 ( .A0(n148), .A1(n73), .B0(n29), .B1(n553), .Y(n300) );
  INVX1 U360 ( .A(n93), .Y(n547) );
  INVX1 U361 ( .A(n93), .Y(n549) );
  INVX1 U362 ( .A(n93), .Y(n548) );
  XOR2X1 U363 ( .A(n533), .B(n531), .Y(n358) );
  INVX1 U364 ( .A(n83), .Y(n552) );
  INVX1 U365 ( .A(n83), .Y(n553) );
  NOR2BX1 U366 ( .AN(n93), .B(n554), .Y(n309) );
  AOI22X1 U367 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U368 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI22X1 U369 ( .A0(n347), .A1(n26), .B0(n556), .B1(n90), .Y(n343) );
  AOI22X1 U370 ( .A0(n250), .A1(n21), .B0(n534), .B1(n251), .Y(n249) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  OAI22X1 U373 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U374 ( .A0(n548), .A1(n230), .B0(n556), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U375 ( .A0(n164), .A1(n547), .B0(a[2]), .B1(n227), .C0(n556), .C1(
        n228), .Y(n226) );
  OAI22X1 U376 ( .A0(n35), .A1(n543), .B0(n550), .B1(n537), .Y(n231) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI21XL U383 ( .A0(n66), .A1(n550), .B0(n259), .Y(n257) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI22X1 U385 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U386 ( .A(a[0]), .Y(n75) );
  AOI211X1 U387 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U388 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U389 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U390 ( .A(a[5]), .Y(n533) );
  OAI221XL U391 ( .A0(n536), .A1(n115), .B0(n121), .B1(n545), .C0(n122), .Y(
        n105) );
  AOI22X1 U392 ( .A0(n539), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  AOI33X1 U393 ( .A0(n532), .A1(n540), .A2(n19), .B0(n185), .B1(n181), .B2(
        a[2]), .Y(n184) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_12 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556;

  OAI221X4 U4 ( .A0(n66), .A1(n536), .B0(n61), .B1(n551), .C0(n84), .Y(n81) );
  OAI221X4 U6 ( .A0(n86), .A1(n87), .B0(n88), .B1(n551), .C0(n89), .Y(n80) );
  OAI221X4 U28 ( .A0(n40), .A1(n551), .B0(n58), .B1(n545), .C0(n137), .Y(n136)
         );
  OAI221X4 U35 ( .A0(n145), .A1(n545), .B0(n28), .B1(n551), .C0(n146), .Y(n144) );
  OAI221X4 U70 ( .A0(n46), .A1(n551), .B0(n63), .B1(n545), .C0(n200), .Y(n194)
         );
  OAI221X4 U103 ( .A0(n551), .A1(n87), .B0(n94), .B1(n104), .C0(n246), .Y(n235) );
  OAI221X4 U151 ( .A0(n67), .A1(n551), .B0(n542), .B1(n538), .C0(n294), .Y(
        n282) );
  OAI221X4 U166 ( .A0(n308), .A1(n551), .B0(n545), .B1(n165), .C0(n162), .Y(
        n307) );
  OAI32X4 U280 ( .A0(n551), .A1(n56), .A2(n53), .B0(n542), .B1(n103), .Y(n366)
         );
  AOI221X1 U1 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n103) );
  NAND2X2 U5 ( .A(n531), .B(n532), .Y(n115) );
  NAND2X1 U7 ( .A(n56), .B(n531), .Y(n229) );
  NAND2X2 U8 ( .A(n532), .B(n66), .Y(n181) );
  NAND2X1 U9 ( .A(n531), .B(n539), .Y(n120) );
  NAND2X1 U10 ( .A(n39), .B(n531), .Y(n142) );
  NAND2X2 U11 ( .A(n537), .B(n181), .Y(n113) );
  NAND2X2 U12 ( .A(n66), .B(n535), .Y(n116) );
  NAND2X2 U13 ( .A(n66), .B(n71), .Y(n138) );
  NAND2X1 U14 ( .A(n531), .B(n181), .Y(n102) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n73) );
  NAND2X1 U16 ( .A(n533), .B(n75), .Y(n110) );
  CLKINVX3 U17 ( .A(n533), .Y(n26) );
  NAND2X2 U18 ( .A(n75), .B(n26), .Y(n154) );
  NAND2X2 U19 ( .A(a[0]), .B(n26), .Y(n156) );
  OAI22X2 U20 ( .A0(n534), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  OAI21X2 U21 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  AOI221X1 U22 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76) );
  OAI22X2 U23 ( .A0(n534), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  NAND2X1 U24 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U25 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI21XL U26 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  OAI222X4 U27 ( .A0(n541), .A1(n118), .B0(n119), .B1(n545), .C0(a[4]), .C1(
        n120), .Y(n117) );
  NAND2X1 U29 ( .A(n531), .B(a[4]), .Y(n224) );
  NAND2X1 U30 ( .A(a[4]), .B(n535), .Y(n263) );
  NAND2X2 U31 ( .A(n532), .B(a[4]), .Y(n111) );
  CLKINVX3 U32 ( .A(a[4]), .Y(n66) );
  NAND2X1 U33 ( .A(n53), .B(n16), .Y(n288) );
  CLKINVX3 U34 ( .A(n541), .Y(n540) );
  INVX1 U36 ( .A(n325), .Y(n34) );
  NAND2X1 U37 ( .A(n113), .B(n535), .Y(n214) );
  NAND2X1 U38 ( .A(n56), .B(n535), .Y(n233) );
  NAND2X1 U39 ( .A(n46), .B(n535), .Y(n209) );
  NAND2X1 U40 ( .A(n50), .B(n535), .Y(n301) );
  NAND2X1 U41 ( .A(n538), .B(n268), .Y(n212) );
  NAND2X1 U42 ( .A(n147), .B(n214), .Y(n207) );
  NAND2X1 U43 ( .A(n115), .B(n209), .Y(n210) );
  INVX1 U44 ( .A(n168), .Y(n62) );
  INVX1 U45 ( .A(n538), .Y(n53) );
  INVX1 U46 ( .A(n182), .Y(n57) );
  NOR2X1 U47 ( .A(n535), .B(n39), .Y(n325) );
  CLKINVX3 U48 ( .A(n555), .Y(n550) );
  NAND2X1 U49 ( .A(n535), .B(n71), .Y(n118) );
  NAND2X1 U50 ( .A(n138), .B(n535), .Y(n223) );
  NAND2X1 U51 ( .A(n39), .B(n535), .Y(n248) );
  NAND2X1 U52 ( .A(n181), .B(n535), .Y(n166) );
  NAND2X1 U53 ( .A(n229), .B(n248), .Y(n87) );
  CLKINVX3 U54 ( .A(n110), .Y(n23) );
  INVX1 U55 ( .A(n102), .Y(n61) );
  NAND2X1 U56 ( .A(n115), .B(n223), .Y(n306) );
  INVX1 U57 ( .A(n230), .Y(n69) );
  INVX1 U58 ( .A(n116), .Y(n64) );
  INVX1 U59 ( .A(n103), .Y(n68) );
  BUFX3 U60 ( .A(n74), .Y(n535) );
  NAND2X1 U61 ( .A(n50), .B(n531), .Y(n147) );
  NAND2X1 U62 ( .A(n111), .B(n535), .Y(n268) );
  NAND2X1 U63 ( .A(n531), .B(n113), .Y(n165) );
  NAND2X1 U64 ( .A(n531), .B(n138), .Y(n182) );
  INVX1 U65 ( .A(n537), .Y(n46) );
  NAND2X1 U66 ( .A(n16), .B(n532), .Y(n259) );
  NAND2X1 U67 ( .A(n111), .B(n147), .Y(n96) );
  NOR2X1 U68 ( .A(n537), .B(n535), .Y(n124) );
  CLKINVX3 U69 ( .A(n111), .Y(n39) );
  NAND2X1 U71 ( .A(n531), .B(n71), .Y(n230) );
  NAND2X1 U72 ( .A(n531), .B(n66), .Y(n337) );
  NAND2BX1 U73 ( .AN(n124), .B(n263), .Y(n196) );
  INVX1 U74 ( .A(n156), .Y(n24) );
  NAND2X1 U75 ( .A(n224), .B(n268), .Y(n141) );
  NAND2BX1 U76 ( .AN(n93), .B(n537), .Y(n299) );
  NAND2X1 U77 ( .A(n224), .B(n233), .Y(n104) );
  NAND2X1 U78 ( .A(n263), .B(n142), .Y(n100) );
  CLKINVX3 U79 ( .A(n534), .Y(n21) );
  CLKINVX3 U80 ( .A(n108), .Y(n22) );
  INVX1 U81 ( .A(n249), .Y(d[3]) );
  BUFX3 U82 ( .A(a[1]), .Y(n531) );
  NAND2X1 U83 ( .A(a[7]), .B(a[2]), .Y(n94) );
  NAND2X1 U84 ( .A(n533), .B(a[0]), .Y(n108) );
  INVX1 U85 ( .A(n238), .Y(n15) );
  NAND2X1 U86 ( .A(n59), .B(n540), .Y(n114) );
  NAND2X1 U87 ( .A(n51), .B(n556), .Y(n238) );
  INVX1 U88 ( .A(n288), .Y(n14) );
  NOR2X1 U89 ( .A(n550), .B(n325), .Y(n199) );
  NOR2X1 U90 ( .A(n49), .B(n62), .Y(n247) );
  NAND2X1 U91 ( .A(n222), .B(n540), .Y(n162) );
  INVX1 U92 ( .A(n301), .Y(n49) );
  INVX1 U93 ( .A(n248), .Y(n37) );
  INVX1 U94 ( .A(n166), .Y(n60) );
  INVX1 U95 ( .A(n207), .Y(n48) );
  INVX1 U96 ( .A(n228), .Y(n51) );
  INVX4 U97 ( .A(n536), .Y(n556) );
  NOR2BX1 U98 ( .AN(n214), .B(n69), .Y(n88) );
  NOR2X1 U99 ( .A(n53), .B(n70), .Y(n326) );
  AOI22X1 U100 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  OAI221XL U101 ( .A0(n36), .A1(n550), .B0(n121), .B1(n543), .C0(n140), .Y(
        n135) );
  INVX1 U102 ( .A(n85), .Y(n36) );
  NOR2X1 U104 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U105 ( .A(n34), .B(n223), .Y(n183) );
  INVX1 U106 ( .A(n118), .Y(n70) );
  NAND2X1 U107 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U108 ( .A(n233), .Y(n55) );
  INVX1 U109 ( .A(n223), .Y(n59) );
  NOR2X1 U110 ( .A(n57), .B(n55), .Y(n197) );
  OAI221XL U111 ( .A0(n58), .A1(n545), .B0(n98), .B1(n94), .C0(n18), .Y(n347)
         );
  INVX1 U112 ( .A(n199), .Y(n18) );
  INVX1 U113 ( .A(n127), .Y(n35) );
  NOR2X1 U114 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U115 ( .A(n212), .Y(n41) );
  INVX1 U116 ( .A(n306), .Y(n58) );
  INVX1 U117 ( .A(n158), .Y(n42) );
  INVX1 U118 ( .A(n87), .Y(n38) );
  INVX1 U119 ( .A(n210), .Y(n44) );
  NAND2X1 U120 ( .A(n63), .B(n535), .Y(n243) );
  OAI22X1 U121 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U122 ( .A0(n61), .A1(n548), .B0(n556), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U123 ( .A0(n556), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U124 ( .A(n116), .B(n229), .Y(n244) );
  NOR2X1 U125 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U126 ( .A0(n94), .A1(n207), .B0(n545), .B1(n538), .Y(n242) );
  CLKINVX3 U127 ( .A(n113), .Y(n50) );
  CLKINVX3 U128 ( .A(n181), .Y(n63) );
  AOI22X1 U129 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U130 ( .A0(n98), .A1(n545), .B0(n30), .B1(n543), .C0(n99), .Y(n91)
         );
  OAI221XL U131 ( .A0(n42), .A1(n545), .B0(n51), .B1(n543), .C0(n95), .Y(n92)
         );
  INVX1 U132 ( .A(n104), .Y(n30) );
  NAND2X1 U133 ( .A(n556), .B(n96), .Y(n187) );
  NAND2X1 U134 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U135 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  OAI221XL U136 ( .A0(n536), .A1(n196), .B0(n197), .B1(n545), .C0(n198), .Y(
        n195) );
  AOI211X1 U137 ( .A0(n201), .A1(n556), .B0(n202), .C0(n203), .Y(n200) );
  AOI22X1 U138 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U139 ( .A0(n35), .A1(n545), .B0(n44), .B1(n543), .C0(n333), .Y(n332) );
  OAI211X1 U140 ( .A0(n326), .A1(n550), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U141 ( .A0(n35), .A1(n556), .B0(n39), .B1(n552), .Y(n333) );
  AOI22X1 U142 ( .A0(n548), .A1(n63), .B0(n247), .B1(n539), .Y(n334) );
  AOI21X1 U143 ( .A0(n115), .A1(n243), .B0(n550), .Y(n360) );
  INVX1 U144 ( .A(n120), .Y(n4) );
  AND2X2 U145 ( .A(n165), .B(n166), .Y(n129) );
  OAI21XL U146 ( .A0(n165), .A1(n550), .B0(n187), .Y(n266) );
  INVX1 U147 ( .A(n284), .Y(n10) );
  OAI31X1 U148 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U149 ( .A0(n541), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U150 ( .A(n147), .Y(n47) );
  OAI22X1 U152 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U153 ( .A0(n556), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U154 ( .A0(n11), .A1(n535), .B0(n27), .B1(n556), .C0(n307), .Y(n302) );
  OAI22X1 U155 ( .A0(n64), .A1(n543), .B0(n550), .B1(n306), .Y(n304) );
  AOI222X1 U156 ( .A0(n56), .A1(n540), .B0(n60), .B1(n554), .C0(n547), .C1(n71), .Y(n356) );
  AOI21X1 U157 ( .A0(n50), .A1(n556), .B0(n366), .Y(n365) );
  AOI2BB2X1 U158 ( .B0(n11), .B1(n535), .A0N(n536), .A1N(n247), .Y(n246) );
  CLKINVX8 U159 ( .A(n546), .Y(n545) );
  CLKINVX3 U160 ( .A(n541), .Y(n539) );
  NOR2X1 U161 ( .A(n545), .B(n535), .Y(n202) );
  AOI222X1 U162 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n540), 
        .Y(n198) );
  AOI221X1 U163 ( .A0(n321), .A1(n553), .B0(n540), .B1(n311), .C0(n327), .Y(
        n315) );
  OAI221XL U164 ( .A0(n536), .A1(n209), .B0(n545), .B1(n103), .C0(n288), .Y(
        n327) );
  AOI221X1 U165 ( .A0(n4), .A1(n71), .B0(n553), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI2BB1X1 U167 ( .A0N(n142), .A1N(n548), .B0(n187), .Y(n186) );
  NOR2X1 U168 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U169 ( .A0(n54), .A1(n545), .B0(n33), .B1(n543), .C0(n232), .Y(n217) );
  INVX1 U170 ( .A(n234), .Y(n54) );
  AOI32X1 U171 ( .A0(n34), .A1(n181), .A2(n556), .B0(n553), .B1(n233), .Y(n232) );
  INVX1 U172 ( .A(n115), .Y(n67) );
  AOI211X1 U173 ( .A0(n48), .A1(n556), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U174 ( .A(n114), .Y(n6) );
  AOI211X1 U175 ( .A0(n60), .A1(n540), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U176 ( .A(n545), .B(n39), .C(n61), .Y(n364) );
  INVX1 U177 ( .A(n259), .Y(n13) );
  OAI221XL U178 ( .A0(n536), .A1(n168), .B0(n164), .B1(n551), .C0(n169), .Y(
        n150) );
  AOI22X1 U179 ( .A0(n549), .A1(n34), .B0(n48), .B1(n539), .Y(n169) );
  AOI211X1 U180 ( .A0(n554), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  AOI211X1 U181 ( .A0(n45), .A1(n540), .B0(n204), .C0(n205), .Y(n192) );
  INVX1 U182 ( .A(n209), .Y(n45) );
  NAND2BX1 U183 ( .AN(n97), .B(n206), .Y(n205) );
  OAI222X1 U184 ( .A0(n551), .A1(n207), .B0(n181), .B1(n120), .C0(n545), .C1(
        n208), .Y(n204) );
  CLKINVX3 U185 ( .A(n555), .Y(n551) );
  INVX1 U186 ( .A(n125), .Y(n7) );
  AOI221X1 U187 ( .A0(n126), .A1(n552), .B0(n127), .B1(n549), .C0(n128), .Y(
        n125) );
  OAI21XL U188 ( .A0(n536), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U189 ( .A(n536), .Y(n16) );
  NOR2X1 U190 ( .A(n39), .B(n57), .Y(n179) );
  NAND3X1 U191 ( .A(n538), .B(n113), .C(n540), .Y(n89) );
  NAND2X1 U192 ( .A(n214), .B(n142), .Y(n90) );
  NAND2X1 U193 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U194 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U195 ( .A(n538), .B(n166), .Y(n311) );
  NOR2BX1 U196 ( .AN(n229), .B(n68), .Y(n164) );
  AOI21X1 U197 ( .A0(n181), .A1(n182), .B0(n536), .Y(n180) );
  AOI22X1 U198 ( .A0(n49), .A1(n548), .B0(n556), .B1(n141), .Y(n140) );
  AOI22X1 U199 ( .A0(n57), .A1(n546), .B0(n555), .B1(n113), .Y(n239) );
  AOI22X1 U200 ( .A0(n547), .A1(n311), .B0(n50), .B1(n539), .Y(n350) );
  NOR2X1 U201 ( .A(n138), .B(n536), .Y(n97) );
  NAND2X1 U202 ( .A(n243), .B(n142), .Y(n127) );
  INVX1 U203 ( .A(n154), .Y(n25) );
  NAND2X1 U204 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U205 ( .A(n138), .Y(n56) );
  NAND2X1 U206 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U207 ( .A(n64), .B(n124), .Y(n121) );
  AOI211X1 U208 ( .A0(n556), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  OAI2BB2X1 U209 ( .B0(n545), .B1(n183), .A0N(n188), .A1N(n540), .Y(n335) );
  AOI21X1 U210 ( .A0(n301), .A1(n337), .B0(n550), .Y(n336) );
  NAND2X1 U211 ( .A(n538), .B(n214), .Y(n126) );
  NAND2X1 U212 ( .A(n138), .B(n102), .Y(n227) );
  NAND2X1 U213 ( .A(n103), .B(n165), .Y(n188) );
  AOI21X1 U214 ( .A0(n556), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U215 ( .A0(n102), .A1(n103), .B0(n550), .Y(n101) );
  OAI221XL U216 ( .A0(n65), .A1(n551), .B0(n31), .B1(n536), .C0(n149), .Y(n143) );
  AOI2BB2X1 U217 ( .B0(n539), .B1(n87), .A0N(n545), .A1N(n121), .Y(n149) );
  INVX1 U218 ( .A(n337), .Y(n65) );
  INVX1 U219 ( .A(n208), .Y(n29) );
  INVX1 U220 ( .A(n299), .Y(n11) );
  INVX1 U221 ( .A(n100), .Y(n33) );
  AOI221XL U222 ( .A0(n556), .A1(n52), .B0(n548), .B1(n123), .C0(n324), .Y(
        n316) );
  INVX1 U223 ( .A(n326), .Y(n52) );
  OAI32X1 U224 ( .A0(n542), .A1(n63), .A2(n325), .B0(n37), .B1(n551), .Y(n324)
         );
  INVX1 U225 ( .A(n196), .Y(n31) );
  OAI221XL U226 ( .A0(n56), .A1(n545), .B0(n32), .B1(n542), .C0(n163), .Y(n151) );
  INVX1 U227 ( .A(n167), .Y(n32) );
  AOI22X1 U228 ( .A0(n164), .A1(n556), .B0(n129), .B1(n552), .Y(n163) );
  INVX1 U229 ( .A(n141), .Y(n27) );
  INVX1 U230 ( .A(n96), .Y(n40) );
  AOI31X1 U231 ( .A0(n102), .A1(n138), .A2(n556), .B0(n8), .Y(n137) );
  INVX1 U232 ( .A(n89), .Y(n8) );
  INVX1 U233 ( .A(n185), .Y(n19) );
  INVX1 U234 ( .A(n540), .Y(n542) );
  INVX1 U235 ( .A(n540), .Y(n543) );
  AOI211X1 U236 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U237 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI2BB2X1 U238 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  AOI211X1 U239 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U240 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U241 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  OAI21X2 U242 ( .A0(n534), .A1(n131), .B0(n132), .Y(d[6]) );
  OAI2BB1X1 U243 ( .A0N(n133), .A1N(n134), .B0(n534), .Y(n132) );
  AOI221X1 U244 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131) );
  AOI22X1 U245 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  OAI2BB1X1 U246 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI22X1 U247 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  AOI22X1 U248 ( .A0(n533), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U249 ( .A0(n61), .A1(n551), .B0(n545), .B1(n260), .C0(n261), .Y(
        n254) );
  OAI221XL U250 ( .A0(n41), .A1(n545), .B0(n543), .B1(n181), .C0(n256), .Y(
        n255) );
  AOI21X1 U251 ( .A0(n33), .A1(n16), .B0(n262), .Y(n261) );
  AOI22X1 U252 ( .A0(n348), .A1(n26), .B0(n533), .B1(n349), .Y(n342) );
  OAI221XL U253 ( .A0(n536), .A1(n166), .B0(n286), .B1(n545), .C0(n351), .Y(
        n348) );
  OAI211X1 U254 ( .A0(n88), .A1(n550), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U255 ( .B0(n539), .B1(n196), .A0N(n550), .A1N(n179), .Y(n351) );
  OAI22X1 U256 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U257 ( .A0(n549), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U258 ( .A0(n56), .A1(n4), .B0(n547), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U259 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U260 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U261 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U262 ( .A0(n61), .A1(n554), .B0(n547), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U263 ( .A0(n542), .A1(n71), .B0(n37), .B1(n550), .Y(n157) );
  OAI22X1 U264 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U265 ( .A0(n549), .A1(n111), .B0(n47), .B1(n540), .C0(n112), .Y(
        n109) );
  AOI221X1 U266 ( .A0(n556), .A1(n115), .B0(n553), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U267 ( .A0(n536), .A1(n113), .B0(n44), .B1(n551), .C0(n114), .Y(
        n112) );
  AOI211X1 U268 ( .A0(n55), .A1(n556), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U269 ( .A0(n114), .A1(n206), .A2(n273), .B0(n533), .Y(n272) );
  OAI22X1 U270 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U271 ( .B0(n70), .B1(n554), .A0N(n90), .A1N(n545), .Y(n273) );
  AOI2BB2X1 U272 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  OAI221XL U273 ( .A0(n46), .A1(n551), .B0(n545), .B1(n116), .C0(n267), .Y(
        n264) );
  AOI221XL U274 ( .A0(n548), .A1(n247), .B0(n212), .B1(n540), .C0(n266), .Y(
        n265) );
  AOI22X1 U275 ( .A0(n539), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  AOI22X1 U276 ( .A0(n554), .A1(n532), .B0(n539), .B1(n66), .Y(n292) );
  AOI22X1 U277 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U278 ( .A0(n63), .A1(n545), .B0(n542), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U279 ( .A0(n38), .A1(n536), .B0(n545), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U281 ( .A0(n179), .A1(n552), .B0(n180), .Y(n178) );
  AOI22X1 U282 ( .A0(n533), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U283 ( .A0(n43), .A1(n545), .B0(n541), .B1(n34), .C0(n365), .Y(n361) );
  OAI221XL U284 ( .A0(n532), .A1(n120), .B0(n201), .B1(n551), .C0(n363), .Y(
        n362) );
  INVX1 U285 ( .A(n260), .Y(n43) );
  AOI22X1 U286 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  OAI21XL U287 ( .A0(n321), .A1(n536), .B0(n322), .Y(n318) );
  OAI221XL U288 ( .A0(n551), .A1(n113), .B0(n88), .B1(n545), .C0(n320), .Y(
        n319) );
  AOI31X1 U289 ( .A0(n538), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  INVX1 U290 ( .A(n312), .Y(d[1]) );
  AOI22X1 U291 ( .A0(n534), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U292 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  OAI221XL U293 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  INVX1 U294 ( .A(n170), .Y(d[5]) );
  AOI22X1 U295 ( .A0(n171), .A1(n21), .B0(n534), .B1(n172), .Y(n170) );
  OAI221XL U296 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  OAI221XL U297 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  CLKINVX3 U298 ( .A(n532), .Y(n71) );
  OAI21XL U299 ( .A0(n545), .A1(n537), .B0(n120), .Y(n276) );
  NAND2X1 U300 ( .A(n63), .B(n531), .Y(n168) );
  AOI21X1 U301 ( .A0(n224), .A1(n243), .B0(n545), .Y(n295) );
  INVX1 U302 ( .A(n531), .Y(n74) );
  OAI21XL U303 ( .A0(n73), .A1(n301), .B0(n550), .Y(n323) );
  OAI21XL U304 ( .A0(n536), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U305 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U306 ( .A(n162), .Y(n5) );
  AOI211X1 U307 ( .A0(n39), .A1(n540), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U308 ( .A0(n551), .A1(n116), .B0(n73), .B1(n230), .C0(n545), .C1(
        n102), .Y(n275) );
  NAND2X1 U309 ( .A(n62), .B(n552), .Y(n287) );
  NOR2BX1 U310 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U311 ( .A(n82), .Y(n536) );
  NAND2X1 U312 ( .A(n73), .B(n20), .Y(n82) );
  OAI221XL U313 ( .A0(n531), .A1(n259), .B0(n94), .B1(n214), .C0(n287), .Y(
        n293) );
  BUFX3 U314 ( .A(n139), .Y(n538) );
  NAND2X1 U315 ( .A(n531), .B(n537), .Y(n139) );
  AOI211X1 U316 ( .A0(n540), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  OAI222X1 U317 ( .A0(n551), .A1(n167), .B0(n339), .B1(n536), .C0(n545), .C1(
        n34), .Y(n338) );
  AOI21X1 U318 ( .A0(n537), .A1(n535), .B0(n65), .Y(n339) );
  AOI211X1 U319 ( .A0(n533), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  OAI221XL U320 ( .A0(n545), .A1(n116), .B0(n321), .B1(n94), .C0(n359), .Y(
        n354) );
  AOI21X1 U321 ( .A0(n356), .A1(n357), .B0(n533), .Y(n355) );
  AOI31X1 U322 ( .A0(n556), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  INVX1 U323 ( .A(n93), .Y(n546) );
  INVX1 U324 ( .A(n83), .Y(n554) );
  INVX1 U325 ( .A(n83), .Y(n555) );
  INVX1 U326 ( .A(n544), .Y(n541) );
  INVX1 U327 ( .A(n94), .Y(n544) );
  AOI22X1 U328 ( .A0(n533), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U329 ( .A0(n545), .A1(n141), .B0(n551), .B1(n263), .C0(n29), .C1(
        n542), .Y(n277) );
  OAI221XL U330 ( .A0(n31), .A1(n536), .B0(n551), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U331 ( .B0(n88), .B1(n539), .A0N(n545), .A1N(n197), .Y(n279) );
  NAND2X1 U332 ( .A(n224), .B(n301), .Y(n148) );
  NOR2BX1 U333 ( .AN(n263), .B(n61), .Y(n321) );
  AOI21X1 U334 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI22X1 U335 ( .A0(n549), .A1(n85), .B0(n41), .B1(n539), .Y(n84) );
  AOI31X1 U336 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U337 ( .A0N(n223), .A1N(n224), .B0(n553), .Y(n220) );
  AOI22X1 U338 ( .A0(n29), .A1(n556), .B0(n222), .B1(n547), .Y(n221) );
  NAND2X1 U339 ( .A(n224), .B(n118), .Y(n208) );
  NAND2X1 U340 ( .A(n263), .B(n337), .Y(n167) );
  AOI21X1 U341 ( .A0(n263), .A1(n182), .B0(n545), .Y(n305) );
  AOI21X1 U342 ( .A0(n111), .A1(n538), .B0(n94), .Y(n203) );
  NAND2X1 U343 ( .A(n16), .B(n531), .Y(n206) );
  OAI21XL U344 ( .A0(n73), .A1(n243), .B0(n550), .Y(n245) );
  XNOR2X1 U345 ( .A(n20), .B(n531), .Y(n185) );
  NAND2X1 U346 ( .A(n539), .B(n537), .Y(n130) );
  XNOR2X1 U347 ( .A(n73), .B(n531), .Y(n161) );
  AOI21X1 U348 ( .A0(n90), .A1(n73), .B0(n556), .Y(n86) );
  AOI221X1 U349 ( .A0(n46), .A1(n540), .B0(n552), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U350 ( .A0(n536), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U351 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  AOI222X1 U352 ( .A0(n549), .A1(n210), .B0(n211), .B1(n212), .C0(n556), .C1(
        n537), .Y(n191) );
  OAI21XL U353 ( .A0(n73), .A1(n214), .B0(n550), .Y(n211) );
  NOR2X1 U354 ( .A(n62), .B(n55), .Y(n145) );
  AOI22X1 U355 ( .A0(n16), .A1(n66), .B0(n539), .B1(n147), .Y(n146) );
  INVX1 U356 ( .A(n148), .Y(n28) );
  AOI31X1 U357 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U358 ( .A0(n148), .A1(n73), .B0(n29), .B1(n553), .Y(n300) );
  INVX1 U359 ( .A(n93), .Y(n547) );
  INVX1 U360 ( .A(n93), .Y(n549) );
  INVX1 U361 ( .A(n93), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n358) );
  INVX1 U363 ( .A(n83), .Y(n552) );
  INVX1 U364 ( .A(n83), .Y(n553) );
  NOR2BX1 U365 ( .AN(n93), .B(n554), .Y(n309) );
  OAI22X2 U366 ( .A0(n340), .A1(n21), .B0(n534), .B1(n341), .Y(d[0]) );
  AOI22X1 U367 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U368 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI22X1 U369 ( .A0(n347), .A1(n26), .B0(n556), .B1(n90), .Y(n343) );
  AOI22X1 U370 ( .A0(n250), .A1(n21), .B0(n534), .B1(n251), .Y(n249) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  OAI22X1 U373 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U374 ( .A0(n548), .A1(n230), .B0(n556), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U375 ( .A0(n164), .A1(n547), .B0(a[2]), .B1(n227), .C0(n556), .C1(
        n228), .Y(n226) );
  OAI22X1 U376 ( .A0(n35), .A1(n543), .B0(n550), .B1(n537), .Y(n231) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI21XL U383 ( .A0(n66), .A1(n550), .B0(n259), .Y(n257) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI33X1 U385 ( .A0(n532), .A1(n540), .A2(n19), .B0(n185), .B1(n181), .B2(
        a[2]), .Y(n184) );
  AOI22X1 U386 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U387 ( .A(a[0]), .Y(n75) );
  AOI211X1 U388 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U389 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U390 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U391 ( .A(a[5]), .Y(n533) );
  OAI221XL U392 ( .A0(n536), .A1(n115), .B0(n121), .B1(n545), .C0(n122), .Y(
        n105) );
  AOI22X1 U393 ( .A0(n539), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_10 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556;

  OAI221X4 U4 ( .A0(n66), .A1(n536), .B0(n61), .B1(n551), .C0(n84), .Y(n81) );
  OAI221X4 U6 ( .A0(n86), .A1(n87), .B0(n88), .B1(n551), .C0(n89), .Y(n80) );
  OAI221X4 U28 ( .A0(n40), .A1(n551), .B0(n58), .B1(n545), .C0(n137), .Y(n136)
         );
  OAI221X4 U35 ( .A0(n145), .A1(n545), .B0(n28), .B1(n551), .C0(n146), .Y(n144) );
  OAI221X4 U70 ( .A0(n46), .A1(n551), .B0(n63), .B1(n545), .C0(n200), .Y(n194)
         );
  OAI221X4 U103 ( .A0(n551), .A1(n87), .B0(n94), .B1(n104), .C0(n246), .Y(n235) );
  OAI221X4 U151 ( .A0(n67), .A1(n551), .B0(n542), .B1(n538), .C0(n294), .Y(
        n282) );
  OAI221X4 U166 ( .A0(n308), .A1(n551), .B0(n545), .B1(n165), .C0(n162), .Y(
        n307) );
  OAI32X4 U280 ( .A0(n551), .A1(n56), .A2(n53), .B0(n542), .B1(n103), .Y(n366)
         );
  NAND2X4 U285 ( .A(n532), .B(n66), .Y(n181) );
  AOI221X1 U1 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n103) );
  NAND2X2 U5 ( .A(n531), .B(n532), .Y(n115) );
  NAND2X1 U7 ( .A(n56), .B(n531), .Y(n229) );
  NAND2X2 U8 ( .A(n66), .B(n71), .Y(n138) );
  NAND2X1 U9 ( .A(n531), .B(n181), .Y(n102) );
  NAND2X1 U10 ( .A(n533), .B(n75), .Y(n110) );
  NAND2X1 U11 ( .A(n531), .B(n539), .Y(n120) );
  NAND2X1 U12 ( .A(n39), .B(n531), .Y(n142) );
  NAND2X2 U13 ( .A(n537), .B(n181), .Y(n113) );
  NAND2X2 U14 ( .A(n66), .B(n535), .Y(n116) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n73) );
  CLKINVX3 U16 ( .A(n533), .Y(n26) );
  NAND2X2 U17 ( .A(a[0]), .B(n26), .Y(n156) );
  NAND2X2 U18 ( .A(n75), .B(n26), .Y(n154) );
  OAI22X2 U19 ( .A0(n534), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  OAI21X2 U20 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  AOI221X1 U21 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76) );
  OAI22X2 U22 ( .A0(n534), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  NAND2X1 U23 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U24 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI21XL U25 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  OAI222X4 U26 ( .A0(n541), .A1(n118), .B0(n119), .B1(n545), .C0(a[4]), .C1(
        n120), .Y(n117) );
  NAND2X1 U27 ( .A(n531), .B(a[4]), .Y(n224) );
  NAND2X1 U29 ( .A(a[4]), .B(n535), .Y(n263) );
  NAND2X2 U30 ( .A(n532), .B(a[4]), .Y(n111) );
  CLKINVX3 U31 ( .A(a[4]), .Y(n66) );
  NAND2X1 U32 ( .A(n53), .B(n16), .Y(n288) );
  CLKINVX3 U33 ( .A(n541), .Y(n540) );
  INVX1 U34 ( .A(n325), .Y(n34) );
  NAND2X1 U36 ( .A(n113), .B(n535), .Y(n214) );
  NAND2X1 U37 ( .A(n56), .B(n535), .Y(n233) );
  NAND2X1 U38 ( .A(n46), .B(n535), .Y(n209) );
  NAND2X1 U39 ( .A(n50), .B(n535), .Y(n301) );
  NAND2X1 U40 ( .A(n538), .B(n268), .Y(n212) );
  NAND2X1 U41 ( .A(n147), .B(n214), .Y(n207) );
  NAND2X1 U42 ( .A(n115), .B(n209), .Y(n210) );
  INVX1 U43 ( .A(n168), .Y(n62) );
  INVX1 U44 ( .A(n538), .Y(n53) );
  INVX1 U45 ( .A(n182), .Y(n57) );
  NOR2X1 U46 ( .A(n535), .B(n39), .Y(n325) );
  CLKINVX3 U47 ( .A(n555), .Y(n550) );
  NAND2X1 U48 ( .A(n535), .B(n71), .Y(n118) );
  NAND2X1 U49 ( .A(n138), .B(n535), .Y(n223) );
  NAND2X1 U50 ( .A(n39), .B(n535), .Y(n248) );
  NAND2X1 U51 ( .A(n181), .B(n535), .Y(n166) );
  NAND2X1 U52 ( .A(n229), .B(n248), .Y(n87) );
  CLKINVX3 U53 ( .A(n110), .Y(n23) );
  INVX1 U54 ( .A(n102), .Y(n61) );
  NAND2X1 U55 ( .A(n115), .B(n223), .Y(n306) );
  INVX1 U56 ( .A(n230), .Y(n69) );
  INVX1 U57 ( .A(n116), .Y(n64) );
  INVX1 U58 ( .A(n103), .Y(n68) );
  BUFX3 U59 ( .A(n74), .Y(n535) );
  NAND2X1 U60 ( .A(n50), .B(n531), .Y(n147) );
  NAND2X1 U61 ( .A(n111), .B(n535), .Y(n268) );
  NAND2X1 U62 ( .A(n531), .B(n113), .Y(n165) );
  NAND2X1 U63 ( .A(n531), .B(n138), .Y(n182) );
  INVX1 U64 ( .A(n537), .Y(n46) );
  NAND2X1 U65 ( .A(n16), .B(n532), .Y(n259) );
  NAND2X1 U66 ( .A(n111), .B(n147), .Y(n96) );
  NOR2X1 U67 ( .A(n537), .B(n535), .Y(n124) );
  CLKINVX3 U68 ( .A(n111), .Y(n39) );
  NAND2X1 U69 ( .A(n531), .B(n71), .Y(n230) );
  NAND2X1 U71 ( .A(n531), .B(n66), .Y(n337) );
  NAND2BX1 U72 ( .AN(n124), .B(n263), .Y(n196) );
  INVX1 U73 ( .A(n156), .Y(n24) );
  NAND2X1 U74 ( .A(n224), .B(n268), .Y(n141) );
  NAND2BX1 U75 ( .AN(n93), .B(n537), .Y(n299) );
  NAND2X1 U76 ( .A(n224), .B(n233), .Y(n104) );
  NAND2X1 U77 ( .A(n263), .B(n142), .Y(n100) );
  CLKINVX3 U78 ( .A(n534), .Y(n21) );
  CLKINVX3 U79 ( .A(n108), .Y(n22) );
  INVX1 U80 ( .A(n249), .Y(d[3]) );
  BUFX3 U81 ( .A(a[1]), .Y(n531) );
  NAND2X1 U82 ( .A(a[7]), .B(a[2]), .Y(n94) );
  NAND2X1 U83 ( .A(n533), .B(a[0]), .Y(n108) );
  INVX1 U84 ( .A(n238), .Y(n15) );
  NAND2X1 U85 ( .A(n59), .B(n540), .Y(n114) );
  NAND2X1 U86 ( .A(n51), .B(n556), .Y(n238) );
  INVX1 U87 ( .A(n288), .Y(n14) );
  NOR2X1 U88 ( .A(n550), .B(n325), .Y(n199) );
  NOR2X1 U89 ( .A(n49), .B(n62), .Y(n247) );
  NAND2X1 U90 ( .A(n222), .B(n540), .Y(n162) );
  INVX1 U91 ( .A(n301), .Y(n49) );
  INVX1 U92 ( .A(n248), .Y(n37) );
  INVX1 U93 ( .A(n166), .Y(n60) );
  INVX1 U94 ( .A(n207), .Y(n48) );
  INVX1 U95 ( .A(n228), .Y(n51) );
  INVX4 U96 ( .A(n536), .Y(n556) );
  NOR2BX1 U97 ( .AN(n214), .B(n69), .Y(n88) );
  NOR2X1 U98 ( .A(n53), .B(n70), .Y(n326) );
  AOI22X1 U99 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  OAI221XL U100 ( .A0(n36), .A1(n550), .B0(n121), .B1(n543), .C0(n140), .Y(
        n135) );
  INVX1 U101 ( .A(n85), .Y(n36) );
  NOR2X1 U102 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U104 ( .A(n34), .B(n223), .Y(n183) );
  INVX1 U105 ( .A(n118), .Y(n70) );
  NAND2X1 U106 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U107 ( .A(n233), .Y(n55) );
  INVX1 U108 ( .A(n223), .Y(n59) );
  NOR2X1 U109 ( .A(n57), .B(n55), .Y(n197) );
  OAI221XL U110 ( .A0(n58), .A1(n545), .B0(n98), .B1(n94), .C0(n18), .Y(n347)
         );
  INVX1 U111 ( .A(n199), .Y(n18) );
  INVX1 U112 ( .A(n127), .Y(n35) );
  NOR2X1 U113 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U114 ( .A(n212), .Y(n41) );
  INVX1 U115 ( .A(n306), .Y(n58) );
  INVX1 U116 ( .A(n158), .Y(n42) );
  INVX1 U117 ( .A(n87), .Y(n38) );
  INVX1 U118 ( .A(n210), .Y(n44) );
  NAND2X1 U119 ( .A(n63), .B(n535), .Y(n243) );
  OAI22X1 U120 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U121 ( .A0(n61), .A1(n548), .B0(n556), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U122 ( .A0(n556), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U123 ( .A(n116), .B(n229), .Y(n244) );
  NOR2X1 U124 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U125 ( .A0(n94), .A1(n207), .B0(n545), .B1(n538), .Y(n242) );
  CLKINVX3 U126 ( .A(n113), .Y(n50) );
  CLKINVX3 U127 ( .A(n181), .Y(n63) );
  AOI22X1 U128 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U129 ( .A0(n98), .A1(n545), .B0(n30), .B1(n543), .C0(n99), .Y(n91)
         );
  OAI221XL U130 ( .A0(n42), .A1(n545), .B0(n51), .B1(n543), .C0(n95), .Y(n92)
         );
  INVX1 U131 ( .A(n104), .Y(n30) );
  NAND2X1 U132 ( .A(n556), .B(n96), .Y(n187) );
  NAND2X1 U133 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U134 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  OAI221XL U135 ( .A0(n536), .A1(n196), .B0(n197), .B1(n545), .C0(n198), .Y(
        n195) );
  AOI211X1 U136 ( .A0(n201), .A1(n556), .B0(n202), .C0(n203), .Y(n200) );
  AOI22X1 U137 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U138 ( .A0(n35), .A1(n545), .B0(n44), .B1(n543), .C0(n333), .Y(n332) );
  OAI211X1 U139 ( .A0(n326), .A1(n550), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U140 ( .A0(n35), .A1(n556), .B0(n39), .B1(n552), .Y(n333) );
  AOI22X1 U141 ( .A0(n548), .A1(n63), .B0(n247), .B1(n539), .Y(n334) );
  AOI21X1 U142 ( .A0(n115), .A1(n243), .B0(n550), .Y(n360) );
  INVX1 U143 ( .A(n120), .Y(n4) );
  AND2X2 U144 ( .A(n165), .B(n166), .Y(n129) );
  OAI21XL U145 ( .A0(n165), .A1(n550), .B0(n187), .Y(n266) );
  INVX1 U146 ( .A(n284), .Y(n10) );
  OAI31X1 U147 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U148 ( .A0(n541), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U149 ( .A(n147), .Y(n47) );
  OAI22X1 U150 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U152 ( .A0(n556), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U153 ( .A0(n11), .A1(n535), .B0(n27), .B1(n556), .C0(n307), .Y(n302) );
  OAI22X1 U154 ( .A0(n64), .A1(n543), .B0(n550), .B1(n306), .Y(n304) );
  AOI222X1 U155 ( .A0(n56), .A1(n540), .B0(n60), .B1(n554), .C0(n547), .C1(n71), .Y(n356) );
  AOI21X1 U156 ( .A0(n50), .A1(n556), .B0(n366), .Y(n365) );
  AOI2BB2X1 U157 ( .B0(n11), .B1(n535), .A0N(n536), .A1N(n247), .Y(n246) );
  CLKINVX8 U158 ( .A(n546), .Y(n545) );
  CLKINVX3 U159 ( .A(n541), .Y(n539) );
  NOR2X1 U160 ( .A(n545), .B(n535), .Y(n202) );
  AOI222X1 U161 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n540), 
        .Y(n198) );
  AOI221X1 U162 ( .A0(n321), .A1(n553), .B0(n540), .B1(n311), .C0(n327), .Y(
        n315) );
  OAI221XL U163 ( .A0(n536), .A1(n209), .B0(n545), .B1(n103), .C0(n288), .Y(
        n327) );
  AOI221X1 U164 ( .A0(n4), .A1(n71), .B0(n553), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI2BB1X1 U165 ( .A0N(n142), .A1N(n548), .B0(n187), .Y(n186) );
  NOR2X1 U167 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U168 ( .A0(n54), .A1(n545), .B0(n33), .B1(n543), .C0(n232), .Y(n217) );
  INVX1 U169 ( .A(n234), .Y(n54) );
  AOI32X1 U170 ( .A0(n34), .A1(n181), .A2(n556), .B0(n553), .B1(n233), .Y(n232) );
  INVX1 U171 ( .A(n115), .Y(n67) );
  AOI211X1 U172 ( .A0(n48), .A1(n556), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U173 ( .A(n114), .Y(n6) );
  AOI211X1 U174 ( .A0(n60), .A1(n540), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U175 ( .A(n545), .B(n39), .C(n61), .Y(n364) );
  INVX1 U176 ( .A(n259), .Y(n13) );
  OAI221XL U177 ( .A0(n536), .A1(n168), .B0(n164), .B1(n551), .C0(n169), .Y(
        n150) );
  AOI22X1 U178 ( .A0(n549), .A1(n34), .B0(n48), .B1(n539), .Y(n169) );
  AOI211X1 U179 ( .A0(n554), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  AOI211X1 U180 ( .A0(n45), .A1(n540), .B0(n204), .C0(n205), .Y(n192) );
  INVX1 U181 ( .A(n209), .Y(n45) );
  NAND2BX1 U182 ( .AN(n97), .B(n206), .Y(n205) );
  OAI222X1 U183 ( .A0(n551), .A1(n207), .B0(n181), .B1(n120), .C0(n545), .C1(
        n208), .Y(n204) );
  CLKINVX3 U184 ( .A(n555), .Y(n551) );
  INVX1 U185 ( .A(n125), .Y(n7) );
  AOI221X1 U186 ( .A0(n126), .A1(n552), .B0(n127), .B1(n549), .C0(n128), .Y(
        n125) );
  OAI21XL U187 ( .A0(n536), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U188 ( .A(n536), .Y(n16) );
  NOR2X1 U189 ( .A(n39), .B(n57), .Y(n179) );
  NAND3X1 U190 ( .A(n538), .B(n113), .C(n540), .Y(n89) );
  NAND2X1 U191 ( .A(n214), .B(n142), .Y(n90) );
  NAND2X1 U192 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U193 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U194 ( .A(n538), .B(n166), .Y(n311) );
  NOR2BX1 U195 ( .AN(n229), .B(n68), .Y(n164) );
  AOI21X1 U196 ( .A0(n181), .A1(n182), .B0(n536), .Y(n180) );
  AOI22X1 U197 ( .A0(n49), .A1(n548), .B0(n556), .B1(n141), .Y(n140) );
  AOI22X1 U198 ( .A0(n57), .A1(n546), .B0(n555), .B1(n113), .Y(n239) );
  AOI22X1 U199 ( .A0(n547), .A1(n311), .B0(n50), .B1(n539), .Y(n350) );
  NOR2X1 U200 ( .A(n138), .B(n536), .Y(n97) );
  NAND2X1 U201 ( .A(n243), .B(n142), .Y(n127) );
  INVX1 U202 ( .A(n154), .Y(n25) );
  NAND2X1 U203 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U204 ( .A(n138), .Y(n56) );
  NAND2X1 U205 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U206 ( .A(n64), .B(n124), .Y(n121) );
  AOI211X1 U207 ( .A0(n556), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  OAI2BB2X1 U208 ( .B0(n545), .B1(n183), .A0N(n188), .A1N(n540), .Y(n335) );
  AOI21X1 U209 ( .A0(n301), .A1(n337), .B0(n550), .Y(n336) );
  NAND2X1 U210 ( .A(n538), .B(n214), .Y(n126) );
  NAND2X1 U211 ( .A(n138), .B(n102), .Y(n227) );
  NAND2X1 U212 ( .A(n103), .B(n165), .Y(n188) );
  AOI21X1 U213 ( .A0(n556), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U214 ( .A0(n102), .A1(n103), .B0(n550), .Y(n101) );
  OAI221XL U215 ( .A0(n65), .A1(n551), .B0(n31), .B1(n536), .C0(n149), .Y(n143) );
  AOI2BB2X1 U216 ( .B0(n539), .B1(n87), .A0N(n545), .A1N(n121), .Y(n149) );
  INVX1 U217 ( .A(n337), .Y(n65) );
  INVX1 U218 ( .A(n208), .Y(n29) );
  INVX1 U219 ( .A(n299), .Y(n11) );
  INVX1 U220 ( .A(n100), .Y(n33) );
  AOI221XL U221 ( .A0(n556), .A1(n52), .B0(n548), .B1(n123), .C0(n324), .Y(
        n316) );
  INVX1 U222 ( .A(n326), .Y(n52) );
  OAI32X1 U223 ( .A0(n542), .A1(n63), .A2(n325), .B0(n37), .B1(n551), .Y(n324)
         );
  INVX1 U224 ( .A(n196), .Y(n31) );
  OAI221XL U225 ( .A0(n56), .A1(n545), .B0(n32), .B1(n542), .C0(n163), .Y(n151) );
  INVX1 U226 ( .A(n167), .Y(n32) );
  AOI22X1 U227 ( .A0(n164), .A1(n556), .B0(n129), .B1(n552), .Y(n163) );
  INVX1 U228 ( .A(n141), .Y(n27) );
  INVX1 U229 ( .A(n96), .Y(n40) );
  AOI31X1 U230 ( .A0(n102), .A1(n138), .A2(n556), .B0(n8), .Y(n137) );
  INVX1 U231 ( .A(n89), .Y(n8) );
  INVX1 U232 ( .A(n185), .Y(n19) );
  INVX1 U233 ( .A(n540), .Y(n542) );
  INVX1 U234 ( .A(n540), .Y(n543) );
  AOI211X1 U235 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U236 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI2BB2X1 U237 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  AOI211X1 U238 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U239 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U240 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  OAI21X2 U241 ( .A0(n534), .A1(n131), .B0(n132), .Y(d[6]) );
  OAI2BB1X1 U242 ( .A0N(n133), .A1N(n134), .B0(n534), .Y(n132) );
  AOI221X1 U243 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131) );
  AOI22X1 U244 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  OAI2BB1X1 U245 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI22X1 U246 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  AOI22X1 U247 ( .A0(n533), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U248 ( .A0(n61), .A1(n551), .B0(n545), .B1(n260), .C0(n261), .Y(
        n254) );
  OAI221XL U249 ( .A0(n41), .A1(n545), .B0(n543), .B1(n181), .C0(n256), .Y(
        n255) );
  AOI21X1 U250 ( .A0(n33), .A1(n16), .B0(n262), .Y(n261) );
  AOI22X1 U251 ( .A0(n348), .A1(n26), .B0(n533), .B1(n349), .Y(n342) );
  OAI221XL U252 ( .A0(n536), .A1(n166), .B0(n286), .B1(n545), .C0(n351), .Y(
        n348) );
  OAI211X1 U253 ( .A0(n88), .A1(n550), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U254 ( .B0(n539), .B1(n196), .A0N(n550), .A1N(n179), .Y(n351) );
  OAI22X1 U255 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U256 ( .A0(n549), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U257 ( .A0(n56), .A1(n4), .B0(n547), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U258 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U259 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U260 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U261 ( .A0(n61), .A1(n554), .B0(n547), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U262 ( .A0(n542), .A1(n71), .B0(n37), .B1(n550), .Y(n157) );
  OAI22X1 U263 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U264 ( .A0(n549), .A1(n111), .B0(n47), .B1(n540), .C0(n112), .Y(
        n109) );
  AOI221X1 U265 ( .A0(n556), .A1(n115), .B0(n553), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U266 ( .A0(n536), .A1(n113), .B0(n44), .B1(n551), .C0(n114), .Y(
        n112) );
  AOI211X1 U267 ( .A0(n55), .A1(n556), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U268 ( .A0(n114), .A1(n206), .A2(n273), .B0(n533), .Y(n272) );
  OAI22X1 U269 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U270 ( .B0(n70), .B1(n554), .A0N(n90), .A1N(n545), .Y(n273) );
  AOI2BB2X1 U271 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  OAI221XL U272 ( .A0(n46), .A1(n551), .B0(n545), .B1(n116), .C0(n267), .Y(
        n264) );
  AOI221XL U273 ( .A0(n548), .A1(n247), .B0(n212), .B1(n540), .C0(n266), .Y(
        n265) );
  AOI22X1 U274 ( .A0(n539), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  AOI22X1 U275 ( .A0(n554), .A1(n532), .B0(n539), .B1(n66), .Y(n292) );
  AOI22X1 U276 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U277 ( .A0(n63), .A1(n545), .B0(n542), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U278 ( .A0(n38), .A1(n536), .B0(n545), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U279 ( .A0(n179), .A1(n552), .B0(n180), .Y(n178) );
  AOI22X1 U281 ( .A0(n533), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U282 ( .A0(n43), .A1(n545), .B0(n541), .B1(n34), .C0(n365), .Y(n361) );
  OAI221XL U283 ( .A0(n532), .A1(n120), .B0(n201), .B1(n551), .C0(n363), .Y(
        n362) );
  INVX1 U284 ( .A(n260), .Y(n43) );
  AOI22X1 U286 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  OAI21XL U287 ( .A0(n321), .A1(n536), .B0(n322), .Y(n318) );
  OAI221XL U288 ( .A0(n551), .A1(n113), .B0(n88), .B1(n545), .C0(n320), .Y(
        n319) );
  AOI31X1 U289 ( .A0(n538), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  INVX1 U290 ( .A(n312), .Y(d[1]) );
  AOI22X1 U291 ( .A0(n534), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U292 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  OAI221XL U293 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  INVX1 U294 ( .A(n170), .Y(d[5]) );
  AOI22X1 U295 ( .A0(n171), .A1(n21), .B0(n534), .B1(n172), .Y(n170) );
  OAI221XL U296 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  OAI221XL U297 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  CLKINVX3 U298 ( .A(n532), .Y(n71) );
  OAI21XL U299 ( .A0(n545), .A1(n537), .B0(n120), .Y(n276) );
  NAND2X1 U300 ( .A(n63), .B(n531), .Y(n168) );
  AOI21X1 U301 ( .A0(n224), .A1(n243), .B0(n545), .Y(n295) );
  INVX1 U302 ( .A(n531), .Y(n74) );
  OAI21XL U303 ( .A0(n73), .A1(n301), .B0(n550), .Y(n323) );
  OAI21XL U304 ( .A0(n536), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U305 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U306 ( .A(n162), .Y(n5) );
  AOI211X1 U307 ( .A0(n39), .A1(n540), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U308 ( .A0(n551), .A1(n116), .B0(n73), .B1(n230), .C0(n545), .C1(
        n102), .Y(n275) );
  NAND2X1 U309 ( .A(n62), .B(n552), .Y(n287) );
  NOR2BX1 U310 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U311 ( .A(n82), .Y(n536) );
  NAND2X1 U312 ( .A(n73), .B(n20), .Y(n82) );
  OAI221XL U313 ( .A0(n531), .A1(n259), .B0(n94), .B1(n214), .C0(n287), .Y(
        n293) );
  BUFX3 U314 ( .A(n139), .Y(n538) );
  NAND2X1 U315 ( .A(n531), .B(n537), .Y(n139) );
  AOI211X1 U316 ( .A0(n540), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  OAI222X1 U317 ( .A0(n551), .A1(n167), .B0(n339), .B1(n536), .C0(n545), .C1(
        n34), .Y(n338) );
  AOI21X1 U318 ( .A0(n537), .A1(n535), .B0(n65), .Y(n339) );
  AOI211X1 U319 ( .A0(n533), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  OAI221XL U320 ( .A0(n545), .A1(n116), .B0(n321), .B1(n94), .C0(n359), .Y(
        n354) );
  AOI21X1 U321 ( .A0(n356), .A1(n357), .B0(n533), .Y(n355) );
  AOI31X1 U322 ( .A0(n556), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  INVX1 U323 ( .A(n93), .Y(n546) );
  INVX1 U324 ( .A(n83), .Y(n554) );
  INVX1 U325 ( .A(n83), .Y(n555) );
  INVX1 U326 ( .A(n544), .Y(n541) );
  INVX1 U327 ( .A(n94), .Y(n544) );
  AOI22X1 U328 ( .A0(n533), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U329 ( .A0(n545), .A1(n141), .B0(n551), .B1(n263), .C0(n29), .C1(
        n542), .Y(n277) );
  OAI221XL U330 ( .A0(n31), .A1(n536), .B0(n551), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U331 ( .B0(n88), .B1(n539), .A0N(n545), .A1N(n197), .Y(n279) );
  NAND2X1 U332 ( .A(n224), .B(n301), .Y(n148) );
  NOR2BX1 U333 ( .AN(n263), .B(n61), .Y(n321) );
  AOI21X1 U334 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI22X1 U335 ( .A0(n549), .A1(n85), .B0(n41), .B1(n539), .Y(n84) );
  AOI31X1 U336 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U337 ( .A0N(n223), .A1N(n224), .B0(n553), .Y(n220) );
  AOI22X1 U338 ( .A0(n29), .A1(n556), .B0(n222), .B1(n547), .Y(n221) );
  NAND2X1 U339 ( .A(n224), .B(n118), .Y(n208) );
  NAND2X1 U340 ( .A(n263), .B(n337), .Y(n167) );
  AOI21X1 U341 ( .A0(n263), .A1(n182), .B0(n545), .Y(n305) );
  AOI21X1 U342 ( .A0(n111), .A1(n538), .B0(n94), .Y(n203) );
  NAND2X1 U343 ( .A(n16), .B(n531), .Y(n206) );
  OAI21XL U344 ( .A0(n73), .A1(n243), .B0(n550), .Y(n245) );
  XNOR2X1 U345 ( .A(n20), .B(n531), .Y(n185) );
  NAND2X1 U346 ( .A(n539), .B(n537), .Y(n130) );
  XNOR2X1 U347 ( .A(n73), .B(n531), .Y(n161) );
  AOI21X1 U348 ( .A0(n90), .A1(n73), .B0(n556), .Y(n86) );
  AOI221X1 U349 ( .A0(n46), .A1(n540), .B0(n552), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U350 ( .A0(n536), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U351 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  AOI222X1 U352 ( .A0(n549), .A1(n210), .B0(n211), .B1(n212), .C0(n556), .C1(
        n537), .Y(n191) );
  OAI21XL U353 ( .A0(n73), .A1(n214), .B0(n550), .Y(n211) );
  NOR2X1 U354 ( .A(n62), .B(n55), .Y(n145) );
  AOI22X1 U355 ( .A0(n16), .A1(n66), .B0(n539), .B1(n147), .Y(n146) );
  INVX1 U356 ( .A(n148), .Y(n28) );
  AOI31X1 U357 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U358 ( .A0(n148), .A1(n73), .B0(n29), .B1(n553), .Y(n300) );
  INVX1 U359 ( .A(n93), .Y(n547) );
  INVX1 U360 ( .A(n93), .Y(n549) );
  INVX1 U361 ( .A(n93), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n358) );
  INVX1 U363 ( .A(n83), .Y(n552) );
  INVX1 U364 ( .A(n83), .Y(n553) );
  NOR2BX1 U365 ( .AN(n93), .B(n554), .Y(n309) );
  OAI22X2 U366 ( .A0(n340), .A1(n21), .B0(n534), .B1(n341), .Y(d[0]) );
  AOI22X1 U367 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U368 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI22X1 U369 ( .A0(n347), .A1(n26), .B0(n556), .B1(n90), .Y(n343) );
  AOI22X1 U370 ( .A0(n250), .A1(n21), .B0(n534), .B1(n251), .Y(n249) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  OAI22X1 U373 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U374 ( .A0(n548), .A1(n230), .B0(n556), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U375 ( .A0(n164), .A1(n547), .B0(a[2]), .B1(n227), .C0(n556), .C1(
        n228), .Y(n226) );
  OAI22X1 U376 ( .A0(n35), .A1(n543), .B0(n550), .B1(n537), .Y(n231) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI21XL U383 ( .A0(n66), .A1(n550), .B0(n259), .Y(n257) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI33X1 U385 ( .A0(n532), .A1(n540), .A2(n19), .B0(n185), .B1(n181), .B2(
        a[2]), .Y(n184) );
  AOI22X1 U386 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U387 ( .A(a[0]), .Y(n75) );
  AOI211X1 U388 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U389 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U390 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U391 ( .A(a[5]), .Y(n533) );
  OAI221XL U392 ( .A0(n536), .A1(n115), .B0(n121), .B1(n545), .C0(n122), .Y(
        n105) );
  AOI22X1 U393 ( .A0(n539), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_8 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556;

  OAI221X4 U4 ( .A0(n66), .A1(n536), .B0(n61), .B1(n551), .C0(n84), .Y(n81) );
  OAI221X4 U6 ( .A0(n86), .A1(n87), .B0(n88), .B1(n551), .C0(n89), .Y(n80) );
  OAI222X4 U75 ( .A0(n551), .A1(n207), .B0(n181), .B1(n120), .C0(n545), .C1(
        n208), .Y(n204) );
  OAI32X4 U280 ( .A0(n551), .A1(n56), .A2(n53), .B0(n94), .B1(n103), .Y(n366)
         );
  AOI221X1 U1 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n103) );
  OAI222X1 U5 ( .A0(n94), .A1(n118), .B0(n119), .B1(n545), .C0(a[4]), .C1(n120), .Y(n117) );
  NAND2X2 U7 ( .A(n531), .B(n532), .Y(n115) );
  NAND2X1 U8 ( .A(n56), .B(n531), .Y(n229) );
  NAND2X2 U9 ( .A(n532), .B(n66), .Y(n181) );
  NAND2X1 U10 ( .A(n39), .B(n531), .Y(n142) );
  NAND2X2 U11 ( .A(n537), .B(n181), .Y(n113) );
  NAND2X2 U12 ( .A(n66), .B(n535), .Y(n116) );
  CLKINVX3 U13 ( .A(n533), .Y(n26) );
  NAND2X2 U14 ( .A(n66), .B(n71), .Y(n138) );
  NAND2X1 U15 ( .A(n531), .B(n181), .Y(n102) );
  CLKINVX3 U16 ( .A(a[2]), .Y(n73) );
  NAND2X1 U17 ( .A(n533), .B(n75), .Y(n110) );
  NAND2X2 U18 ( .A(n75), .B(n26), .Y(n154) );
  NAND2X2 U19 ( .A(a[0]), .B(n26), .Y(n156) );
  CLKINVX3 U20 ( .A(n534), .Y(n21) );
  OAI22X2 U21 ( .A0(n340), .A1(n21), .B0(n534), .B1(n341), .Y(d[0]) );
  OAI22X2 U22 ( .A0(n534), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  OAI21X2 U23 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  AOI221X1 U24 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76) );
  OAI22X2 U25 ( .A0(n534), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  OAI21X2 U26 ( .A0(n534), .A1(n131), .B0(n132), .Y(d[6]) );
  AOI221X1 U27 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131)
         );
  NAND2X1 U28 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U29 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI21XL U30 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  NAND2X1 U31 ( .A(a[4]), .B(n535), .Y(n263) );
  NAND2X1 U32 ( .A(n531), .B(a[4]), .Y(n224) );
  NAND2X2 U33 ( .A(n532), .B(a[4]), .Y(n111) );
  CLKINVX3 U34 ( .A(a[4]), .Y(n66) );
  CLKINVX3 U35 ( .A(n542), .Y(n540) );
  NAND2X1 U36 ( .A(n53), .B(n16), .Y(n288) );
  INVX1 U37 ( .A(n325), .Y(n34) );
  NAND2X1 U38 ( .A(n113), .B(n535), .Y(n214) );
  CLKINVX3 U39 ( .A(n555), .Y(n550) );
  NAND2X1 U40 ( .A(n56), .B(n535), .Y(n233) );
  NAND2X1 U41 ( .A(n50), .B(n535), .Y(n301) );
  NAND2X1 U42 ( .A(n538), .B(n268), .Y(n212) );
  NAND2X1 U43 ( .A(n115), .B(n209), .Y(n210) );
  NAND2X1 U44 ( .A(n147), .B(n214), .Y(n207) );
  INVX1 U45 ( .A(n168), .Y(n62) );
  INVX1 U46 ( .A(n538), .Y(n53) );
  INVX1 U47 ( .A(n182), .Y(n57) );
  NOR2X1 U48 ( .A(n535), .B(n39), .Y(n325) );
  NAND2X1 U49 ( .A(n535), .B(n71), .Y(n118) );
  NAND2X1 U50 ( .A(n138), .B(n535), .Y(n223) );
  NAND2X1 U51 ( .A(n39), .B(n535), .Y(n248) );
  NAND2X1 U52 ( .A(n181), .B(n535), .Y(n166) );
  NAND2X1 U53 ( .A(n229), .B(n248), .Y(n87) );
  INVX1 U54 ( .A(n102), .Y(n61) );
  NAND2X1 U55 ( .A(n115), .B(n223), .Y(n306) );
  INVX1 U56 ( .A(n230), .Y(n69) );
  INVX1 U57 ( .A(n116), .Y(n64) );
  INVX1 U58 ( .A(n103), .Y(n68) );
  BUFX3 U59 ( .A(n74), .Y(n535) );
  NAND2X1 U60 ( .A(n50), .B(n531), .Y(n147) );
  NAND2X1 U61 ( .A(n531), .B(n539), .Y(n120) );
  NAND2X1 U62 ( .A(n111), .B(n535), .Y(n268) );
  NAND2X1 U63 ( .A(n531), .B(n113), .Y(n165) );
  NAND2X1 U64 ( .A(n531), .B(n138), .Y(n182) );
  INVX1 U65 ( .A(n312), .Y(d[1]) );
  INVX1 U66 ( .A(n170), .Y(d[5]) );
  NAND2X1 U67 ( .A(n16), .B(n532), .Y(n259) );
  INVX1 U68 ( .A(n537), .Y(n46) );
  NAND2X1 U69 ( .A(n111), .B(n147), .Y(n96) );
  NOR2X1 U70 ( .A(n537), .B(n535), .Y(n124) );
  CLKINVX3 U71 ( .A(n111), .Y(n39) );
  NAND2X1 U72 ( .A(n531), .B(n71), .Y(n230) );
  NAND2X1 U73 ( .A(n531), .B(n66), .Y(n337) );
  NAND2BX1 U74 ( .AN(n124), .B(n263), .Y(n196) );
  INVX1 U76 ( .A(n156), .Y(n24) );
  NAND2X1 U77 ( .A(n224), .B(n268), .Y(n141) );
  NAND2BX1 U78 ( .AN(n93), .B(n537), .Y(n299) );
  NAND2X1 U79 ( .A(n224), .B(n233), .Y(n104) );
  NAND2X1 U80 ( .A(n263), .B(n142), .Y(n100) );
  CLKINVX3 U81 ( .A(n108), .Y(n22) );
  BUFX3 U82 ( .A(a[1]), .Y(n531) );
  NAND2X1 U83 ( .A(a[7]), .B(a[2]), .Y(n94) );
  INVX1 U84 ( .A(n249), .Y(d[3]) );
  NAND2X1 U85 ( .A(n533), .B(a[0]), .Y(n108) );
  INVX1 U86 ( .A(n238), .Y(n15) );
  NAND2X1 U87 ( .A(n59), .B(n540), .Y(n114) );
  NAND2X1 U88 ( .A(n51), .B(n556), .Y(n238) );
  INVX1 U89 ( .A(n288), .Y(n14) );
  NOR2X1 U90 ( .A(n550), .B(n325), .Y(n199) );
  NOR2X1 U91 ( .A(n49), .B(n62), .Y(n247) );
  NAND2X1 U92 ( .A(n222), .B(n540), .Y(n162) );
  INVX1 U93 ( .A(n301), .Y(n49) );
  INVX1 U94 ( .A(n248), .Y(n37) );
  INVX1 U95 ( .A(n166), .Y(n60) );
  INVX1 U96 ( .A(n207), .Y(n48) );
  INVX1 U97 ( .A(n228), .Y(n51) );
  INVX1 U98 ( .A(n210), .Y(n44) );
  INVX4 U99 ( .A(n536), .Y(n556) );
  NOR2BX1 U100 ( .AN(n214), .B(n69), .Y(n88) );
  NOR2X1 U101 ( .A(n53), .B(n70), .Y(n326) );
  NOR2X1 U102 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U103 ( .A(n34), .B(n223), .Y(n183) );
  INVX1 U104 ( .A(n118), .Y(n70) );
  NAND2X1 U105 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U106 ( .A(n233), .Y(n55) );
  INVX1 U107 ( .A(n223), .Y(n59) );
  NOR2X1 U108 ( .A(n57), .B(n55), .Y(n197) );
  OAI221XL U109 ( .A0(n58), .A1(n545), .B0(n98), .B1(n543), .C0(n18), .Y(n347)
         );
  INVX1 U110 ( .A(n199), .Y(n18) );
  INVX1 U111 ( .A(n127), .Y(n35) );
  NOR2X1 U112 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U113 ( .A(n212), .Y(n41) );
  NOR2X1 U114 ( .A(n62), .B(n55), .Y(n145) );
  INVX1 U115 ( .A(n306), .Y(n58) );
  INVX1 U116 ( .A(n158), .Y(n42) );
  INVX1 U117 ( .A(n87), .Y(n38) );
  NAND2X1 U118 ( .A(n63), .B(n535), .Y(n243) );
  NAND2X1 U119 ( .A(n46), .B(n535), .Y(n209) );
  OAI22X1 U120 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U121 ( .A0(n61), .A1(n548), .B0(n556), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U122 ( .A0(n556), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U123 ( .A(n116), .B(n229), .Y(n244) );
  NOR2X1 U124 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U125 ( .A0(n542), .A1(n207), .B0(n545), .B1(n538), .Y(n242) );
  CLKINVX3 U126 ( .A(n113), .Y(n50) );
  NAND2X1 U127 ( .A(n214), .B(n142), .Y(n90) );
  CLKINVX3 U128 ( .A(n181), .Y(n63) );
  AOI22X1 U129 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U130 ( .A0(n98), .A1(n545), .B0(n30), .B1(n541), .C0(n99), .Y(n91)
         );
  OAI221XL U131 ( .A0(n42), .A1(n545), .B0(n51), .B1(n542), .C0(n95), .Y(n92)
         );
  INVX1 U132 ( .A(n104), .Y(n30) );
  NAND2X1 U133 ( .A(n556), .B(n96), .Y(n187) );
  NAND2X1 U134 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U135 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  OAI221XL U136 ( .A0(n46), .A1(n551), .B0(n63), .B1(n545), .C0(n200), .Y(n194) );
  OAI221XL U137 ( .A0(n536), .A1(n196), .B0(n197), .B1(n545), .C0(n198), .Y(
        n195) );
  AOI211X1 U138 ( .A0(n201), .A1(n556), .B0(n202), .C0(n203), .Y(n200) );
  AOI22X1 U139 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U140 ( .A0(n35), .A1(n545), .B0(n44), .B1(n542), .C0(n333), .Y(n332) );
  OAI211X1 U141 ( .A0(n326), .A1(n550), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U142 ( .A0(n35), .A1(n16), .B0(n39), .B1(n553), .Y(n333) );
  AOI22X1 U143 ( .A0(n548), .A1(n63), .B0(n247), .B1(n539), .Y(n334) );
  AOI21X1 U144 ( .A0(n115), .A1(n243), .B0(n550), .Y(n360) );
  INVX1 U145 ( .A(n120), .Y(n4) );
  AND2X2 U146 ( .A(n165), .B(n166), .Y(n129) );
  NAND2X1 U147 ( .A(n538), .B(n214), .Y(n126) );
  OAI21XL U148 ( .A0(n165), .A1(n550), .B0(n187), .Y(n266) );
  INVX1 U149 ( .A(n284), .Y(n10) );
  OAI31X1 U150 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U151 ( .A0(n541), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U152 ( .A(n147), .Y(n47) );
  OAI22X1 U153 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U154 ( .A0(n556), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U155 ( .A0(n11), .A1(n535), .B0(n27), .B1(n556), .C0(n307), .Y(n302) );
  OAI22X1 U156 ( .A0(n64), .A1(n542), .B0(n550), .B1(n306), .Y(n304) );
  AOI222X1 U157 ( .A0(n56), .A1(n540), .B0(n60), .B1(n552), .C0(n547), .C1(n71), .Y(n356) );
  AOI21X1 U158 ( .A0(n50), .A1(n556), .B0(n366), .Y(n365) );
  OAI221XL U159 ( .A0(n551), .A1(n87), .B0(n543), .B1(n104), .C0(n246), .Y(
        n235) );
  AOI2BB2X1 U160 ( .B0(n11), .B1(n535), .A0N(n536), .A1N(n247), .Y(n246) );
  CLKINVX8 U161 ( .A(n546), .Y(n545) );
  CLKINVX3 U162 ( .A(n541), .Y(n539) );
  NOR2X1 U163 ( .A(n545), .B(n535), .Y(n202) );
  AOI211X1 U164 ( .A0(n45), .A1(n540), .B0(n204), .C0(n205), .Y(n192) );
  INVX1 U165 ( .A(n209), .Y(n45) );
  NAND2BX1 U166 ( .AN(n97), .B(n206), .Y(n205) );
  AOI222X1 U167 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n540), 
        .Y(n198) );
  AOI221X1 U168 ( .A0(n321), .A1(n554), .B0(n540), .B1(n311), .C0(n327), .Y(
        n315) );
  OAI221XL U169 ( .A0(n536), .A1(n209), .B0(n545), .B1(n103), .C0(n288), .Y(
        n327) );
  AOI221X1 U170 ( .A0(n4), .A1(n71), .B0(n554), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI2BB1X1 U171 ( .A0N(n142), .A1N(n547), .B0(n187), .Y(n186) );
  OAI221XL U172 ( .A0(n308), .A1(n551), .B0(n545), .B1(n165), .C0(n162), .Y(
        n307) );
  NOR2X1 U173 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U174 ( .A0(n54), .A1(n545), .B0(n33), .B1(n94), .C0(n232), .Y(n217)
         );
  INVX1 U175 ( .A(n234), .Y(n54) );
  AOI32X1 U176 ( .A0(n34), .A1(n181), .A2(n556), .B0(n554), .B1(n233), .Y(n232) );
  OAI221XL U177 ( .A0(n67), .A1(n551), .B0(n541), .B1(n538), .C0(n294), .Y(
        n282) );
  INVX1 U178 ( .A(n115), .Y(n67) );
  AOI211X1 U179 ( .A0(n48), .A1(n556), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U180 ( .A(n114), .Y(n6) );
  AOI211X1 U181 ( .A0(n60), .A1(n540), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U182 ( .A(n545), .B(n39), .C(n61), .Y(n364) );
  INVX1 U183 ( .A(n259), .Y(n13) );
  OAI221XL U184 ( .A0(n536), .A1(n168), .B0(n164), .B1(n551), .C0(n169), .Y(
        n150) );
  AOI22X1 U185 ( .A0(n549), .A1(n34), .B0(n48), .B1(n539), .Y(n169) );
  AOI211X1 U186 ( .A0(n554), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  CLKINVX3 U187 ( .A(n555), .Y(n551) );
  INVX1 U188 ( .A(n544), .Y(n542) );
  INVX1 U189 ( .A(n125), .Y(n7) );
  AOI221X1 U190 ( .A0(n126), .A1(n553), .B0(n127), .B1(n549), .C0(n128), .Y(
        n125) );
  OAI21XL U191 ( .A0(n536), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U192 ( .A(n536), .Y(n16) );
  NOR2X1 U193 ( .A(n39), .B(n57), .Y(n179) );
  CLKINVX3 U194 ( .A(n110), .Y(n23) );
  NAND3X1 U195 ( .A(n538), .B(n113), .C(n540), .Y(n89) );
  NAND2X1 U196 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U197 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U198 ( .A(n538), .B(n166), .Y(n311) );
  NOR2BX1 U199 ( .AN(n229), .B(n68), .Y(n164) );
  AOI21X1 U200 ( .A0(n181), .A1(n182), .B0(n536), .Y(n180) );
  OAI221XL U201 ( .A0(n36), .A1(n550), .B0(n121), .B1(n541), .C0(n140), .Y(
        n135) );
  INVX1 U202 ( .A(n85), .Y(n36) );
  AOI22X1 U203 ( .A0(n49), .A1(n548), .B0(n556), .B1(n141), .Y(n140) );
  AOI22X1 U204 ( .A0(n57), .A1(n546), .B0(n552), .B1(n113), .Y(n239) );
  AOI22X1 U205 ( .A0(n547), .A1(n311), .B0(n50), .B1(n539), .Y(n350) );
  NOR2X1 U206 ( .A(n138), .B(n536), .Y(n97) );
  NAND2X1 U207 ( .A(n243), .B(n142), .Y(n127) );
  INVX1 U208 ( .A(n154), .Y(n25) );
  NAND2X1 U209 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U210 ( .A(n138), .Y(n56) );
  NAND2X1 U211 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U212 ( .A(n64), .B(n124), .Y(n121) );
  AOI211X1 U213 ( .A0(n556), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  OAI2BB2X1 U214 ( .B0(n545), .B1(n183), .A0N(n188), .A1N(n540), .Y(n335) );
  AOI21X1 U215 ( .A0(n301), .A1(n337), .B0(n550), .Y(n336) );
  NAND2X1 U216 ( .A(n138), .B(n102), .Y(n227) );
  NAND2X1 U217 ( .A(n103), .B(n165), .Y(n188) );
  AOI21X1 U218 ( .A0(n556), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U219 ( .A0(n102), .A1(n103), .B0(n550), .Y(n101) );
  INVX1 U220 ( .A(n337), .Y(n65) );
  AOI22X1 U221 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  OAI221XL U222 ( .A0(n65), .A1(n551), .B0(n31), .B1(n536), .C0(n149), .Y(n143) );
  OAI221XL U223 ( .A0(n145), .A1(n545), .B0(n28), .B1(n551), .C0(n146), .Y(
        n144) );
  AOI2BB2X1 U224 ( .B0(n539), .B1(n87), .A0N(n545), .A1N(n121), .Y(n149) );
  INVX1 U225 ( .A(n208), .Y(n29) );
  INVX1 U226 ( .A(n299), .Y(n11) );
  INVX1 U227 ( .A(n100), .Y(n33) );
  AOI221XL U228 ( .A0(n556), .A1(n52), .B0(n548), .B1(n123), .C0(n324), .Y(
        n316) );
  INVX1 U229 ( .A(n326), .Y(n52) );
  OAI32X1 U230 ( .A0(n94), .A1(n63), .A2(n325), .B0(n37), .B1(n551), .Y(n324)
         );
  INVX1 U231 ( .A(n196), .Y(n31) );
  OAI221XL U232 ( .A0(n56), .A1(n545), .B0(n32), .B1(n94), .C0(n163), .Y(n151)
         );
  INVX1 U233 ( .A(n167), .Y(n32) );
  AOI22X1 U234 ( .A0(n164), .A1(n556), .B0(n129), .B1(n553), .Y(n163) );
  INVX1 U235 ( .A(n141), .Y(n27) );
  INVX1 U236 ( .A(n148), .Y(n28) );
  OAI221XL U237 ( .A0(n40), .A1(n551), .B0(n58), .B1(n545), .C0(n137), .Y(n136) );
  INVX1 U238 ( .A(n96), .Y(n40) );
  AOI31X1 U239 ( .A0(n102), .A1(n138), .A2(n556), .B0(n8), .Y(n137) );
  INVX1 U240 ( .A(n89), .Y(n8) );
  INVX1 U241 ( .A(n185), .Y(n19) );
  INVX1 U242 ( .A(n540), .Y(n543) );
  AOI211X1 U243 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U244 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U245 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  OAI2BB1X1 U246 ( .A0N(n133), .A1N(n134), .B0(n534), .Y(n132) );
  AOI22X1 U247 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  AOI22X1 U248 ( .A0(n171), .A1(n21), .B0(n534), .B1(n172), .Y(n170) );
  OAI221XL U249 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  OAI221XL U250 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  AOI22X1 U251 ( .A0(n533), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U252 ( .A0(n61), .A1(n551), .B0(n545), .B1(n260), .C0(n261), .Y(
        n254) );
  OAI221XL U253 ( .A0(n41), .A1(n545), .B0(n94), .B1(n181), .C0(n256), .Y(n255) );
  AOI21X1 U254 ( .A0(n33), .A1(n16), .B0(n262), .Y(n261) );
  AOI22X1 U255 ( .A0(n348), .A1(n26), .B0(n533), .B1(n349), .Y(n342) );
  OAI221XL U256 ( .A0(n536), .A1(n166), .B0(n286), .B1(n545), .C0(n351), .Y(
        n348) );
  OAI211X1 U257 ( .A0(n88), .A1(n550), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U258 ( .B0(n539), .B1(n196), .A0N(n550), .A1N(n179), .Y(n351) );
  OAI22X1 U259 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U260 ( .A0(n549), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U261 ( .A0(n56), .A1(n4), .B0(n547), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U262 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U263 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U264 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U265 ( .A0(n61), .A1(n552), .B0(n547), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U266 ( .A0(n543), .A1(n71), .B0(n37), .B1(n550), .Y(n157) );
  OAI22X1 U267 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U268 ( .A0(n549), .A1(n111), .B0(n47), .B1(n540), .C0(n112), .Y(
        n109) );
  AOI221X1 U269 ( .A0(n556), .A1(n115), .B0(n553), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U270 ( .A0(n536), .A1(n113), .B0(n44), .B1(n551), .C0(n114), .Y(
        n112) );
  AOI211X1 U271 ( .A0(n55), .A1(n556), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U272 ( .A0(n114), .A1(n206), .A2(n273), .B0(n533), .Y(n272) );
  OAI22X1 U273 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U274 ( .B0(n70), .B1(n552), .A0N(n90), .A1N(n545), .Y(n273) );
  AOI22X1 U275 ( .A0(n534), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U276 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  OAI221XL U277 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  AOI2BB2X1 U278 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  OAI221XL U279 ( .A0(n46), .A1(n551), .B0(n545), .B1(n116), .C0(n267), .Y(
        n264) );
  AOI221XL U281 ( .A0(n548), .A1(n247), .B0(n212), .B1(n540), .C0(n266), .Y(
        n265) );
  AOI22X1 U282 ( .A0(n539), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  AOI22X1 U283 ( .A0(n553), .A1(n532), .B0(n539), .B1(n66), .Y(n292) );
  AOI22X1 U284 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U285 ( .A0(n63), .A1(n545), .B0(n541), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U286 ( .A0(n38), .A1(n536), .B0(n545), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U287 ( .A0(n179), .A1(n552), .B0(n180), .Y(n178) );
  AOI22X1 U288 ( .A0(n533), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U289 ( .A0(n43), .A1(n545), .B0(n541), .B1(n34), .C0(n365), .Y(n361) );
  OAI221XL U290 ( .A0(n532), .A1(n120), .B0(n201), .B1(n551), .C0(n363), .Y(
        n362) );
  INVX1 U291 ( .A(n260), .Y(n43) );
  AOI22X1 U292 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  OAI21XL U293 ( .A0(n321), .A1(n536), .B0(n322), .Y(n318) );
  OAI221XL U294 ( .A0(n551), .A1(n113), .B0(n88), .B1(n545), .C0(n320), .Y(
        n319) );
  AOI31X1 U295 ( .A0(n538), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  CLKINVX3 U296 ( .A(n532), .Y(n71) );
  OAI21XL U297 ( .A0(n545), .A1(n537), .B0(n120), .Y(n276) );
  NAND2X1 U298 ( .A(n63), .B(n531), .Y(n168) );
  AOI21X1 U299 ( .A0(n224), .A1(n243), .B0(n545), .Y(n295) );
  INVX1 U300 ( .A(n531), .Y(n74) );
  OAI21XL U301 ( .A0(n73), .A1(n301), .B0(n550), .Y(n323) );
  OAI21XL U302 ( .A0(n73), .A1(n243), .B0(n550), .Y(n245) );
  OAI21XL U303 ( .A0(n536), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U304 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U305 ( .A(n162), .Y(n5) );
  OAI2BB1X1 U306 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI22X1 U307 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  AOI211X1 U308 ( .A0(n39), .A1(n540), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U309 ( .A0(n551), .A1(n116), .B0(n73), .B1(n230), .C0(n545), .C1(
        n102), .Y(n275) );
  AOI211X1 U310 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U311 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI2BB2X1 U312 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  NAND2X1 U313 ( .A(n62), .B(n552), .Y(n287) );
  NOR2BX1 U314 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U315 ( .A(n82), .Y(n536) );
  NAND2X1 U316 ( .A(n73), .B(n20), .Y(n82) );
  OAI221XL U317 ( .A0(n531), .A1(n259), .B0(n543), .B1(n214), .C0(n287), .Y(
        n293) );
  BUFX3 U318 ( .A(n139), .Y(n538) );
  NAND2X1 U319 ( .A(n531), .B(n537), .Y(n139) );
  AOI211X1 U320 ( .A0(n540), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  OAI222X1 U321 ( .A0(n551), .A1(n167), .B0(n339), .B1(n536), .C0(n545), .C1(
        n34), .Y(n338) );
  AOI21X1 U322 ( .A0(n537), .A1(n535), .B0(n65), .Y(n339) );
  AOI211X1 U323 ( .A0(n533), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  OAI221XL U324 ( .A0(n545), .A1(n116), .B0(n321), .B1(n543), .C0(n359), .Y(
        n354) );
  AOI21X1 U325 ( .A0(n356), .A1(n357), .B0(n533), .Y(n355) );
  AOI31X1 U326 ( .A0(n556), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  INVX1 U327 ( .A(n93), .Y(n546) );
  INVX1 U328 ( .A(n83), .Y(n555) );
  INVX1 U329 ( .A(n544), .Y(n541) );
  INVX1 U330 ( .A(n94), .Y(n544) );
  AOI22X1 U331 ( .A0(n533), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U332 ( .A0(n545), .A1(n141), .B0(n551), .B1(n263), .C0(n29), .C1(
        n543), .Y(n277) );
  OAI221XL U333 ( .A0(n31), .A1(n536), .B0(n551), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U334 ( .B0(n88), .B1(n539), .A0N(n545), .A1N(n197), .Y(n279) );
  NAND2X1 U335 ( .A(n224), .B(n301), .Y(n148) );
  NOR2BX1 U336 ( .AN(n263), .B(n61), .Y(n321) );
  AOI21X1 U337 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI22X1 U338 ( .A0(n556), .A1(n66), .B0(n539), .B1(n147), .Y(n146) );
  AOI22X1 U339 ( .A0(n549), .A1(n85), .B0(n41), .B1(n539), .Y(n84) );
  NAND2X1 U340 ( .A(n224), .B(n118), .Y(n208) );
  NAND2X1 U341 ( .A(n263), .B(n337), .Y(n167) );
  AOI21X1 U342 ( .A0(n263), .A1(n182), .B0(n545), .Y(n305) );
  AOI21X1 U343 ( .A0(n111), .A1(n538), .B0(n543), .Y(n203) );
  NAND2X1 U344 ( .A(n16), .B(n531), .Y(n206) );
  XNOR2X1 U345 ( .A(n20), .B(n531), .Y(n185) );
  NAND2X1 U346 ( .A(n539), .B(n537), .Y(n130) );
  XNOR2X1 U347 ( .A(n73), .B(n531), .Y(n161) );
  AOI21X1 U348 ( .A0(n90), .A1(n73), .B0(n556), .Y(n86) );
  AOI221X1 U349 ( .A0(n46), .A1(n540), .B0(n555), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U350 ( .A0(n536), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U351 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  AOI222X1 U352 ( .A0(n549), .A1(n210), .B0(n211), .B1(n212), .C0(n556), .C1(
        n537), .Y(n191) );
  OAI21XL U353 ( .A0(n73), .A1(n214), .B0(n550), .Y(n211) );
  AOI31X1 U354 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U355 ( .A0(n148), .A1(n73), .B0(n29), .B1(n554), .Y(n300) );
  AOI31X1 U356 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U357 ( .A0N(n223), .A1N(n224), .B0(n554), .Y(n220) );
  AOI22X1 U358 ( .A0(n29), .A1(n556), .B0(n222), .B1(n547), .Y(n221) );
  INVX1 U359 ( .A(n93), .Y(n547) );
  INVX1 U360 ( .A(n93), .Y(n549) );
  INVX1 U361 ( .A(n93), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n358) );
  INVX1 U363 ( .A(n83), .Y(n553) );
  INVX1 U364 ( .A(n83), .Y(n554) );
  INVX1 U365 ( .A(n83), .Y(n552) );
  NOR2BX1 U366 ( .AN(n93), .B(n553), .Y(n309) );
  AOI22X1 U367 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U368 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI22X1 U369 ( .A0(n347), .A1(n26), .B0(n556), .B1(n90), .Y(n343) );
  AOI22X1 U370 ( .A0(n250), .A1(n21), .B0(n534), .B1(n251), .Y(n249) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  OAI22X1 U373 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U374 ( .A0(n548), .A1(n230), .B0(n556), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U375 ( .A0(n164), .A1(n547), .B0(a[2]), .B1(n227), .C0(n556), .C1(
        n228), .Y(n226) );
  OAI22X1 U376 ( .A0(n35), .A1(n542), .B0(n550), .B1(n537), .Y(n231) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI21XL U383 ( .A0(n66), .A1(n550), .B0(n259), .Y(n257) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI33X1 U385 ( .A0(n532), .A1(n540), .A2(n19), .B0(n185), .B1(n181), .B2(
        a[2]), .Y(n184) );
  AOI22X1 U386 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U387 ( .A(a[0]), .Y(n75) );
  AOI211X1 U388 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U389 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U390 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U391 ( .A(a[5]), .Y(n533) );
  OAI221XL U392 ( .A0(n536), .A1(n115), .B0(n121), .B1(n545), .C0(n122), .Y(
        n105) );
  AOI22X1 U393 ( .A0(n539), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_5 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n4, n5, n6, n7, n8, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556;

  OAI221X4 U4 ( .A0(n66), .A1(n536), .B0(n61), .B1(n551), .C0(n84), .Y(n81) );
  OAI221X4 U6 ( .A0(n86), .A1(n87), .B0(n88), .B1(n551), .C0(n89), .Y(n80) );
  OAI222X4 U75 ( .A0(n551), .A1(n207), .B0(n181), .B1(n120), .C0(n545), .C1(
        n208), .Y(n204) );
  OAI32X4 U280 ( .A0(n551), .A1(n56), .A2(n53), .B0(n94), .B1(n103), .Y(n366)
         );
  AOI221X1 U1 ( .A0(n65), .A1(a[2]), .B0(n97), .B1(n358), .C0(n4), .Y(n357) );
  INVX1 U2 ( .A(a[7]), .Y(n20) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n103) );
  OAI222X1 U5 ( .A0(n94), .A1(n118), .B0(n119), .B1(n545), .C0(a[4]), .C1(n120), .Y(n117) );
  NAND2X2 U7 ( .A(n531), .B(n532), .Y(n115) );
  NAND2X1 U8 ( .A(n56), .B(n531), .Y(n229) );
  NAND2X2 U9 ( .A(n532), .B(n66), .Y(n181) );
  NAND2X1 U10 ( .A(n39), .B(n531), .Y(n142) );
  NAND2X2 U11 ( .A(n537), .B(n181), .Y(n113) );
  NAND2X2 U12 ( .A(n66), .B(n535), .Y(n116) );
  CLKINVX3 U13 ( .A(n533), .Y(n26) );
  NAND2X2 U14 ( .A(n66), .B(n71), .Y(n138) );
  NAND2X1 U15 ( .A(n531), .B(n181), .Y(n102) );
  CLKINVX3 U16 ( .A(a[2]), .Y(n73) );
  NAND2X1 U17 ( .A(n533), .B(n75), .Y(n110) );
  NAND2X2 U18 ( .A(n75), .B(n26), .Y(n154) );
  NAND2X2 U19 ( .A(a[0]), .B(n26), .Y(n156) );
  CLKINVX3 U20 ( .A(n534), .Y(n21) );
  OAI22X2 U21 ( .A0(n340), .A1(n21), .B0(n534), .B1(n341), .Y(d[0]) );
  OAI22X2 U22 ( .A0(n534), .A1(n280), .B0(n281), .B1(n21), .Y(d[2]) );
  OAI21X2 U23 ( .A0(n76), .A1(n21), .B0(n77), .Y(d[7]) );
  AOI221X1 U24 ( .A0(n24), .A1(n7), .B0(n25), .B1(n105), .C0(n106), .Y(n76) );
  OAI22X2 U25 ( .A0(n534), .A1(n215), .B0(n216), .B1(n21), .Y(d[4]) );
  OAI21X2 U26 ( .A0(n534), .A1(n131), .B0(n132), .Y(d[6]) );
  AOI221X1 U27 ( .A0(n23), .A1(n150), .B0(n22), .B1(n151), .C0(n152), .Y(n131)
         );
  NAND2X1 U28 ( .A(a[2]), .B(n20), .Y(n83) );
  NAND2X1 U29 ( .A(a[7]), .B(n73), .Y(n93) );
  AOI21XL U30 ( .A0(n4), .A1(a[4]), .B0(n15), .Y(n320) );
  NAND2X1 U31 ( .A(a[4]), .B(n535), .Y(n263) );
  NAND2X1 U32 ( .A(n531), .B(a[4]), .Y(n224) );
  NAND2X2 U33 ( .A(n532), .B(a[4]), .Y(n111) );
  CLKINVX3 U34 ( .A(a[4]), .Y(n66) );
  CLKINVX3 U35 ( .A(n542), .Y(n540) );
  NAND2X1 U36 ( .A(n53), .B(n16), .Y(n288) );
  INVX1 U37 ( .A(n325), .Y(n34) );
  NAND2X1 U38 ( .A(n113), .B(n535), .Y(n214) );
  CLKINVX3 U39 ( .A(n555), .Y(n550) );
  NAND2X1 U40 ( .A(n56), .B(n535), .Y(n233) );
  NAND2X1 U41 ( .A(n50), .B(n535), .Y(n301) );
  NAND2X1 U42 ( .A(n538), .B(n268), .Y(n212) );
  NAND2X1 U43 ( .A(n115), .B(n209), .Y(n210) );
  NAND2X1 U44 ( .A(n147), .B(n214), .Y(n207) );
  INVX1 U45 ( .A(n168), .Y(n62) );
  INVX1 U46 ( .A(n538), .Y(n53) );
  INVX1 U47 ( .A(n182), .Y(n57) );
  NOR2X1 U48 ( .A(n535), .B(n39), .Y(n325) );
  NAND2X1 U49 ( .A(n535), .B(n71), .Y(n118) );
  NAND2X1 U50 ( .A(n138), .B(n535), .Y(n223) );
  NAND2X1 U51 ( .A(n39), .B(n535), .Y(n248) );
  NAND2X1 U52 ( .A(n181), .B(n535), .Y(n166) );
  NAND2X1 U53 ( .A(n229), .B(n248), .Y(n87) );
  INVX1 U54 ( .A(n102), .Y(n61) );
  NAND2X1 U55 ( .A(n115), .B(n223), .Y(n306) );
  INVX1 U56 ( .A(n230), .Y(n69) );
  INVX1 U57 ( .A(n116), .Y(n64) );
  INVX1 U58 ( .A(n103), .Y(n68) );
  BUFX3 U59 ( .A(n74), .Y(n535) );
  NAND2X1 U60 ( .A(n50), .B(n531), .Y(n147) );
  NAND2X1 U61 ( .A(n531), .B(n539), .Y(n120) );
  NAND2X1 U62 ( .A(n111), .B(n535), .Y(n268) );
  NAND2X1 U63 ( .A(n531), .B(n113), .Y(n165) );
  NAND2X1 U64 ( .A(n531), .B(n138), .Y(n182) );
  INVX1 U65 ( .A(n312), .Y(d[1]) );
  INVX1 U66 ( .A(n170), .Y(d[5]) );
  NAND2X1 U67 ( .A(n16), .B(n532), .Y(n259) );
  INVX1 U68 ( .A(n537), .Y(n46) );
  NAND2X1 U69 ( .A(n111), .B(n147), .Y(n96) );
  NOR2X1 U70 ( .A(n537), .B(n535), .Y(n124) );
  CLKINVX3 U71 ( .A(n111), .Y(n39) );
  NAND2X1 U72 ( .A(n531), .B(n71), .Y(n230) );
  NAND2X1 U73 ( .A(n531), .B(n66), .Y(n337) );
  NAND2BX1 U74 ( .AN(n124), .B(n263), .Y(n196) );
  INVX1 U76 ( .A(n156), .Y(n24) );
  NAND2X1 U77 ( .A(n224), .B(n268), .Y(n141) );
  NAND2BX1 U78 ( .AN(n93), .B(n537), .Y(n299) );
  NAND2X1 U79 ( .A(n224), .B(n233), .Y(n104) );
  NAND2X1 U80 ( .A(n263), .B(n142), .Y(n100) );
  CLKINVX3 U81 ( .A(n108), .Y(n22) );
  BUFX3 U82 ( .A(a[1]), .Y(n531) );
  NAND2X1 U83 ( .A(a[7]), .B(a[2]), .Y(n94) );
  INVX1 U84 ( .A(n249), .Y(d[3]) );
  NAND2X1 U85 ( .A(n533), .B(a[0]), .Y(n108) );
  INVX1 U86 ( .A(n238), .Y(n15) );
  NAND2X1 U87 ( .A(n59), .B(n540), .Y(n114) );
  NAND2X1 U88 ( .A(n51), .B(n556), .Y(n238) );
  INVX1 U89 ( .A(n288), .Y(n14) );
  NOR2X1 U90 ( .A(n550), .B(n325), .Y(n199) );
  NOR2X1 U91 ( .A(n49), .B(n62), .Y(n247) );
  NAND2X1 U92 ( .A(n222), .B(n540), .Y(n162) );
  INVX1 U93 ( .A(n301), .Y(n49) );
  INVX1 U94 ( .A(n248), .Y(n37) );
  INVX1 U95 ( .A(n166), .Y(n60) );
  INVX1 U96 ( .A(n207), .Y(n48) );
  INVX1 U97 ( .A(n228), .Y(n51) );
  INVX1 U98 ( .A(n210), .Y(n44) );
  INVX4 U99 ( .A(n536), .Y(n556) );
  NOR2BX1 U100 ( .AN(n214), .B(n69), .Y(n88) );
  NOR2X1 U101 ( .A(n53), .B(n70), .Y(n326) );
  NOR2X1 U102 ( .A(n50), .B(n61), .Y(n286) );
  NAND2X1 U103 ( .A(n34), .B(n223), .Y(n183) );
  INVX1 U104 ( .A(n118), .Y(n70) );
  NAND2X1 U105 ( .A(n34), .B(n248), .Y(n123) );
  INVX1 U106 ( .A(n233), .Y(n55) );
  INVX1 U107 ( .A(n223), .Y(n59) );
  NOR2X1 U108 ( .A(n57), .B(n55), .Y(n197) );
  OAI221XL U109 ( .A0(n58), .A1(n545), .B0(n98), .B1(n543), .C0(n18), .Y(n347)
         );
  INVX1 U110 ( .A(n199), .Y(n18) );
  INVX1 U111 ( .A(n127), .Y(n35) );
  NOR2X1 U112 ( .A(n59), .B(n69), .Y(n98) );
  INVX1 U113 ( .A(n212), .Y(n41) );
  NOR2X1 U114 ( .A(n62), .B(n55), .Y(n145) );
  INVX1 U115 ( .A(n306), .Y(n58) );
  INVX1 U116 ( .A(n158), .Y(n42) );
  INVX1 U117 ( .A(n87), .Y(n38) );
  NAND2X1 U118 ( .A(n63), .B(n535), .Y(n243) );
  NAND2X1 U119 ( .A(n46), .B(n535), .Y(n209) );
  OAI22X1 U120 ( .A0(n240), .A1(n110), .B0(n241), .B1(n154), .Y(n236) );
  AOI222X1 U121 ( .A0(n61), .A1(n548), .B0(n556), .B1(n244), .C0(n245), .C1(
        n212), .Y(n240) );
  AOI211X1 U122 ( .A0(n556), .A1(n234), .B0(n242), .C0(n199), .Y(n241) );
  NAND2X1 U123 ( .A(n116), .B(n229), .Y(n244) );
  NOR2X1 U124 ( .A(n46), .B(n57), .Y(n222) );
  OAI22X1 U125 ( .A0(n542), .A1(n207), .B0(n545), .B1(n538), .Y(n242) );
  CLKINVX3 U126 ( .A(n113), .Y(n50) );
  NAND2X1 U127 ( .A(n214), .B(n142), .Y(n90) );
  CLKINVX3 U128 ( .A(n181), .Y(n63) );
  AOI22X1 U129 ( .A0(n24), .A1(n91), .B0(n23), .B1(n92), .Y(n78) );
  OAI221XL U130 ( .A0(n98), .A1(n545), .B0(n30), .B1(n541), .C0(n99), .Y(n91)
         );
  OAI221XL U131 ( .A0(n42), .A1(n545), .B0(n51), .B1(n542), .C0(n95), .Y(n92)
         );
  INVX1 U132 ( .A(n104), .Y(n30) );
  NAND2X1 U133 ( .A(n556), .B(n96), .Y(n187) );
  NAND2X1 U134 ( .A(n115), .B(n214), .Y(n228) );
  AOI22X1 U135 ( .A0(n23), .A1(n194), .B0(n22), .B1(n195), .Y(n193) );
  OAI221XL U136 ( .A0(n46), .A1(n551), .B0(n63), .B1(n545), .C0(n200), .Y(n194) );
  OAI221XL U137 ( .A0(n536), .A1(n196), .B0(n197), .B1(n545), .C0(n198), .Y(
        n195) );
  AOI211X1 U138 ( .A0(n201), .A1(n556), .B0(n202), .C0(n203), .Y(n200) );
  AOI22X1 U139 ( .A0(n23), .A1(n331), .B0(n22), .B1(n332), .Y(n330) );
  OAI221XL U140 ( .A0(n35), .A1(n545), .B0(n44), .B1(n542), .C0(n333), .Y(n332) );
  OAI211X1 U141 ( .A0(n326), .A1(n550), .B0(n288), .C0(n334), .Y(n331) );
  AOI22X1 U142 ( .A0(n35), .A1(n16), .B0(n39), .B1(n553), .Y(n333) );
  AOI22X1 U143 ( .A0(n548), .A1(n63), .B0(n247), .B1(n539), .Y(n334) );
  AOI21X1 U144 ( .A0(n115), .A1(n243), .B0(n550), .Y(n360) );
  INVX1 U145 ( .A(n120), .Y(n4) );
  AND2X2 U146 ( .A(n165), .B(n166), .Y(n129) );
  NAND2X1 U147 ( .A(n538), .B(n214), .Y(n126) );
  OAI21XL U148 ( .A0(n165), .A1(n550), .B0(n187), .Y(n266) );
  INVX1 U149 ( .A(n284), .Y(n10) );
  OAI31X1 U150 ( .A0(n202), .A1(n14), .A2(n285), .B0(n25), .Y(n284) );
  OAI21XL U151 ( .A0(n541), .A1(n286), .B0(n287), .Y(n285) );
  INVX1 U152 ( .A(n147), .Y(n47) );
  OAI22X1 U153 ( .A0(n302), .A1(n154), .B0(n303), .B1(n110), .Y(n297) );
  AOI211X1 U154 ( .A0(n556), .A1(n102), .B0(n304), .C0(n305), .Y(n303) );
  AOI221X1 U155 ( .A0(n11), .A1(n535), .B0(n27), .B1(n556), .C0(n307), .Y(n302) );
  OAI22X1 U156 ( .A0(n64), .A1(n542), .B0(n550), .B1(n306), .Y(n304) );
  AOI222X1 U157 ( .A0(n56), .A1(n540), .B0(n60), .B1(n552), .C0(n547), .C1(n71), .Y(n356) );
  AOI21X1 U158 ( .A0(n50), .A1(n556), .B0(n366), .Y(n365) );
  OAI221XL U159 ( .A0(n551), .A1(n87), .B0(n543), .B1(n104), .C0(n246), .Y(
        n235) );
  AOI2BB2X1 U160 ( .B0(n11), .B1(n535), .A0N(n536), .A1N(n247), .Y(n246) );
  CLKINVX8 U161 ( .A(n546), .Y(n545) );
  CLKINVX3 U162 ( .A(n541), .Y(n539) );
  NOR2X1 U163 ( .A(n545), .B(n535), .Y(n202) );
  AOI211X1 U164 ( .A0(n45), .A1(n540), .B0(n204), .C0(n205), .Y(n192) );
  INVX1 U165 ( .A(n209), .Y(n45) );
  NAND2BX1 U166 ( .AN(n97), .B(n206), .Y(n205) );
  AOI222X1 U167 ( .A0(n4), .A1(n113), .B0(n199), .B1(n50), .C0(n37), .C1(n540), 
        .Y(n198) );
  AOI221X1 U168 ( .A0(n321), .A1(n554), .B0(n540), .B1(n311), .C0(n327), .Y(
        n315) );
  OAI221XL U169 ( .A0(n536), .A1(n209), .B0(n545), .B1(n103), .C0(n288), .Y(
        n327) );
  AOI221X1 U170 ( .A0(n4), .A1(n71), .B0(n554), .B1(n113), .C0(n186), .Y(n174)
         );
  OAI2BB1X1 U171 ( .A0N(n142), .A1N(n547), .B0(n187), .Y(n186) );
  OAI221XL U172 ( .A0(n308), .A1(n551), .B0(n545), .B1(n165), .C0(n162), .Y(
        n307) );
  NOR2X1 U173 ( .A(n69), .B(n68), .Y(n308) );
  OAI221XL U174 ( .A0(n54), .A1(n545), .B0(n33), .B1(n94), .C0(n232), .Y(n217)
         );
  INVX1 U175 ( .A(n234), .Y(n54) );
  AOI32X1 U176 ( .A0(n34), .A1(n181), .A2(n556), .B0(n554), .B1(n233), .Y(n232) );
  OAI221XL U177 ( .A0(n67), .A1(n551), .B0(n541), .B1(n538), .C0(n294), .Y(
        n282) );
  INVX1 U178 ( .A(n115), .Y(n67) );
  AOI211X1 U179 ( .A0(n48), .A1(n556), .B0(n6), .C0(n295), .Y(n294) );
  INVX1 U180 ( .A(n114), .Y(n6) );
  AOI211X1 U181 ( .A0(n60), .A1(n540), .B0(n13), .C0(n364), .Y(n363) );
  NOR3X1 U182 ( .A(n545), .B(n39), .C(n61), .Y(n364) );
  INVX1 U183 ( .A(n259), .Y(n13) );
  OAI221XL U184 ( .A0(n536), .A1(n168), .B0(n164), .B1(n551), .C0(n169), .Y(
        n150) );
  AOI22X1 U185 ( .A0(n549), .A1(n34), .B0(n48), .B1(n539), .Y(n169) );
  AOI211X1 U186 ( .A0(n554), .A1(n96), .B0(n14), .C0(n97), .Y(n95) );
  CLKINVX3 U187 ( .A(n555), .Y(n551) );
  INVX1 U188 ( .A(n544), .Y(n542) );
  INVX1 U189 ( .A(n125), .Y(n7) );
  AOI221X1 U190 ( .A0(n126), .A1(n553), .B0(n127), .B1(n549), .C0(n128), .Y(
        n125) );
  OAI21XL U191 ( .A0(n536), .A1(n129), .B0(n130), .Y(n128) );
  INVX1 U192 ( .A(n536), .Y(n16) );
  NOR2X1 U193 ( .A(n39), .B(n57), .Y(n179) );
  CLKINVX3 U194 ( .A(n110), .Y(n23) );
  NAND3X1 U195 ( .A(n538), .B(n113), .C(n540), .Y(n89) );
  NAND2X1 U196 ( .A(n116), .B(n142), .Y(n85) );
  NAND2X1 U197 ( .A(n115), .B(n268), .Y(n158) );
  NAND2X1 U198 ( .A(n538), .B(n166), .Y(n311) );
  NOR2BX1 U199 ( .AN(n229), .B(n68), .Y(n164) );
  AOI21X1 U200 ( .A0(n181), .A1(n182), .B0(n536), .Y(n180) );
  OAI221XL U201 ( .A0(n36), .A1(n550), .B0(n121), .B1(n541), .C0(n140), .Y(
        n135) );
  INVX1 U202 ( .A(n85), .Y(n36) );
  AOI22X1 U203 ( .A0(n49), .A1(n548), .B0(n556), .B1(n141), .Y(n140) );
  AOI22X1 U204 ( .A0(n57), .A1(n546), .B0(n552), .B1(n113), .Y(n239) );
  AOI22X1 U205 ( .A0(n547), .A1(n311), .B0(n50), .B1(n539), .Y(n350) );
  NOR2X1 U206 ( .A(n138), .B(n536), .Y(n97) );
  NAND2X1 U207 ( .A(n243), .B(n142), .Y(n127) );
  INVX1 U208 ( .A(n154), .Y(n25) );
  NAND2X1 U209 ( .A(n229), .B(n243), .Y(n234) );
  CLKINVX3 U210 ( .A(n138), .Y(n56) );
  NAND2X1 U211 ( .A(n229), .B(n209), .Y(n260) );
  NOR2X1 U212 ( .A(n64), .B(n124), .Y(n121) );
  AOI211X1 U213 ( .A0(n556), .A1(n306), .B0(n335), .C0(n336), .Y(n329) );
  OAI2BB2X1 U214 ( .B0(n545), .B1(n183), .A0N(n188), .A1N(n540), .Y(n335) );
  AOI21X1 U215 ( .A0(n301), .A1(n337), .B0(n550), .Y(n336) );
  NAND2X1 U216 ( .A(n138), .B(n102), .Y(n227) );
  NAND2X1 U217 ( .A(n103), .B(n165), .Y(n188) );
  AOI21X1 U218 ( .A0(n556), .A1(n100), .B0(n101), .Y(n99) );
  AOI21X1 U219 ( .A0(n102), .A1(n103), .B0(n550), .Y(n101) );
  INVX1 U220 ( .A(n337), .Y(n65) );
  AOI22X1 U221 ( .A0(n24), .A1(n143), .B0(n22), .B1(n144), .Y(n133) );
  OAI221XL U222 ( .A0(n65), .A1(n551), .B0(n31), .B1(n536), .C0(n149), .Y(n143) );
  OAI221XL U223 ( .A0(n145), .A1(n545), .B0(n28), .B1(n551), .C0(n146), .Y(
        n144) );
  AOI2BB2X1 U224 ( .B0(n539), .B1(n87), .A0N(n545), .A1N(n121), .Y(n149) );
  INVX1 U225 ( .A(n208), .Y(n29) );
  INVX1 U226 ( .A(n299), .Y(n11) );
  INVX1 U227 ( .A(n100), .Y(n33) );
  AOI221XL U228 ( .A0(n556), .A1(n52), .B0(n548), .B1(n123), .C0(n324), .Y(
        n316) );
  INVX1 U229 ( .A(n326), .Y(n52) );
  OAI32X1 U230 ( .A0(n94), .A1(n63), .A2(n325), .B0(n37), .B1(n551), .Y(n324)
         );
  INVX1 U231 ( .A(n196), .Y(n31) );
  OAI221XL U232 ( .A0(n56), .A1(n545), .B0(n32), .B1(n94), .C0(n163), .Y(n151)
         );
  INVX1 U233 ( .A(n167), .Y(n32) );
  AOI22X1 U234 ( .A0(n164), .A1(n556), .B0(n129), .B1(n553), .Y(n163) );
  INVX1 U235 ( .A(n141), .Y(n27) );
  INVX1 U236 ( .A(n148), .Y(n28) );
  OAI221XL U237 ( .A0(n40), .A1(n551), .B0(n58), .B1(n545), .C0(n137), .Y(n136) );
  INVX1 U238 ( .A(n96), .Y(n40) );
  AOI31X1 U239 ( .A0(n102), .A1(n138), .A2(n556), .B0(n8), .Y(n137) );
  INVX1 U240 ( .A(n89), .Y(n8) );
  INVX1 U241 ( .A(n185), .Y(n19) );
  INVX1 U242 ( .A(n540), .Y(n543) );
  AOI211X1 U243 ( .A0(n22), .A1(n235), .B0(n236), .C0(n237), .Y(n215) );
  AOI211X1 U244 ( .A0(n23), .A1(n217), .B0(n218), .C0(n219), .Y(n216) );
  AOI31X1 U245 ( .A0(n238), .A1(n130), .A2(n239), .B0(n156), .Y(n237) );
  OAI2BB1X1 U246 ( .A0N(n133), .A1N(n134), .B0(n534), .Y(n132) );
  AOI22X1 U247 ( .A0(n23), .A1(n135), .B0(n25), .B1(n136), .Y(n134) );
  AOI22X1 U248 ( .A0(n171), .A1(n21), .B0(n534), .B1(n172), .Y(n170) );
  OAI221XL U249 ( .A0(n173), .A1(n108), .B0(n174), .B1(n154), .C0(n175), .Y(
        n172) );
  OAI221XL U250 ( .A0(n191), .A1(n154), .B0(n192), .B1(n156), .C0(n193), .Y(
        n171) );
  AOI22X1 U251 ( .A0(n533), .A1(n254), .B0(n255), .B1(n26), .Y(n253) );
  OAI221XL U252 ( .A0(n61), .A1(n551), .B0(n545), .B1(n260), .C0(n261), .Y(
        n254) );
  OAI221XL U253 ( .A0(n41), .A1(n545), .B0(n94), .B1(n181), .C0(n256), .Y(n255) );
  AOI21X1 U254 ( .A0(n33), .A1(n16), .B0(n262), .Y(n261) );
  AOI22X1 U255 ( .A0(n348), .A1(n26), .B0(n533), .B1(n349), .Y(n342) );
  OAI221XL U256 ( .A0(n536), .A1(n166), .B0(n286), .B1(n545), .C0(n351), .Y(
        n348) );
  OAI211X1 U257 ( .A0(n88), .A1(n550), .B0(n187), .C0(n350), .Y(n349) );
  AOI2BB2X1 U258 ( .B0(n539), .B1(n196), .A0N(n550), .A1N(n179), .Y(n351) );
  OAI22X1 U259 ( .A0(n289), .A1(n110), .B0(n290), .B1(n156), .Y(n283) );
  AOI221XL U260 ( .A0(n549), .A1(n183), .B0(n124), .B1(n73), .C0(n291), .Y(
        n290) );
  AOI221XL U261 ( .A0(n56), .A1(n4), .B0(n547), .B1(n210), .C0(n293), .Y(n289)
         );
  OAI32X1 U262 ( .A0(n185), .A1(n63), .A2(n73), .B0(n292), .B1(n19), .Y(n291)
         );
  OAI22X1 U263 ( .A0(n153), .A1(n154), .B0(n155), .B1(n156), .Y(n152) );
  AOI211X1 U264 ( .A0(n42), .A1(n73), .B0(n157), .C0(n15), .Y(n155) );
  AOI221XL U265 ( .A0(n61), .A1(n552), .B0(n547), .B1(n147), .C0(n159), .Y(
        n153) );
  OAI22X1 U266 ( .A0(n543), .A1(n71), .B0(n37), .B1(n550), .Y(n157) );
  OAI22X1 U267 ( .A0(n107), .A1(n108), .B0(n109), .B1(n110), .Y(n106) );
  AOI221XL U268 ( .A0(n549), .A1(n111), .B0(n47), .B1(n540), .C0(n112), .Y(
        n109) );
  AOI221X1 U269 ( .A0(n556), .A1(n115), .B0(n553), .B1(n116), .C0(n117), .Y(
        n107) );
  OAI221XL U270 ( .A0(n536), .A1(n113), .B0(n44), .B1(n551), .C0(n114), .Y(
        n112) );
  AOI211X1 U271 ( .A0(n55), .A1(n556), .B0(n271), .C0(n272), .Y(n270) );
  AOI31X1 U272 ( .A0(n114), .A1(n206), .A2(n273), .B0(n533), .Y(n272) );
  OAI22X1 U273 ( .A0(n66), .A1(n120), .B0(n274), .B1(n26), .Y(n271) );
  AOI2BB2X1 U274 ( .B0(n70), .B1(n552), .A0N(n90), .A1N(n545), .Y(n273) );
  AOI22X1 U275 ( .A0(n534), .A1(n313), .B0(n314), .B1(n21), .Y(n312) );
  OAI221XL U276 ( .A0(n328), .A1(n156), .B0(n329), .B1(n154), .C0(n330), .Y(
        n313) );
  OAI221XL U277 ( .A0(n315), .A1(n156), .B0(n316), .B1(n154), .C0(n317), .Y(
        n314) );
  AOI2BB2X1 U278 ( .B0(n264), .B1(n26), .A0N(n26), .A1N(n265), .Y(n252) );
  OAI221XL U279 ( .A0(n46), .A1(n551), .B0(n545), .B1(n116), .C0(n267), .Y(
        n264) );
  AOI221XL U281 ( .A0(n548), .A1(n247), .B0(n212), .B1(n540), .C0(n266), .Y(
        n265) );
  AOI22X1 U282 ( .A0(n539), .A1(n158), .B0(n50), .B1(n20), .Y(n267) );
  AOI22X1 U283 ( .A0(n553), .A1(n532), .B0(n539), .B1(n66), .Y(n292) );
  AOI22X1 U284 ( .A0(n23), .A1(n176), .B0(n24), .B1(n177), .Y(n175) );
  OAI221XL U285 ( .A0(n63), .A1(n545), .B0(n541), .B1(n116), .C0(n178), .Y(
        n177) );
  OAI221XL U286 ( .A0(n38), .A1(n536), .B0(n545), .B1(n183), .C0(n184), .Y(
        n176) );
  AOI21X1 U287 ( .A0(n179), .A1(n552), .B0(n180), .Y(n178) );
  AOI22X1 U288 ( .A0(n533), .A1(n361), .B0(n362), .B1(n26), .Y(n352) );
  OAI221XL U289 ( .A0(n43), .A1(n545), .B0(n541), .B1(n34), .C0(n365), .Y(n361) );
  OAI221XL U290 ( .A0(n532), .A1(n120), .B0(n201), .B1(n551), .C0(n363), .Y(
        n362) );
  INVX1 U291 ( .A(n260), .Y(n43) );
  AOI22X1 U292 ( .A0(n22), .A1(n318), .B0(n23), .B1(n319), .Y(n317) );
  OAI21XL U293 ( .A0(n321), .A1(n536), .B0(n322), .Y(n318) );
  OAI221XL U294 ( .A0(n551), .A1(n113), .B0(n88), .B1(n545), .C0(n320), .Y(
        n319) );
  AOI31X1 U295 ( .A0(n538), .A1(n181), .A2(n323), .B0(n11), .Y(n322) );
  CLKINVX3 U296 ( .A(n532), .Y(n71) );
  OAI21XL U297 ( .A0(n545), .A1(n537), .B0(n120), .Y(n276) );
  NAND2X1 U298 ( .A(n63), .B(n531), .Y(n168) );
  AOI21X1 U299 ( .A0(n224), .A1(n243), .B0(n545), .Y(n295) );
  INVX1 U300 ( .A(n531), .Y(n74) );
  OAI21XL U301 ( .A0(n73), .A1(n301), .B0(n550), .Y(n323) );
  OAI21XL U302 ( .A0(n73), .A1(n243), .B0(n550), .Y(n245) );
  OAI21XL U303 ( .A0(n536), .A1(n118), .B0(n160), .Y(n159) );
  AOI31X1 U304 ( .A0(n111), .A1(n20), .A2(n161), .B0(n5), .Y(n160) );
  INVX1 U305 ( .A(n162), .Y(n5) );
  OAI2BB1X1 U306 ( .A0N(n78), .A1N(n79), .B0(n21), .Y(n77) );
  AOI22X1 U307 ( .A0(n22), .A1(n80), .B0(n25), .B1(n81), .Y(n79) );
  AOI211X1 U308 ( .A0(n39), .A1(n540), .B0(n275), .C0(n276), .Y(n274) );
  OAI222X1 U309 ( .A0(n551), .A1(n116), .B0(n73), .B1(n230), .C0(n545), .C1(
        n102), .Y(n275) );
  AOI211X1 U310 ( .A0(n22), .A1(n296), .B0(n297), .C0(n298), .Y(n280) );
  AOI211X1 U311 ( .A0(n22), .A1(n282), .B0(n283), .C0(n10), .Y(n281) );
  OAI2BB2X1 U312 ( .B0(n309), .B1(n310), .A0N(n179), .A1N(n309), .Y(n296) );
  NAND2X1 U313 ( .A(n62), .B(n552), .Y(n287) );
  NOR2BX1 U314 ( .AN(n263), .B(n47), .Y(n201) );
  BUFX3 U315 ( .A(n82), .Y(n536) );
  NAND2X1 U316 ( .A(n73), .B(n20), .Y(n82) );
  OAI221XL U317 ( .A0(n531), .A1(n259), .B0(n543), .B1(n214), .C0(n287), .Y(
        n293) );
  BUFX3 U318 ( .A(n139), .Y(n538) );
  NAND2X1 U319 ( .A(n531), .B(n537), .Y(n139) );
  AOI211X1 U320 ( .A0(n540), .A1(n71), .B0(n338), .C0(n276), .Y(n328) );
  OAI222X1 U321 ( .A0(n551), .A1(n167), .B0(n339), .B1(n536), .C0(n545), .C1(
        n34), .Y(n338) );
  AOI21X1 U322 ( .A0(n537), .A1(n535), .B0(n65), .Y(n339) );
  AOI211X1 U323 ( .A0(n533), .A1(n354), .B0(n75), .C0(n355), .Y(n353) );
  OAI221XL U324 ( .A0(n545), .A1(n116), .B0(n321), .B1(n543), .C0(n359), .Y(
        n354) );
  AOI21X1 U325 ( .A0(n356), .A1(n357), .B0(n533), .Y(n355) );
  AOI31X1 U326 ( .A0(n556), .A1(n358), .A2(n39), .B0(n360), .Y(n359) );
  INVX1 U327 ( .A(n93), .Y(n546) );
  INVX1 U328 ( .A(n83), .Y(n555) );
  INVX1 U329 ( .A(n544), .Y(n541) );
  INVX1 U330 ( .A(n94), .Y(n544) );
  AOI22X1 U331 ( .A0(n533), .A1(n277), .B0(n278), .B1(n26), .Y(n269) );
  OAI222X1 U332 ( .A0(n545), .A1(n141), .B0(n551), .B1(n263), .C0(n29), .C1(
        n543), .Y(n277) );
  OAI221XL U333 ( .A0(n31), .A1(n536), .B0(n551), .B1(n104), .C0(n279), .Y(
        n278) );
  AOI2BB2X1 U334 ( .B0(n88), .B1(n539), .A0N(n545), .A1N(n197), .Y(n279) );
  NAND2X1 U335 ( .A(n224), .B(n301), .Y(n148) );
  NOR2BX1 U336 ( .AN(n263), .B(n61), .Y(n321) );
  AOI21X1 U337 ( .A0(n233), .A1(n165), .B0(n20), .Y(n262) );
  AOI22X1 U338 ( .A0(n556), .A1(n66), .B0(n539), .B1(n147), .Y(n146) );
  AOI22X1 U339 ( .A0(n549), .A1(n85), .B0(n41), .B1(n539), .Y(n84) );
  NAND2X1 U340 ( .A(n224), .B(n118), .Y(n208) );
  NAND2X1 U341 ( .A(n263), .B(n337), .Y(n167) );
  AOI21X1 U342 ( .A0(n263), .A1(n182), .B0(n545), .Y(n305) );
  AOI21X1 U343 ( .A0(n111), .A1(n538), .B0(n543), .Y(n203) );
  NAND2X1 U344 ( .A(n16), .B(n531), .Y(n206) );
  XNOR2X1 U345 ( .A(n20), .B(n531), .Y(n185) );
  NAND2X1 U346 ( .A(n539), .B(n537), .Y(n130) );
  XNOR2X1 U347 ( .A(n73), .B(n531), .Y(n161) );
  AOI21X1 U348 ( .A0(n90), .A1(n73), .B0(n556), .Y(n86) );
  AOI221X1 U349 ( .A0(n46), .A1(n540), .B0(n555), .B1(n188), .C0(n189), .Y(
        n173) );
  AOI21X1 U350 ( .A0(n536), .A1(n190), .B0(n124), .Y(n189) );
  OAI21XL U351 ( .A0(n62), .A1(n70), .B0(n73), .Y(n190) );
  AOI222X1 U352 ( .A0(n549), .A1(n210), .B0(n211), .B1(n212), .C0(n556), .C1(
        n537), .Y(n191) );
  OAI21XL U353 ( .A0(n73), .A1(n214), .B0(n550), .Y(n211) );
  AOI31X1 U354 ( .A0(n162), .A1(n299), .A2(n300), .B0(n156), .Y(n298) );
  AOI22X1 U355 ( .A0(n148), .A1(n73), .B0(n29), .B1(n554), .Y(n300) );
  AOI31X1 U356 ( .A0(n220), .A1(n130), .A2(n221), .B0(n108), .Y(n219) );
  OAI2BB1X1 U357 ( .A0N(n223), .A1N(n224), .B0(n554), .Y(n220) );
  AOI22X1 U358 ( .A0(n29), .A1(n556), .B0(n222), .B1(n547), .Y(n221) );
  INVX1 U359 ( .A(n93), .Y(n547) );
  INVX1 U360 ( .A(n93), .Y(n549) );
  INVX1 U361 ( .A(n93), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n358) );
  INVX1 U363 ( .A(n83), .Y(n553) );
  INVX1 U364 ( .A(n83), .Y(n554) );
  INVX1 U365 ( .A(n83), .Y(n552) );
  NOR2BX1 U366 ( .AN(n93), .B(n553), .Y(n309) );
  AOI22X1 U367 ( .A0(n342), .A1(a[0]), .B0(n343), .B1(n344), .Y(n341) );
  AOI31X1 U368 ( .A0(n206), .A1(n75), .A2(n352), .B0(n353), .Y(n340) );
  AOI22X1 U369 ( .A0(n347), .A1(n26), .B0(n556), .B1(n90), .Y(n343) );
  AOI22X1 U370 ( .A0(n250), .A1(n21), .B0(n534), .B1(n251), .Y(n249) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n269), .B0(n270), .B1(n75), .Y(n250) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n252), .B0(n253), .B1(n75), .Y(n251) );
  OAI22X1 U373 ( .A0(n225), .A1(n156), .B0(n226), .B1(n154), .Y(n218) );
  AOI221X1 U374 ( .A0(n548), .A1(n230), .B0(n556), .B1(n126), .C0(n231), .Y(
        n225) );
  AOI222X1 U375 ( .A0(n164), .A1(n547), .B0(a[2]), .B1(n227), .C0(n556), .C1(
        n228), .Y(n226) );
  OAI22X1 U376 ( .A0(n35), .A1(n542), .B0(n550), .B1(n537), .Y(n231) );
  NOR2X1 U377 ( .A(n60), .B(n62), .Y(n119) );
  BUFX3 U378 ( .A(n213), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n71), .Y(n213) );
  AOI221X1 U380 ( .A0(n4), .A1(n138), .B0(n72), .B1(n257), .C0(n258), .Y(n256)
         );
  NOR3X1 U381 ( .A(n72), .B(a[7]), .C(n63), .Y(n258) );
  INVX1 U382 ( .A(n161), .Y(n72) );
  OAI21XL U383 ( .A0(n66), .A1(n550), .B0(n259), .Y(n257) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI33X1 U385 ( .A0(n532), .A1(n540), .A2(n19), .B0(n185), .B1(n181), .B2(
        a[2]), .Y(n184) );
  AOI22X1 U386 ( .A0(n41), .A1(n73), .B0(a[2]), .B1(n311), .Y(n310) );
  CLKINVX3 U387 ( .A(a[0]), .Y(n75) );
  AOI211X1 U388 ( .A0(n199), .A1(n345), .B0(n346), .C0(a[0]), .Y(n344) );
  NAND2X1 U389 ( .A(n142), .B(n118), .Y(n345) );
  AOI21X1 U390 ( .A0(n120), .A1(n299), .B0(n26), .Y(n346) );
  BUFX3 U391 ( .A(a[5]), .Y(n533) );
  OAI221XL U392 ( .A0(n536), .A1(n115), .B0(n121), .B1(n545), .C0(n122), .Y(
        n105) );
  AOI22X1 U393 ( .A0(n539), .A1(n123), .B0(n124), .B1(a[2]), .Y(n122) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_6 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916;

  OAI221X4 U4 ( .A0(n857), .A1(n536), .B0(n862), .B1(n551), .C0(n839), .Y(n842) );
  OAI221X4 U6 ( .A0(n837), .A1(n836), .B0(n835), .B1(n551), .C0(n834), .Y(n843) );
  OAI222X4 U75 ( .A0(n551), .A1(n716), .B0(n742), .B1(n803), .C0(n545), .C1(
        n715), .Y(n719) );
  OAI32X4 U280 ( .A0(n551), .A1(n867), .A2(n870), .B0(n829), .B1(n820), .Y(
        n557) );
  AOI221X1 U1 ( .A0(n858), .A1(a[2]), .B0(n826), .B1(n565), .C0(n916), .Y(n566) );
  INVX1 U2 ( .A(a[7]), .Y(n903) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n820) );
  OAI222X1 U5 ( .A0(n829), .A1(n805), .B0(n804), .B1(n545), .C0(a[4]), .C1(
        n803), .Y(n806) );
  NAND2X2 U7 ( .A(n531), .B(n532), .Y(n808) );
  NAND2X1 U8 ( .A(n867), .B(n531), .Y(n694) );
  NAND2X2 U9 ( .A(n532), .B(n857), .Y(n742) );
  NAND2X1 U10 ( .A(n884), .B(n531), .Y(n781) );
  NAND2X2 U11 ( .A(n537), .B(n742), .Y(n810) );
  NAND2X2 U12 ( .A(n857), .B(n535), .Y(n807) );
  CLKINVX3 U13 ( .A(n533), .Y(n897) );
  NAND2X2 U14 ( .A(n857), .B(n852), .Y(n785) );
  NAND2X1 U15 ( .A(n531), .B(n742), .Y(n821) );
  CLKINVX3 U16 ( .A(a[2]), .Y(n850) );
  NAND2X1 U17 ( .A(n533), .B(n848), .Y(n813) );
  NAND2X2 U18 ( .A(n848), .B(n897), .Y(n769) );
  NAND2X2 U19 ( .A(a[0]), .B(n897), .Y(n767) );
  CLKINVX3 U20 ( .A(n534), .Y(n902) );
  OAI22X2 U21 ( .A0(n583), .A1(n902), .B0(n534), .B1(n582), .Y(d[0]) );
  OAI22X2 U22 ( .A0(n534), .A1(n643), .B0(n642), .B1(n902), .Y(d[2]) );
  OAI21X2 U23 ( .A0(n847), .A1(n902), .B0(n846), .Y(d[7]) );
  AOI221X1 U24 ( .A0(n899), .A1(n913), .B0(n898), .B1(n818), .C0(n817), .Y(
        n847) );
  OAI22X2 U25 ( .A0(n534), .A1(n708), .B0(n707), .B1(n902), .Y(d[4]) );
  OAI21X2 U26 ( .A0(n534), .A1(n792), .B0(n791), .Y(d[6]) );
  AOI221X1 U27 ( .A0(n900), .A1(n773), .B0(n901), .B1(n772), .C0(n771), .Y(
        n792) );
  NAND2X1 U28 ( .A(a[2]), .B(n903), .Y(n840) );
  NAND2X1 U29 ( .A(a[7]), .B(n850), .Y(n830) );
  AOI21XL U30 ( .A0(n916), .A1(a[4]), .B0(n907), .Y(n603) );
  NAND2X1 U31 ( .A(a[4]), .B(n535), .Y(n660) );
  NAND2X1 U32 ( .A(n531), .B(a[4]), .Y(n699) );
  NAND2X2 U33 ( .A(n532), .B(a[4]), .Y(n812) );
  CLKINVX3 U34 ( .A(a[4]), .Y(n857) );
  CLKINVX3 U35 ( .A(n542), .Y(n540) );
  NAND2X1 U36 ( .A(n870), .B(n906), .Y(n635) );
  INVX1 U37 ( .A(n598), .Y(n889) );
  NAND2X1 U38 ( .A(n810), .B(n535), .Y(n709) );
  CLKINVX3 U39 ( .A(n555), .Y(n550) );
  NAND2X1 U40 ( .A(n867), .B(n535), .Y(n690) );
  NAND2X1 U41 ( .A(n873), .B(n535), .Y(n622) );
  NAND2X1 U42 ( .A(n538), .B(n655), .Y(n711) );
  NAND2X1 U43 ( .A(n808), .B(n714), .Y(n713) );
  NAND2X1 U44 ( .A(n776), .B(n709), .Y(n716) );
  INVX1 U45 ( .A(n755), .Y(n861) );
  INVX1 U46 ( .A(n538), .Y(n870) );
  INVX1 U47 ( .A(n741), .Y(n866) );
  NOR2X1 U48 ( .A(n535), .B(n884), .Y(n598) );
  NAND2X1 U49 ( .A(n535), .B(n852), .Y(n805) );
  NAND2X1 U50 ( .A(n785), .B(n535), .Y(n700) );
  NAND2X1 U51 ( .A(n884), .B(n535), .Y(n675) );
  NAND2X1 U52 ( .A(n742), .B(n535), .Y(n757) );
  NAND2X1 U53 ( .A(n694), .B(n675), .Y(n836) );
  INVX1 U54 ( .A(n821), .Y(n862) );
  NAND2X1 U55 ( .A(n808), .B(n700), .Y(n617) );
  INVX1 U56 ( .A(n693), .Y(n854) );
  INVX1 U57 ( .A(n807), .Y(n859) );
  INVX1 U58 ( .A(n820), .Y(n855) );
  BUFX3 U59 ( .A(n849), .Y(n535) );
  NAND2X1 U60 ( .A(n873), .B(n531), .Y(n776) );
  NAND2X1 U61 ( .A(n531), .B(n539), .Y(n803) );
  NAND2X1 U62 ( .A(n812), .B(n535), .Y(n655) );
  NAND2X1 U63 ( .A(n531), .B(n810), .Y(n758) );
  NAND2X1 U64 ( .A(n531), .B(n785), .Y(n741) );
  INVX1 U65 ( .A(n611), .Y(d[1]) );
  INVX1 U66 ( .A(n753), .Y(d[5]) );
  NAND2X1 U67 ( .A(n906), .B(n532), .Y(n664) );
  INVX1 U68 ( .A(n537), .Y(n877) );
  NAND2X1 U69 ( .A(n812), .B(n776), .Y(n827) );
  NOR2X1 U70 ( .A(n537), .B(n535), .Y(n799) );
  CLKINVX3 U71 ( .A(n812), .Y(n884) );
  NAND2X1 U72 ( .A(n531), .B(n852), .Y(n693) );
  NAND2X1 U73 ( .A(n531), .B(n857), .Y(n586) );
  NAND2BX1 U74 ( .AN(n799), .B(n660), .Y(n727) );
  INVX1 U76 ( .A(n767), .Y(n899) );
  NAND2X1 U77 ( .A(n699), .B(n655), .Y(n782) );
  NAND2BX1 U78 ( .AN(n830), .B(n537), .Y(n624) );
  NAND2X1 U79 ( .A(n699), .B(n690), .Y(n819) );
  NAND2X1 U80 ( .A(n660), .B(n781), .Y(n823) );
  CLKINVX3 U81 ( .A(n815), .Y(n901) );
  BUFX3 U82 ( .A(a[1]), .Y(n531) );
  NAND2X1 U83 ( .A(a[7]), .B(a[2]), .Y(n829) );
  INVX1 U84 ( .A(n674), .Y(d[3]) );
  NAND2X1 U85 ( .A(n533), .B(a[0]), .Y(n815) );
  INVX1 U86 ( .A(n685), .Y(n907) );
  NAND2X1 U87 ( .A(n864), .B(n540), .Y(n809) );
  NAND2X1 U88 ( .A(n872), .B(n556), .Y(n685) );
  INVX1 U89 ( .A(n635), .Y(n908) );
  NOR2X1 U90 ( .A(n550), .B(n598), .Y(n724) );
  NOR2X1 U91 ( .A(n874), .B(n861), .Y(n676) );
  NAND2X1 U92 ( .A(n701), .B(n540), .Y(n761) );
  INVX1 U93 ( .A(n622), .Y(n874) );
  INVX1 U94 ( .A(n675), .Y(n886) );
  INVX1 U95 ( .A(n757), .Y(n863) );
  INVX1 U96 ( .A(n716), .Y(n875) );
  INVX1 U97 ( .A(n695), .Y(n872) );
  INVX1 U98 ( .A(n713), .Y(n879) );
  INVX4 U99 ( .A(n536), .Y(n556) );
  NOR2BX1 U100 ( .AN(n709), .B(n854), .Y(n835) );
  NOR2X1 U101 ( .A(n870), .B(n853), .Y(n597) );
  NOR2X1 U102 ( .A(n873), .B(n862), .Y(n637) );
  NAND2X1 U103 ( .A(n889), .B(n700), .Y(n740) );
  INVX1 U104 ( .A(n805), .Y(n853) );
  NAND2X1 U105 ( .A(n889), .B(n675), .Y(n800) );
  INVX1 U106 ( .A(n690), .Y(n868) );
  INVX1 U107 ( .A(n700), .Y(n864) );
  NOR2X1 U108 ( .A(n866), .B(n868), .Y(n726) );
  OAI221XL U109 ( .A0(n865), .A1(n545), .B0(n825), .B1(n543), .C0(n905), .Y(
        n576) );
  INVX1 U110 ( .A(n724), .Y(n905) );
  INVX1 U111 ( .A(n796), .Y(n888) );
  NOR2X1 U112 ( .A(n864), .B(n854), .Y(n825) );
  INVX1 U113 ( .A(n711), .Y(n882) );
  NOR2X1 U114 ( .A(n861), .B(n868), .Y(n778) );
  INVX1 U115 ( .A(n617), .Y(n865) );
  INVX1 U116 ( .A(n765), .Y(n881) );
  INVX1 U117 ( .A(n836), .Y(n885) );
  NAND2X1 U118 ( .A(n860), .B(n535), .Y(n680) );
  NAND2X1 U119 ( .A(n877), .B(n535), .Y(n714) );
  OAI22X1 U120 ( .A0(n683), .A1(n813), .B0(n682), .B1(n769), .Y(n687) );
  AOI222X1 U121 ( .A0(n862), .A1(n548), .B0(n556), .B1(n679), .C0(n678), .C1(
        n711), .Y(n683) );
  AOI211X1 U122 ( .A0(n556), .A1(n689), .B0(n681), .C0(n724), .Y(n682) );
  NAND2X1 U123 ( .A(n807), .B(n694), .Y(n679) );
  NOR2X1 U124 ( .A(n877), .B(n866), .Y(n701) );
  OAI22X1 U125 ( .A0(n542), .A1(n716), .B0(n545), .B1(n538), .Y(n681) );
  CLKINVX3 U126 ( .A(n810), .Y(n873) );
  NAND2X1 U127 ( .A(n709), .B(n781), .Y(n833) );
  CLKINVX3 U128 ( .A(n742), .Y(n860) );
  AOI22X1 U129 ( .A0(n899), .A1(n832), .B0(n900), .B1(n831), .Y(n845) );
  OAI221XL U130 ( .A0(n825), .A1(n545), .B0(n893), .B1(n541), .C0(n824), .Y(
        n832) );
  OAI221XL U131 ( .A0(n881), .A1(n545), .B0(n872), .B1(n542), .C0(n828), .Y(
        n831) );
  INVX1 U132 ( .A(n819), .Y(n893) );
  NAND2X1 U133 ( .A(n556), .B(n827), .Y(n736) );
  NAND2X1 U134 ( .A(n808), .B(n709), .Y(n695) );
  AOI22X1 U135 ( .A0(n900), .A1(n729), .B0(n901), .B1(n728), .Y(n730) );
  OAI221XL U136 ( .A0(n877), .A1(n551), .B0(n860), .B1(n545), .C0(n723), .Y(
        n729) );
  OAI221XL U137 ( .A0(n536), .A1(n727), .B0(n726), .B1(n545), .C0(n725), .Y(
        n728) );
  AOI211X1 U138 ( .A0(n722), .A1(n556), .B0(n721), .C0(n720), .Y(n723) );
  AOI22X1 U139 ( .A0(n900), .A1(n592), .B0(n901), .B1(n591), .Y(n593) );
  OAI221XL U140 ( .A0(n888), .A1(n545), .B0(n879), .B1(n542), .C0(n590), .Y(
        n591) );
  OAI211X1 U141 ( .A0(n597), .A1(n550), .B0(n635), .C0(n589), .Y(n592) );
  AOI22X1 U142 ( .A0(n888), .A1(n906), .B0(n884), .B1(n553), .Y(n590) );
  AOI22X1 U143 ( .A0(n548), .A1(n860), .B0(n676), .B1(n539), .Y(n589) );
  AOI21X1 U144 ( .A0(n808), .A1(n680), .B0(n550), .Y(n563) );
  INVX1 U145 ( .A(n803), .Y(n916) );
  AND2X2 U146 ( .A(n758), .B(n757), .Y(n794) );
  NAND2X1 U147 ( .A(n538), .B(n709), .Y(n797) );
  OAI21XL U148 ( .A0(n758), .A1(n550), .B0(n736), .Y(n657) );
  INVX1 U149 ( .A(n639), .Y(n911) );
  OAI31X1 U150 ( .A0(n721), .A1(n908), .A2(n638), .B0(n898), .Y(n639) );
  OAI21XL U151 ( .A0(n541), .A1(n637), .B0(n636), .Y(n638) );
  INVX1 U152 ( .A(n776), .Y(n876) );
  OAI22X1 U153 ( .A0(n621), .A1(n769), .B0(n620), .B1(n813), .Y(n626) );
  AOI211X1 U154 ( .A0(n556), .A1(n821), .B0(n619), .C0(n618), .Y(n620) );
  AOI221X1 U155 ( .A0(n910), .A1(n535), .B0(n896), .B1(n556), .C0(n616), .Y(
        n621) );
  OAI22X1 U156 ( .A0(n859), .A1(n542), .B0(n550), .B1(n617), .Y(n619) );
  AOI222X1 U157 ( .A0(n867), .A1(n540), .B0(n863), .B1(n552), .C0(n547), .C1(
        n852), .Y(n567) );
  AOI21X1 U158 ( .A0(n873), .A1(n556), .B0(n557), .Y(n558) );
  OAI221XL U159 ( .A0(n551), .A1(n836), .B0(n543), .B1(n819), .C0(n677), .Y(
        n688) );
  AOI2BB2X1 U160 ( .B0(n910), .B1(n535), .A0N(n536), .A1N(n676), .Y(n677) );
  CLKINVX8 U161 ( .A(n546), .Y(n545) );
  CLKINVX3 U162 ( .A(n541), .Y(n539) );
  NOR2X1 U163 ( .A(n545), .B(n535), .Y(n721) );
  AOI211X1 U164 ( .A0(n878), .A1(n540), .B0(n719), .C0(n718), .Y(n731) );
  INVX1 U165 ( .A(n714), .Y(n878) );
  NAND2BX1 U166 ( .AN(n826), .B(n717), .Y(n718) );
  AOI222X1 U167 ( .A0(n916), .A1(n810), .B0(n724), .B1(n873), .C0(n886), .C1(
        n540), .Y(n725) );
  AOI221X1 U168 ( .A0(n602), .A1(n554), .B0(n540), .B1(n612), .C0(n596), .Y(
        n608) );
  OAI221XL U169 ( .A0(n536), .A1(n714), .B0(n545), .B1(n820), .C0(n635), .Y(
        n596) );
  AOI221X1 U170 ( .A0(n916), .A1(n852), .B0(n554), .B1(n810), .C0(n737), .Y(
        n749) );
  OAI2BB1X1 U171 ( .A0N(n781), .A1N(n547), .B0(n736), .Y(n737) );
  OAI221XL U172 ( .A0(n615), .A1(n551), .B0(n545), .B1(n758), .C0(n761), .Y(
        n616) );
  NOR2X1 U173 ( .A(n854), .B(n855), .Y(n615) );
  OAI221XL U174 ( .A0(n869), .A1(n545), .B0(n890), .B1(n829), .C0(n691), .Y(
        n706) );
  INVX1 U175 ( .A(n689), .Y(n869) );
  AOI32X1 U176 ( .A0(n889), .A1(n742), .A2(n556), .B0(n554), .B1(n690), .Y(
        n691) );
  OAI221XL U177 ( .A0(n856), .A1(n551), .B0(n541), .B1(n538), .C0(n629), .Y(
        n641) );
  INVX1 U178 ( .A(n808), .Y(n856) );
  AOI211X1 U179 ( .A0(n875), .A1(n556), .B0(n914), .C0(n628), .Y(n629) );
  INVX1 U180 ( .A(n809), .Y(n914) );
  AOI211X1 U181 ( .A0(n863), .A1(n540), .B0(n909), .C0(n559), .Y(n560) );
  NOR3X1 U182 ( .A(n545), .B(n884), .C(n862), .Y(n559) );
  INVX1 U183 ( .A(n664), .Y(n909) );
  OAI221XL U184 ( .A0(n536), .A1(n755), .B0(n759), .B1(n551), .C0(n754), .Y(
        n773) );
  AOI22X1 U185 ( .A0(n549), .A1(n889), .B0(n875), .B1(n539), .Y(n754) );
  AOI211X1 U186 ( .A0(n554), .A1(n827), .B0(n908), .C0(n826), .Y(n828) );
  CLKINVX3 U187 ( .A(n555), .Y(n551) );
  INVX1 U188 ( .A(n544), .Y(n542) );
  INVX1 U189 ( .A(n798), .Y(n913) );
  AOI221X1 U190 ( .A0(n797), .A1(n553), .B0(n796), .B1(n549), .C0(n795), .Y(
        n798) );
  OAI21XL U191 ( .A0(n536), .A1(n794), .B0(n793), .Y(n795) );
  INVX1 U192 ( .A(n536), .Y(n906) );
  NOR2X1 U193 ( .A(n884), .B(n866), .Y(n744) );
  CLKINVX3 U194 ( .A(n813), .Y(n900) );
  NAND3X1 U195 ( .A(n538), .B(n810), .C(n540), .Y(n834) );
  NAND2X1 U196 ( .A(n807), .B(n781), .Y(n838) );
  NAND2X1 U197 ( .A(n808), .B(n655), .Y(n765) );
  NAND2X1 U198 ( .A(n538), .B(n757), .Y(n612) );
  NOR2BX1 U199 ( .AN(n694), .B(n855), .Y(n759) );
  AOI21X1 U200 ( .A0(n742), .A1(n741), .B0(n536), .Y(n743) );
  OAI221XL U201 ( .A0(n887), .A1(n550), .B0(n802), .B1(n541), .C0(n783), .Y(
        n788) );
  INVX1 U202 ( .A(n838), .Y(n887) );
  AOI22X1 U203 ( .A0(n874), .A1(n548), .B0(n556), .B1(n782), .Y(n783) );
  AOI22X1 U204 ( .A0(n866), .A1(n546), .B0(n552), .B1(n810), .Y(n684) );
  AOI22X1 U205 ( .A0(n547), .A1(n612), .B0(n873), .B1(n539), .Y(n573) );
  NOR2X1 U206 ( .A(n785), .B(n536), .Y(n826) );
  NAND2X1 U207 ( .A(n680), .B(n781), .Y(n796) );
  INVX1 U208 ( .A(n769), .Y(n898) );
  NAND2X1 U209 ( .A(n694), .B(n680), .Y(n689) );
  CLKINVX3 U210 ( .A(n785), .Y(n867) );
  NAND2X1 U211 ( .A(n694), .B(n714), .Y(n663) );
  NOR2X1 U212 ( .A(n859), .B(n799), .Y(n802) );
  AOI211X1 U213 ( .A0(n556), .A1(n617), .B0(n588), .C0(n587), .Y(n594) );
  OAI2BB2X1 U214 ( .B0(n545), .B1(n740), .A0N(n735), .A1N(n540), .Y(n588) );
  AOI21X1 U215 ( .A0(n622), .A1(n586), .B0(n550), .Y(n587) );
  NAND2X1 U216 ( .A(n785), .B(n821), .Y(n696) );
  NAND2X1 U217 ( .A(n820), .B(n758), .Y(n735) );
  AOI21X1 U218 ( .A0(n556), .A1(n823), .B0(n822), .Y(n824) );
  AOI21X1 U219 ( .A0(n821), .A1(n820), .B0(n550), .Y(n822) );
  INVX1 U220 ( .A(n586), .Y(n858) );
  AOI22X1 U221 ( .A0(n899), .A1(n780), .B0(n901), .B1(n779), .Y(n790) );
  OAI221XL U222 ( .A0(n858), .A1(n551), .B0(n892), .B1(n536), .C0(n774), .Y(
        n780) );
  OAI221XL U223 ( .A0(n778), .A1(n545), .B0(n895), .B1(n551), .C0(n777), .Y(
        n779) );
  AOI2BB2X1 U224 ( .B0(n539), .B1(n836), .A0N(n545), .A1N(n802), .Y(n774) );
  INVX1 U225 ( .A(n715), .Y(n894) );
  INVX1 U226 ( .A(n624), .Y(n910) );
  INVX1 U227 ( .A(n823), .Y(n890) );
  AOI221XL U228 ( .A0(n556), .A1(n871), .B0(n548), .B1(n800), .C0(n599), .Y(
        n607) );
  INVX1 U229 ( .A(n597), .Y(n871) );
  OAI32X1 U230 ( .A0(n829), .A1(n860), .A2(n598), .B0(n886), .B1(n551), .Y(
        n599) );
  INVX1 U231 ( .A(n727), .Y(n892) );
  OAI221XL U232 ( .A0(n867), .A1(n545), .B0(n891), .B1(n829), .C0(n760), .Y(
        n772) );
  INVX1 U233 ( .A(n756), .Y(n891) );
  AOI22X1 U234 ( .A0(n759), .A1(n556), .B0(n794), .B1(n553), .Y(n760) );
  INVX1 U235 ( .A(n782), .Y(n896) );
  INVX1 U236 ( .A(n775), .Y(n895) );
  OAI221XL U237 ( .A0(n883), .A1(n551), .B0(n865), .B1(n545), .C0(n786), .Y(
        n787) );
  INVX1 U238 ( .A(n827), .Y(n883) );
  AOI31X1 U239 ( .A0(n821), .A1(n785), .A2(n556), .B0(n912), .Y(n786) );
  INVX1 U240 ( .A(n834), .Y(n912) );
  INVX1 U241 ( .A(n738), .Y(n904) );
  INVX1 U242 ( .A(n540), .Y(n543) );
  AOI211X1 U243 ( .A0(n901), .A1(n688), .B0(n687), .C0(n686), .Y(n708) );
  AOI211X1 U244 ( .A0(n900), .A1(n706), .B0(n705), .C0(n704), .Y(n707) );
  AOI31X1 U245 ( .A0(n685), .A1(n793), .A2(n684), .B0(n767), .Y(n686) );
  OAI2BB1X1 U246 ( .A0N(n790), .A1N(n789), .B0(n534), .Y(n791) );
  AOI22X1 U247 ( .A0(n900), .A1(n788), .B0(n898), .B1(n787), .Y(n789) );
  AOI22X1 U248 ( .A0(n752), .A1(n902), .B0(n534), .B1(n751), .Y(n753) );
  OAI221XL U249 ( .A0(n750), .A1(n815), .B0(n749), .B1(n769), .C0(n748), .Y(
        n751) );
  OAI221XL U250 ( .A0(n732), .A1(n769), .B0(n731), .B1(n767), .C0(n730), .Y(
        n752) );
  AOI22X1 U251 ( .A0(n533), .A1(n669), .B0(n668), .B1(n897), .Y(n670) );
  OAI221XL U252 ( .A0(n862), .A1(n551), .B0(n545), .B1(n663), .C0(n662), .Y(
        n669) );
  OAI221XL U253 ( .A0(n882), .A1(n545), .B0(n829), .B1(n742), .C0(n667), .Y(
        n668) );
  AOI21X1 U254 ( .A0(n890), .A1(n906), .B0(n661), .Y(n662) );
  AOI22X1 U255 ( .A0(n575), .A1(n897), .B0(n533), .B1(n574), .Y(n581) );
  OAI221XL U256 ( .A0(n536), .A1(n757), .B0(n637), .B1(n545), .C0(n572), .Y(
        n575) );
  OAI211X1 U257 ( .A0(n835), .A1(n550), .B0(n736), .C0(n573), .Y(n574) );
  AOI2BB2X1 U258 ( .B0(n539), .B1(n727), .A0N(n550), .A1N(n744), .Y(n572) );
  OAI22X1 U259 ( .A0(n634), .A1(n813), .B0(n633), .B1(n767), .Y(n640) );
  AOI221XL U260 ( .A0(n549), .A1(n740), .B0(n799), .B1(n850), .C0(n632), .Y(
        n633) );
  AOI221XL U261 ( .A0(n867), .A1(n916), .B0(n547), .B1(n713), .C0(n630), .Y(
        n634) );
  OAI32X1 U262 ( .A0(n738), .A1(n860), .A2(n850), .B0(n631), .B1(n904), .Y(
        n632) );
  OAI22X1 U263 ( .A0(n770), .A1(n769), .B0(n768), .B1(n767), .Y(n771) );
  AOI211X1 U264 ( .A0(n881), .A1(n850), .B0(n766), .C0(n907), .Y(n768) );
  AOI221XL U265 ( .A0(n862), .A1(n552), .B0(n547), .B1(n776), .C0(n764), .Y(
        n770) );
  OAI22X1 U266 ( .A0(n543), .A1(n852), .B0(n886), .B1(n550), .Y(n766) );
  OAI22X1 U267 ( .A0(n816), .A1(n815), .B0(n814), .B1(n813), .Y(n817) );
  AOI221XL U268 ( .A0(n549), .A1(n812), .B0(n876), .B1(n540), .C0(n811), .Y(
        n814) );
  AOI221X1 U269 ( .A0(n556), .A1(n808), .B0(n553), .B1(n807), .C0(n806), .Y(
        n816) );
  OAI221XL U270 ( .A0(n536), .A1(n810), .B0(n879), .B1(n551), .C0(n809), .Y(
        n811) );
  AOI211X1 U271 ( .A0(n868), .A1(n556), .B0(n652), .C0(n651), .Y(n653) );
  AOI31X1 U272 ( .A0(n809), .A1(n717), .A2(n650), .B0(n533), .Y(n651) );
  OAI22X1 U273 ( .A0(n857), .A1(n803), .B0(n649), .B1(n897), .Y(n652) );
  AOI2BB2X1 U274 ( .B0(n853), .B1(n552), .A0N(n833), .A1N(n545), .Y(n650) );
  AOI22X1 U275 ( .A0(n534), .A1(n610), .B0(n609), .B1(n902), .Y(n611) );
  OAI221XL U276 ( .A0(n595), .A1(n767), .B0(n594), .B1(n769), .C0(n593), .Y(
        n610) );
  OAI221XL U277 ( .A0(n608), .A1(n767), .B0(n607), .B1(n769), .C0(n606), .Y(
        n609) );
  AOI2BB2X1 U278 ( .B0(n659), .B1(n897), .A0N(n897), .A1N(n658), .Y(n671) );
  OAI221XL U279 ( .A0(n877), .A1(n551), .B0(n545), .B1(n807), .C0(n656), .Y(
        n659) );
  AOI221XL U281 ( .A0(n548), .A1(n676), .B0(n711), .B1(n540), .C0(n657), .Y(
        n658) );
  AOI22X1 U282 ( .A0(n539), .A1(n765), .B0(n873), .B1(n903), .Y(n656) );
  AOI22X1 U283 ( .A0(n553), .A1(n532), .B0(n539), .B1(n857), .Y(n631) );
  AOI22X1 U284 ( .A0(n900), .A1(n747), .B0(n899), .B1(n746), .Y(n748) );
  OAI221XL U285 ( .A0(n860), .A1(n545), .B0(n541), .B1(n807), .C0(n745), .Y(
        n746) );
  OAI221XL U286 ( .A0(n885), .A1(n536), .B0(n545), .B1(n740), .C0(n739), .Y(
        n747) );
  AOI21X1 U287 ( .A0(n744), .A1(n552), .B0(n743), .Y(n745) );
  AOI22X1 U288 ( .A0(n533), .A1(n562), .B0(n561), .B1(n897), .Y(n571) );
  OAI221XL U289 ( .A0(n880), .A1(n545), .B0(n541), .B1(n889), .C0(n558), .Y(
        n562) );
  OAI221XL U290 ( .A0(n532), .A1(n803), .B0(n722), .B1(n551), .C0(n560), .Y(
        n561) );
  INVX1 U291 ( .A(n663), .Y(n880) );
  AOI22X1 U292 ( .A0(n901), .A1(n605), .B0(n900), .B1(n604), .Y(n606) );
  OAI21XL U293 ( .A0(n602), .A1(n536), .B0(n601), .Y(n605) );
  OAI221XL U294 ( .A0(n551), .A1(n810), .B0(n835), .B1(n545), .C0(n603), .Y(
        n604) );
  AOI31X1 U295 ( .A0(n538), .A1(n742), .A2(n600), .B0(n910), .Y(n601) );
  CLKINVX3 U296 ( .A(n532), .Y(n852) );
  OAI21XL U297 ( .A0(n545), .A1(n537), .B0(n803), .Y(n647) );
  NAND2X1 U298 ( .A(n860), .B(n531), .Y(n755) );
  AOI21X1 U299 ( .A0(n699), .A1(n680), .B0(n545), .Y(n628) );
  INVX1 U300 ( .A(n531), .Y(n849) );
  OAI21XL U301 ( .A0(n850), .A1(n622), .B0(n550), .Y(n600) );
  OAI21XL U302 ( .A0(n850), .A1(n680), .B0(n550), .Y(n678) );
  OAI21XL U303 ( .A0(n536), .A1(n805), .B0(n763), .Y(n764) );
  AOI31X1 U304 ( .A0(n812), .A1(n903), .A2(n762), .B0(n915), .Y(n763) );
  INVX1 U305 ( .A(n761), .Y(n915) );
  OAI2BB1X1 U306 ( .A0N(n845), .A1N(n844), .B0(n902), .Y(n846) );
  AOI22X1 U307 ( .A0(n901), .A1(n843), .B0(n898), .B1(n842), .Y(n844) );
  AOI211X1 U308 ( .A0(n884), .A1(n540), .B0(n648), .C0(n647), .Y(n649) );
  OAI222X1 U309 ( .A0(n551), .A1(n807), .B0(n850), .B1(n693), .C0(n545), .C1(
        n821), .Y(n648) );
  AOI211X1 U310 ( .A0(n901), .A1(n627), .B0(n626), .C0(n625), .Y(n643) );
  AOI211X1 U311 ( .A0(n901), .A1(n641), .B0(n640), .C0(n911), .Y(n642) );
  OAI2BB2X1 U312 ( .B0(n614), .B1(n613), .A0N(n744), .A1N(n614), .Y(n627) );
  NAND2X1 U313 ( .A(n861), .B(n552), .Y(n636) );
  NOR2BX1 U314 ( .AN(n660), .B(n876), .Y(n722) );
  BUFX3 U315 ( .A(n841), .Y(n536) );
  NAND2X1 U316 ( .A(n850), .B(n903), .Y(n841) );
  OAI221XL U317 ( .A0(n531), .A1(n664), .B0(n543), .B1(n709), .C0(n636), .Y(
        n630) );
  BUFX3 U318 ( .A(n784), .Y(n538) );
  NAND2X1 U319 ( .A(n531), .B(n537), .Y(n784) );
  AOI211X1 U320 ( .A0(n540), .A1(n852), .B0(n585), .C0(n647), .Y(n595) );
  OAI222X1 U321 ( .A0(n551), .A1(n756), .B0(n584), .B1(n536), .C0(n545), .C1(
        n889), .Y(n585) );
  AOI21X1 U322 ( .A0(n537), .A1(n535), .B0(n858), .Y(n584) );
  AOI211X1 U323 ( .A0(n533), .A1(n569), .B0(n848), .C0(n568), .Y(n570) );
  OAI221XL U324 ( .A0(n545), .A1(n807), .B0(n602), .B1(n543), .C0(n564), .Y(
        n569) );
  AOI21X1 U325 ( .A0(n567), .A1(n566), .B0(n533), .Y(n568) );
  AOI31X1 U326 ( .A0(n556), .A1(n565), .A2(n884), .B0(n563), .Y(n564) );
  INVX1 U327 ( .A(n830), .Y(n546) );
  INVX1 U328 ( .A(n840), .Y(n555) );
  INVX1 U329 ( .A(n544), .Y(n541) );
  INVX1 U330 ( .A(n829), .Y(n544) );
  AOI22X1 U331 ( .A0(n533), .A1(n646), .B0(n645), .B1(n897), .Y(n654) );
  OAI222X1 U332 ( .A0(n545), .A1(n782), .B0(n551), .B1(n660), .C0(n894), .C1(
        n543), .Y(n646) );
  OAI221XL U333 ( .A0(n892), .A1(n536), .B0(n551), .B1(n819), .C0(n644), .Y(
        n645) );
  AOI2BB2X1 U334 ( .B0(n835), .B1(n539), .A0N(n545), .A1N(n726), .Y(n644) );
  NAND2X1 U335 ( .A(n699), .B(n622), .Y(n775) );
  NOR2BX1 U336 ( .AN(n660), .B(n862), .Y(n602) );
  AOI21X1 U337 ( .A0(n690), .A1(n758), .B0(n903), .Y(n661) );
  AOI22X1 U338 ( .A0(n556), .A1(n857), .B0(n539), .B1(n776), .Y(n777) );
  AOI22X1 U339 ( .A0(n549), .A1(n838), .B0(n882), .B1(n539), .Y(n839) );
  NAND2X1 U340 ( .A(n699), .B(n805), .Y(n715) );
  NAND2X1 U341 ( .A(n660), .B(n586), .Y(n756) );
  AOI21X1 U342 ( .A0(n660), .A1(n741), .B0(n545), .Y(n618) );
  AOI21X1 U343 ( .A0(n812), .A1(n538), .B0(n543), .Y(n720) );
  NAND2X1 U344 ( .A(n906), .B(n531), .Y(n717) );
  XNOR2X1 U345 ( .A(n903), .B(n531), .Y(n738) );
  NAND2X1 U346 ( .A(n539), .B(n537), .Y(n793) );
  XNOR2X1 U347 ( .A(n850), .B(n531), .Y(n762) );
  AOI21X1 U348 ( .A0(n833), .A1(n850), .B0(n556), .Y(n837) );
  AOI221X1 U349 ( .A0(n877), .A1(n540), .B0(n555), .B1(n735), .C0(n734), .Y(
        n750) );
  AOI21X1 U350 ( .A0(n536), .A1(n733), .B0(n799), .Y(n734) );
  OAI21XL U351 ( .A0(n861), .A1(n853), .B0(n850), .Y(n733) );
  AOI222X1 U352 ( .A0(n549), .A1(n713), .B0(n712), .B1(n711), .C0(n556), .C1(
        n537), .Y(n732) );
  OAI21XL U353 ( .A0(n850), .A1(n709), .B0(n550), .Y(n712) );
  AOI31X1 U354 ( .A0(n761), .A1(n624), .A2(n623), .B0(n767), .Y(n625) );
  AOI22X1 U355 ( .A0(n775), .A1(n850), .B0(n894), .B1(n554), .Y(n623) );
  AOI31X1 U356 ( .A0(n703), .A1(n793), .A2(n702), .B0(n815), .Y(n704) );
  OAI2BB1X1 U357 ( .A0N(n700), .A1N(n699), .B0(n554), .Y(n703) );
  AOI22X1 U358 ( .A0(n894), .A1(n556), .B0(n701), .B1(n547), .Y(n702) );
  INVX1 U359 ( .A(n830), .Y(n547) );
  INVX1 U360 ( .A(n830), .Y(n549) );
  INVX1 U361 ( .A(n830), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n565) );
  INVX1 U363 ( .A(n840), .Y(n553) );
  INVX1 U364 ( .A(n840), .Y(n554) );
  INVX1 U365 ( .A(n840), .Y(n552) );
  NOR2BX1 U366 ( .AN(n830), .B(n553), .Y(n614) );
  AOI22X1 U367 ( .A0(n581), .A1(a[0]), .B0(n580), .B1(n579), .Y(n582) );
  AOI31X1 U368 ( .A0(n717), .A1(n848), .A2(n571), .B0(n570), .Y(n583) );
  AOI22X1 U369 ( .A0(n576), .A1(n897), .B0(n556), .B1(n833), .Y(n580) );
  AOI22X1 U370 ( .A0(n673), .A1(n902), .B0(n534), .B1(n672), .Y(n674) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n654), .B0(n653), .B1(n848), .Y(n673) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n671), .B0(n670), .B1(n848), .Y(n672) );
  OAI22X1 U373 ( .A0(n698), .A1(n767), .B0(n697), .B1(n769), .Y(n705) );
  AOI221X1 U374 ( .A0(n548), .A1(n693), .B0(n556), .B1(n797), .C0(n692), .Y(
        n698) );
  AOI222X1 U375 ( .A0(n759), .A1(n547), .B0(a[2]), .B1(n696), .C0(n556), .C1(
        n695), .Y(n697) );
  OAI22X1 U376 ( .A0(n888), .A1(n542), .B0(n550), .B1(n537), .Y(n692) );
  NOR2X1 U377 ( .A(n863), .B(n861), .Y(n804) );
  BUFX3 U378 ( .A(n710), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n852), .Y(n710) );
  AOI221X1 U380 ( .A0(n916), .A1(n785), .B0(n851), .B1(n666), .C0(n665), .Y(
        n667) );
  NOR3X1 U381 ( .A(n851), .B(a[7]), .C(n860), .Y(n665) );
  INVX1 U382 ( .A(n762), .Y(n851) );
  OAI21XL U383 ( .A0(n857), .A1(n550), .B0(n664), .Y(n666) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI33X1 U385 ( .A0(n532), .A1(n540), .A2(n904), .B0(n738), .B1(n742), .B2(
        a[2]), .Y(n739) );
  AOI22X1 U386 ( .A0(n882), .A1(n850), .B0(a[2]), .B1(n612), .Y(n613) );
  CLKINVX3 U387 ( .A(a[0]), .Y(n848) );
  AOI211X1 U388 ( .A0(n724), .A1(n578), .B0(n577), .C0(a[0]), .Y(n579) );
  NAND2X1 U389 ( .A(n781), .B(n805), .Y(n578) );
  AOI21X1 U390 ( .A0(n803), .A1(n624), .B0(n897), .Y(n577) );
  BUFX3 U391 ( .A(a[5]), .Y(n533) );
  OAI221XL U392 ( .A0(n536), .A1(n808), .B0(n802), .B1(n545), .C0(n801), .Y(
        n818) );
  AOI22X1 U393 ( .A0(n539), .A1(n800), .B0(n799), .B1(a[2]), .Y(n801) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_7 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916;

  OAI221X4 U4 ( .A0(n857), .A1(n536), .B0(n862), .B1(n551), .C0(n839), .Y(n842) );
  OAI221X4 U6 ( .A0(n837), .A1(n836), .B0(n835), .B1(n551), .C0(n834), .Y(n843) );
  OAI222X4 U75 ( .A0(n551), .A1(n716), .B0(n742), .B1(n803), .C0(n545), .C1(
        n715), .Y(n719) );
  OAI32X4 U280 ( .A0(n551), .A1(n867), .A2(n870), .B0(n829), .B1(n820), .Y(
        n557) );
  AOI221X1 U1 ( .A0(n858), .A1(a[2]), .B0(n826), .B1(n565), .C0(n916), .Y(n566) );
  INVX1 U2 ( .A(a[7]), .Y(n903) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n820) );
  OAI222X1 U5 ( .A0(n829), .A1(n805), .B0(n804), .B1(n545), .C0(a[4]), .C1(
        n803), .Y(n806) );
  NAND2X2 U7 ( .A(n531), .B(n532), .Y(n808) );
  NAND2X1 U8 ( .A(n867), .B(n531), .Y(n694) );
  NAND2X2 U9 ( .A(n532), .B(n857), .Y(n742) );
  NAND2X1 U10 ( .A(n884), .B(n531), .Y(n781) );
  NAND2X2 U11 ( .A(n537), .B(n742), .Y(n810) );
  NAND2X2 U12 ( .A(n857), .B(n535), .Y(n807) );
  CLKINVX3 U13 ( .A(n533), .Y(n897) );
  NAND2X2 U14 ( .A(n857), .B(n852), .Y(n785) );
  NAND2X1 U15 ( .A(n531), .B(n742), .Y(n821) );
  CLKINVX3 U16 ( .A(a[2]), .Y(n850) );
  NAND2X1 U17 ( .A(n533), .B(n848), .Y(n813) );
  NAND2X2 U18 ( .A(n848), .B(n897), .Y(n769) );
  NAND2X2 U19 ( .A(a[0]), .B(n897), .Y(n767) );
  CLKINVX3 U20 ( .A(n534), .Y(n902) );
  OAI22X2 U21 ( .A0(n583), .A1(n902), .B0(n534), .B1(n582), .Y(d[0]) );
  OAI22X2 U22 ( .A0(n534), .A1(n643), .B0(n642), .B1(n902), .Y(d[2]) );
  OAI21X2 U23 ( .A0(n847), .A1(n902), .B0(n846), .Y(d[7]) );
  AOI221X1 U24 ( .A0(n899), .A1(n913), .B0(n898), .B1(n818), .C0(n817), .Y(
        n847) );
  OAI22X2 U25 ( .A0(n534), .A1(n708), .B0(n707), .B1(n902), .Y(d[4]) );
  OAI21X2 U26 ( .A0(n534), .A1(n792), .B0(n791), .Y(d[6]) );
  AOI221X1 U27 ( .A0(n900), .A1(n773), .B0(n901), .B1(n772), .C0(n771), .Y(
        n792) );
  NAND2X1 U28 ( .A(a[2]), .B(n903), .Y(n840) );
  NAND2X1 U29 ( .A(a[7]), .B(n850), .Y(n830) );
  AOI21XL U30 ( .A0(n916), .A1(a[4]), .B0(n907), .Y(n603) );
  NAND2X1 U31 ( .A(a[4]), .B(n535), .Y(n660) );
  NAND2X1 U32 ( .A(n531), .B(a[4]), .Y(n699) );
  NAND2X2 U33 ( .A(n532), .B(a[4]), .Y(n812) );
  CLKINVX3 U34 ( .A(a[4]), .Y(n857) );
  CLKINVX3 U35 ( .A(n542), .Y(n540) );
  NAND2X1 U36 ( .A(n870), .B(n906), .Y(n635) );
  INVX1 U37 ( .A(n598), .Y(n889) );
  NAND2X1 U38 ( .A(n810), .B(n535), .Y(n709) );
  CLKINVX3 U39 ( .A(n555), .Y(n550) );
  NAND2X1 U40 ( .A(n867), .B(n535), .Y(n690) );
  NAND2X1 U41 ( .A(n873), .B(n535), .Y(n622) );
  NAND2X1 U42 ( .A(n538), .B(n655), .Y(n711) );
  NAND2X1 U43 ( .A(n808), .B(n714), .Y(n713) );
  NAND2X1 U44 ( .A(n776), .B(n709), .Y(n716) );
  INVX1 U45 ( .A(n755), .Y(n861) );
  INVX1 U46 ( .A(n538), .Y(n870) );
  INVX1 U47 ( .A(n741), .Y(n866) );
  NOR2X1 U48 ( .A(n535), .B(n884), .Y(n598) );
  NAND2X1 U49 ( .A(n535), .B(n852), .Y(n805) );
  NAND2X1 U50 ( .A(n785), .B(n535), .Y(n700) );
  NAND2X1 U51 ( .A(n884), .B(n535), .Y(n675) );
  NAND2X1 U52 ( .A(n742), .B(n535), .Y(n757) );
  NAND2X1 U53 ( .A(n694), .B(n675), .Y(n836) );
  INVX1 U54 ( .A(n821), .Y(n862) );
  NAND2X1 U55 ( .A(n808), .B(n700), .Y(n617) );
  INVX1 U56 ( .A(n693), .Y(n854) );
  INVX1 U57 ( .A(n807), .Y(n859) );
  INVX1 U58 ( .A(n820), .Y(n855) );
  BUFX3 U59 ( .A(n849), .Y(n535) );
  NAND2X1 U60 ( .A(n873), .B(n531), .Y(n776) );
  NAND2X1 U61 ( .A(n531), .B(n539), .Y(n803) );
  NAND2X1 U62 ( .A(n812), .B(n535), .Y(n655) );
  NAND2X1 U63 ( .A(n531), .B(n810), .Y(n758) );
  NAND2X1 U64 ( .A(n531), .B(n785), .Y(n741) );
  INVX1 U65 ( .A(n611), .Y(d[1]) );
  INVX1 U66 ( .A(n753), .Y(d[5]) );
  NAND2X1 U67 ( .A(n906), .B(n532), .Y(n664) );
  INVX1 U68 ( .A(n537), .Y(n877) );
  NAND2X1 U69 ( .A(n812), .B(n776), .Y(n827) );
  NOR2X1 U70 ( .A(n537), .B(n535), .Y(n799) );
  CLKINVX3 U71 ( .A(n812), .Y(n884) );
  NAND2X1 U72 ( .A(n531), .B(n852), .Y(n693) );
  NAND2X1 U73 ( .A(n531), .B(n857), .Y(n586) );
  NAND2BX1 U74 ( .AN(n799), .B(n660), .Y(n727) );
  INVX1 U76 ( .A(n767), .Y(n899) );
  NAND2X1 U77 ( .A(n699), .B(n655), .Y(n782) );
  NAND2BX1 U78 ( .AN(n830), .B(n537), .Y(n624) );
  NAND2X1 U79 ( .A(n699), .B(n690), .Y(n819) );
  NAND2X1 U80 ( .A(n660), .B(n781), .Y(n823) );
  CLKINVX3 U81 ( .A(n815), .Y(n901) );
  BUFX3 U82 ( .A(a[1]), .Y(n531) );
  NAND2X1 U83 ( .A(a[7]), .B(a[2]), .Y(n829) );
  INVX1 U84 ( .A(n674), .Y(d[3]) );
  NAND2X1 U85 ( .A(n533), .B(a[0]), .Y(n815) );
  INVX1 U86 ( .A(n685), .Y(n907) );
  NAND2X1 U87 ( .A(n864), .B(n540), .Y(n809) );
  NAND2X1 U88 ( .A(n872), .B(n556), .Y(n685) );
  INVX1 U89 ( .A(n635), .Y(n908) );
  NOR2X1 U90 ( .A(n550), .B(n598), .Y(n724) );
  NOR2X1 U91 ( .A(n874), .B(n861), .Y(n676) );
  NAND2X1 U92 ( .A(n701), .B(n540), .Y(n761) );
  INVX1 U93 ( .A(n622), .Y(n874) );
  INVX1 U94 ( .A(n675), .Y(n886) );
  INVX1 U95 ( .A(n757), .Y(n863) );
  INVX1 U96 ( .A(n716), .Y(n875) );
  INVX1 U97 ( .A(n695), .Y(n872) );
  INVX1 U98 ( .A(n713), .Y(n879) );
  INVX4 U99 ( .A(n536), .Y(n556) );
  NOR2BX1 U100 ( .AN(n709), .B(n854), .Y(n835) );
  NOR2X1 U101 ( .A(n870), .B(n853), .Y(n597) );
  NOR2X1 U102 ( .A(n873), .B(n862), .Y(n637) );
  NAND2X1 U103 ( .A(n889), .B(n700), .Y(n740) );
  INVX1 U104 ( .A(n805), .Y(n853) );
  NAND2X1 U105 ( .A(n889), .B(n675), .Y(n800) );
  INVX1 U106 ( .A(n690), .Y(n868) );
  INVX1 U107 ( .A(n700), .Y(n864) );
  NOR2X1 U108 ( .A(n866), .B(n868), .Y(n726) );
  OAI221XL U109 ( .A0(n865), .A1(n545), .B0(n825), .B1(n543), .C0(n905), .Y(
        n576) );
  INVX1 U110 ( .A(n724), .Y(n905) );
  INVX1 U111 ( .A(n796), .Y(n888) );
  NOR2X1 U112 ( .A(n864), .B(n854), .Y(n825) );
  INVX1 U113 ( .A(n711), .Y(n882) );
  NOR2X1 U114 ( .A(n861), .B(n868), .Y(n778) );
  INVX1 U115 ( .A(n617), .Y(n865) );
  INVX1 U116 ( .A(n765), .Y(n881) );
  INVX1 U117 ( .A(n836), .Y(n885) );
  NAND2X1 U118 ( .A(n860), .B(n535), .Y(n680) );
  NAND2X1 U119 ( .A(n877), .B(n535), .Y(n714) );
  OAI22X1 U120 ( .A0(n683), .A1(n813), .B0(n682), .B1(n769), .Y(n687) );
  AOI222X1 U121 ( .A0(n862), .A1(n548), .B0(n556), .B1(n679), .C0(n678), .C1(
        n711), .Y(n683) );
  AOI211X1 U122 ( .A0(n556), .A1(n689), .B0(n681), .C0(n724), .Y(n682) );
  NAND2X1 U123 ( .A(n807), .B(n694), .Y(n679) );
  NOR2X1 U124 ( .A(n877), .B(n866), .Y(n701) );
  OAI22X1 U125 ( .A0(n542), .A1(n716), .B0(n545), .B1(n538), .Y(n681) );
  CLKINVX3 U126 ( .A(n810), .Y(n873) );
  NAND2X1 U127 ( .A(n709), .B(n781), .Y(n833) );
  CLKINVX3 U128 ( .A(n742), .Y(n860) );
  AOI22X1 U129 ( .A0(n899), .A1(n832), .B0(n900), .B1(n831), .Y(n845) );
  OAI221XL U130 ( .A0(n825), .A1(n545), .B0(n893), .B1(n541), .C0(n824), .Y(
        n832) );
  OAI221XL U131 ( .A0(n881), .A1(n545), .B0(n872), .B1(n542), .C0(n828), .Y(
        n831) );
  INVX1 U132 ( .A(n819), .Y(n893) );
  NAND2X1 U133 ( .A(n556), .B(n827), .Y(n736) );
  NAND2X1 U134 ( .A(n808), .B(n709), .Y(n695) );
  AOI22X1 U135 ( .A0(n900), .A1(n729), .B0(n901), .B1(n728), .Y(n730) );
  OAI221XL U136 ( .A0(n877), .A1(n551), .B0(n860), .B1(n545), .C0(n723), .Y(
        n729) );
  OAI221XL U137 ( .A0(n536), .A1(n727), .B0(n726), .B1(n545), .C0(n725), .Y(
        n728) );
  AOI211X1 U138 ( .A0(n722), .A1(n556), .B0(n721), .C0(n720), .Y(n723) );
  AOI22X1 U139 ( .A0(n900), .A1(n592), .B0(n901), .B1(n591), .Y(n593) );
  OAI221XL U140 ( .A0(n888), .A1(n545), .B0(n879), .B1(n542), .C0(n590), .Y(
        n591) );
  OAI211X1 U141 ( .A0(n597), .A1(n550), .B0(n635), .C0(n589), .Y(n592) );
  AOI22X1 U142 ( .A0(n888), .A1(n906), .B0(n884), .B1(n553), .Y(n590) );
  AOI22X1 U143 ( .A0(n548), .A1(n860), .B0(n676), .B1(n539), .Y(n589) );
  AOI21X1 U144 ( .A0(n808), .A1(n680), .B0(n550), .Y(n563) );
  INVX1 U145 ( .A(n803), .Y(n916) );
  AND2X2 U146 ( .A(n758), .B(n757), .Y(n794) );
  NAND2X1 U147 ( .A(n538), .B(n709), .Y(n797) );
  OAI21XL U148 ( .A0(n758), .A1(n550), .B0(n736), .Y(n657) );
  INVX1 U149 ( .A(n639), .Y(n911) );
  OAI31X1 U150 ( .A0(n721), .A1(n908), .A2(n638), .B0(n898), .Y(n639) );
  OAI21XL U151 ( .A0(n541), .A1(n637), .B0(n636), .Y(n638) );
  INVX1 U152 ( .A(n776), .Y(n876) );
  OAI22X1 U153 ( .A0(n621), .A1(n769), .B0(n620), .B1(n813), .Y(n626) );
  AOI211X1 U154 ( .A0(n556), .A1(n821), .B0(n619), .C0(n618), .Y(n620) );
  AOI221X1 U155 ( .A0(n910), .A1(n535), .B0(n896), .B1(n556), .C0(n616), .Y(
        n621) );
  OAI22X1 U156 ( .A0(n859), .A1(n542), .B0(n550), .B1(n617), .Y(n619) );
  AOI222X1 U157 ( .A0(n867), .A1(n540), .B0(n863), .B1(n552), .C0(n547), .C1(
        n852), .Y(n567) );
  AOI21X1 U158 ( .A0(n873), .A1(n556), .B0(n557), .Y(n558) );
  OAI221XL U159 ( .A0(n551), .A1(n836), .B0(n543), .B1(n819), .C0(n677), .Y(
        n688) );
  AOI2BB2X1 U160 ( .B0(n910), .B1(n535), .A0N(n536), .A1N(n676), .Y(n677) );
  CLKINVX8 U161 ( .A(n546), .Y(n545) );
  CLKINVX3 U162 ( .A(n541), .Y(n539) );
  NOR2X1 U163 ( .A(n545), .B(n535), .Y(n721) );
  AOI211X1 U164 ( .A0(n878), .A1(n540), .B0(n719), .C0(n718), .Y(n731) );
  INVX1 U165 ( .A(n714), .Y(n878) );
  NAND2BX1 U166 ( .AN(n826), .B(n717), .Y(n718) );
  AOI222X1 U167 ( .A0(n916), .A1(n810), .B0(n724), .B1(n873), .C0(n886), .C1(
        n540), .Y(n725) );
  AOI221X1 U168 ( .A0(n602), .A1(n554), .B0(n540), .B1(n612), .C0(n596), .Y(
        n608) );
  OAI221XL U169 ( .A0(n536), .A1(n714), .B0(n545), .B1(n820), .C0(n635), .Y(
        n596) );
  AOI221X1 U170 ( .A0(n916), .A1(n852), .B0(n554), .B1(n810), .C0(n737), .Y(
        n749) );
  OAI2BB1X1 U171 ( .A0N(n781), .A1N(n547), .B0(n736), .Y(n737) );
  OAI221XL U172 ( .A0(n615), .A1(n551), .B0(n545), .B1(n758), .C0(n761), .Y(
        n616) );
  NOR2X1 U173 ( .A(n854), .B(n855), .Y(n615) );
  OAI221XL U174 ( .A0(n869), .A1(n545), .B0(n890), .B1(n829), .C0(n691), .Y(
        n706) );
  INVX1 U175 ( .A(n689), .Y(n869) );
  AOI32X1 U176 ( .A0(n889), .A1(n742), .A2(n556), .B0(n554), .B1(n690), .Y(
        n691) );
  OAI221XL U177 ( .A0(n856), .A1(n551), .B0(n541), .B1(n538), .C0(n629), .Y(
        n641) );
  INVX1 U178 ( .A(n808), .Y(n856) );
  AOI211X1 U179 ( .A0(n875), .A1(n556), .B0(n914), .C0(n628), .Y(n629) );
  INVX1 U180 ( .A(n809), .Y(n914) );
  AOI211X1 U181 ( .A0(n863), .A1(n540), .B0(n909), .C0(n559), .Y(n560) );
  NOR3X1 U182 ( .A(n545), .B(n884), .C(n862), .Y(n559) );
  INVX1 U183 ( .A(n664), .Y(n909) );
  OAI221XL U184 ( .A0(n536), .A1(n755), .B0(n759), .B1(n551), .C0(n754), .Y(
        n773) );
  AOI22X1 U185 ( .A0(n549), .A1(n889), .B0(n875), .B1(n539), .Y(n754) );
  AOI211X1 U186 ( .A0(n554), .A1(n827), .B0(n908), .C0(n826), .Y(n828) );
  CLKINVX3 U187 ( .A(n555), .Y(n551) );
  INVX1 U188 ( .A(n544), .Y(n542) );
  INVX1 U189 ( .A(n798), .Y(n913) );
  AOI221X1 U190 ( .A0(n797), .A1(n553), .B0(n796), .B1(n549), .C0(n795), .Y(
        n798) );
  OAI21XL U191 ( .A0(n536), .A1(n794), .B0(n793), .Y(n795) );
  INVX1 U192 ( .A(n536), .Y(n906) );
  NOR2X1 U193 ( .A(n884), .B(n866), .Y(n744) );
  CLKINVX3 U194 ( .A(n813), .Y(n900) );
  NAND3X1 U195 ( .A(n538), .B(n810), .C(n540), .Y(n834) );
  NAND2X1 U196 ( .A(n807), .B(n781), .Y(n838) );
  NAND2X1 U197 ( .A(n808), .B(n655), .Y(n765) );
  NAND2X1 U198 ( .A(n538), .B(n757), .Y(n612) );
  NOR2BX1 U199 ( .AN(n694), .B(n855), .Y(n759) );
  AOI21X1 U200 ( .A0(n742), .A1(n741), .B0(n536), .Y(n743) );
  OAI221XL U201 ( .A0(n887), .A1(n550), .B0(n802), .B1(n541), .C0(n783), .Y(
        n788) );
  INVX1 U202 ( .A(n838), .Y(n887) );
  AOI22X1 U203 ( .A0(n874), .A1(n548), .B0(n556), .B1(n782), .Y(n783) );
  AOI22X1 U204 ( .A0(n866), .A1(n546), .B0(n552), .B1(n810), .Y(n684) );
  AOI22X1 U205 ( .A0(n547), .A1(n612), .B0(n873), .B1(n539), .Y(n573) );
  NOR2X1 U206 ( .A(n785), .B(n536), .Y(n826) );
  NAND2X1 U207 ( .A(n680), .B(n781), .Y(n796) );
  INVX1 U208 ( .A(n769), .Y(n898) );
  NAND2X1 U209 ( .A(n694), .B(n680), .Y(n689) );
  CLKINVX3 U210 ( .A(n785), .Y(n867) );
  NAND2X1 U211 ( .A(n694), .B(n714), .Y(n663) );
  NOR2X1 U212 ( .A(n859), .B(n799), .Y(n802) );
  AOI211X1 U213 ( .A0(n556), .A1(n617), .B0(n588), .C0(n587), .Y(n594) );
  OAI2BB2X1 U214 ( .B0(n545), .B1(n740), .A0N(n735), .A1N(n540), .Y(n588) );
  AOI21X1 U215 ( .A0(n622), .A1(n586), .B0(n550), .Y(n587) );
  NAND2X1 U216 ( .A(n785), .B(n821), .Y(n696) );
  NAND2X1 U217 ( .A(n820), .B(n758), .Y(n735) );
  AOI21X1 U218 ( .A0(n556), .A1(n823), .B0(n822), .Y(n824) );
  AOI21X1 U219 ( .A0(n821), .A1(n820), .B0(n550), .Y(n822) );
  INVX1 U220 ( .A(n586), .Y(n858) );
  AOI22X1 U221 ( .A0(n899), .A1(n780), .B0(n901), .B1(n779), .Y(n790) );
  OAI221XL U222 ( .A0(n858), .A1(n551), .B0(n892), .B1(n536), .C0(n774), .Y(
        n780) );
  OAI221XL U223 ( .A0(n778), .A1(n545), .B0(n895), .B1(n551), .C0(n777), .Y(
        n779) );
  AOI2BB2X1 U224 ( .B0(n539), .B1(n836), .A0N(n545), .A1N(n802), .Y(n774) );
  INVX1 U225 ( .A(n715), .Y(n894) );
  INVX1 U226 ( .A(n624), .Y(n910) );
  INVX1 U227 ( .A(n823), .Y(n890) );
  AOI221XL U228 ( .A0(n556), .A1(n871), .B0(n548), .B1(n800), .C0(n599), .Y(
        n607) );
  INVX1 U229 ( .A(n597), .Y(n871) );
  OAI32X1 U230 ( .A0(n829), .A1(n860), .A2(n598), .B0(n886), .B1(n551), .Y(
        n599) );
  INVX1 U231 ( .A(n727), .Y(n892) );
  OAI221XL U232 ( .A0(n867), .A1(n545), .B0(n891), .B1(n829), .C0(n760), .Y(
        n772) );
  INVX1 U233 ( .A(n756), .Y(n891) );
  AOI22X1 U234 ( .A0(n759), .A1(n556), .B0(n794), .B1(n553), .Y(n760) );
  INVX1 U235 ( .A(n782), .Y(n896) );
  INVX1 U236 ( .A(n775), .Y(n895) );
  OAI221XL U237 ( .A0(n883), .A1(n551), .B0(n865), .B1(n545), .C0(n786), .Y(
        n787) );
  INVX1 U238 ( .A(n827), .Y(n883) );
  AOI31X1 U239 ( .A0(n821), .A1(n785), .A2(n556), .B0(n912), .Y(n786) );
  INVX1 U240 ( .A(n834), .Y(n912) );
  INVX1 U241 ( .A(n738), .Y(n904) );
  INVX1 U242 ( .A(n540), .Y(n543) );
  AOI211X1 U243 ( .A0(n901), .A1(n688), .B0(n687), .C0(n686), .Y(n708) );
  AOI211X1 U244 ( .A0(n900), .A1(n706), .B0(n705), .C0(n704), .Y(n707) );
  AOI31X1 U245 ( .A0(n685), .A1(n793), .A2(n684), .B0(n767), .Y(n686) );
  OAI2BB1X1 U246 ( .A0N(n790), .A1N(n789), .B0(n534), .Y(n791) );
  AOI22X1 U247 ( .A0(n900), .A1(n788), .B0(n898), .B1(n787), .Y(n789) );
  AOI22X1 U248 ( .A0(n752), .A1(n902), .B0(n534), .B1(n751), .Y(n753) );
  OAI221XL U249 ( .A0(n750), .A1(n815), .B0(n749), .B1(n769), .C0(n748), .Y(
        n751) );
  OAI221XL U250 ( .A0(n732), .A1(n769), .B0(n731), .B1(n767), .C0(n730), .Y(
        n752) );
  AOI22X1 U251 ( .A0(n533), .A1(n669), .B0(n668), .B1(n897), .Y(n670) );
  OAI221XL U252 ( .A0(n862), .A1(n551), .B0(n545), .B1(n663), .C0(n662), .Y(
        n669) );
  OAI221XL U253 ( .A0(n882), .A1(n545), .B0(n829), .B1(n742), .C0(n667), .Y(
        n668) );
  AOI21X1 U254 ( .A0(n890), .A1(n906), .B0(n661), .Y(n662) );
  AOI22X1 U255 ( .A0(n575), .A1(n897), .B0(n533), .B1(n574), .Y(n581) );
  OAI221XL U256 ( .A0(n536), .A1(n757), .B0(n637), .B1(n545), .C0(n572), .Y(
        n575) );
  OAI211X1 U257 ( .A0(n835), .A1(n550), .B0(n736), .C0(n573), .Y(n574) );
  AOI2BB2X1 U258 ( .B0(n539), .B1(n727), .A0N(n550), .A1N(n744), .Y(n572) );
  OAI22X1 U259 ( .A0(n634), .A1(n813), .B0(n633), .B1(n767), .Y(n640) );
  AOI221XL U260 ( .A0(n549), .A1(n740), .B0(n799), .B1(n850), .C0(n632), .Y(
        n633) );
  AOI221XL U261 ( .A0(n867), .A1(n916), .B0(n547), .B1(n713), .C0(n630), .Y(
        n634) );
  OAI32X1 U262 ( .A0(n738), .A1(n860), .A2(n850), .B0(n631), .B1(n904), .Y(
        n632) );
  OAI22X1 U263 ( .A0(n770), .A1(n769), .B0(n768), .B1(n767), .Y(n771) );
  AOI211X1 U264 ( .A0(n881), .A1(n850), .B0(n766), .C0(n907), .Y(n768) );
  AOI221XL U265 ( .A0(n862), .A1(n552), .B0(n547), .B1(n776), .C0(n764), .Y(
        n770) );
  OAI22X1 U266 ( .A0(n543), .A1(n852), .B0(n886), .B1(n550), .Y(n766) );
  OAI22X1 U267 ( .A0(n816), .A1(n815), .B0(n814), .B1(n813), .Y(n817) );
  AOI221XL U268 ( .A0(n549), .A1(n812), .B0(n876), .B1(n540), .C0(n811), .Y(
        n814) );
  AOI221X1 U269 ( .A0(n556), .A1(n808), .B0(n553), .B1(n807), .C0(n806), .Y(
        n816) );
  OAI221XL U270 ( .A0(n536), .A1(n810), .B0(n879), .B1(n551), .C0(n809), .Y(
        n811) );
  AOI211X1 U271 ( .A0(n868), .A1(n556), .B0(n652), .C0(n651), .Y(n653) );
  AOI31X1 U272 ( .A0(n809), .A1(n717), .A2(n650), .B0(n533), .Y(n651) );
  OAI22X1 U273 ( .A0(n857), .A1(n803), .B0(n649), .B1(n897), .Y(n652) );
  AOI2BB2X1 U274 ( .B0(n853), .B1(n552), .A0N(n833), .A1N(n545), .Y(n650) );
  AOI22X1 U275 ( .A0(n534), .A1(n610), .B0(n609), .B1(n902), .Y(n611) );
  OAI221XL U276 ( .A0(n595), .A1(n767), .B0(n594), .B1(n769), .C0(n593), .Y(
        n610) );
  OAI221XL U277 ( .A0(n608), .A1(n767), .B0(n607), .B1(n769), .C0(n606), .Y(
        n609) );
  AOI2BB2X1 U278 ( .B0(n659), .B1(n897), .A0N(n897), .A1N(n658), .Y(n671) );
  OAI221XL U279 ( .A0(n877), .A1(n551), .B0(n545), .B1(n807), .C0(n656), .Y(
        n659) );
  AOI221XL U281 ( .A0(n548), .A1(n676), .B0(n711), .B1(n540), .C0(n657), .Y(
        n658) );
  AOI22X1 U282 ( .A0(n539), .A1(n765), .B0(n873), .B1(n903), .Y(n656) );
  AOI22X1 U283 ( .A0(n553), .A1(n532), .B0(n539), .B1(n857), .Y(n631) );
  AOI22X1 U284 ( .A0(n900), .A1(n747), .B0(n899), .B1(n746), .Y(n748) );
  OAI221XL U285 ( .A0(n860), .A1(n545), .B0(n541), .B1(n807), .C0(n745), .Y(
        n746) );
  OAI221XL U286 ( .A0(n885), .A1(n536), .B0(n545), .B1(n740), .C0(n739), .Y(
        n747) );
  AOI21X1 U287 ( .A0(n744), .A1(n552), .B0(n743), .Y(n745) );
  AOI22X1 U288 ( .A0(n533), .A1(n562), .B0(n561), .B1(n897), .Y(n571) );
  OAI221XL U289 ( .A0(n880), .A1(n545), .B0(n541), .B1(n889), .C0(n558), .Y(
        n562) );
  OAI221XL U290 ( .A0(n532), .A1(n803), .B0(n722), .B1(n551), .C0(n560), .Y(
        n561) );
  INVX1 U291 ( .A(n663), .Y(n880) );
  AOI22X1 U292 ( .A0(n901), .A1(n605), .B0(n900), .B1(n604), .Y(n606) );
  OAI21XL U293 ( .A0(n602), .A1(n536), .B0(n601), .Y(n605) );
  OAI221XL U294 ( .A0(n551), .A1(n810), .B0(n835), .B1(n545), .C0(n603), .Y(
        n604) );
  AOI31X1 U295 ( .A0(n538), .A1(n742), .A2(n600), .B0(n910), .Y(n601) );
  CLKINVX3 U296 ( .A(n532), .Y(n852) );
  OAI21XL U297 ( .A0(n545), .A1(n537), .B0(n803), .Y(n647) );
  NAND2X1 U298 ( .A(n860), .B(n531), .Y(n755) );
  AOI21X1 U299 ( .A0(n699), .A1(n680), .B0(n545), .Y(n628) );
  INVX1 U300 ( .A(n531), .Y(n849) );
  OAI21XL U301 ( .A0(n850), .A1(n622), .B0(n550), .Y(n600) );
  OAI21XL U302 ( .A0(n850), .A1(n680), .B0(n550), .Y(n678) );
  OAI21XL U303 ( .A0(n536), .A1(n805), .B0(n763), .Y(n764) );
  AOI31X1 U304 ( .A0(n812), .A1(n903), .A2(n762), .B0(n915), .Y(n763) );
  INVX1 U305 ( .A(n761), .Y(n915) );
  OAI2BB1X1 U306 ( .A0N(n845), .A1N(n844), .B0(n902), .Y(n846) );
  AOI22X1 U307 ( .A0(n901), .A1(n843), .B0(n898), .B1(n842), .Y(n844) );
  AOI211X1 U308 ( .A0(n884), .A1(n540), .B0(n648), .C0(n647), .Y(n649) );
  OAI222X1 U309 ( .A0(n551), .A1(n807), .B0(n850), .B1(n693), .C0(n545), .C1(
        n821), .Y(n648) );
  AOI211X1 U310 ( .A0(n901), .A1(n627), .B0(n626), .C0(n625), .Y(n643) );
  AOI211X1 U311 ( .A0(n901), .A1(n641), .B0(n640), .C0(n911), .Y(n642) );
  OAI2BB2X1 U312 ( .B0(n614), .B1(n613), .A0N(n744), .A1N(n614), .Y(n627) );
  NAND2X1 U313 ( .A(n861), .B(n552), .Y(n636) );
  NOR2BX1 U314 ( .AN(n660), .B(n876), .Y(n722) );
  BUFX3 U315 ( .A(n841), .Y(n536) );
  NAND2X1 U316 ( .A(n850), .B(n903), .Y(n841) );
  OAI221XL U317 ( .A0(n531), .A1(n664), .B0(n543), .B1(n709), .C0(n636), .Y(
        n630) );
  BUFX3 U318 ( .A(n784), .Y(n538) );
  NAND2X1 U319 ( .A(n531), .B(n537), .Y(n784) );
  AOI211X1 U320 ( .A0(n540), .A1(n852), .B0(n585), .C0(n647), .Y(n595) );
  OAI222X1 U321 ( .A0(n551), .A1(n756), .B0(n584), .B1(n536), .C0(n545), .C1(
        n889), .Y(n585) );
  AOI21X1 U322 ( .A0(n537), .A1(n535), .B0(n858), .Y(n584) );
  AOI211X1 U323 ( .A0(n533), .A1(n569), .B0(n848), .C0(n568), .Y(n570) );
  OAI221XL U324 ( .A0(n545), .A1(n807), .B0(n602), .B1(n543), .C0(n564), .Y(
        n569) );
  AOI21X1 U325 ( .A0(n567), .A1(n566), .B0(n533), .Y(n568) );
  AOI31X1 U326 ( .A0(n556), .A1(n565), .A2(n884), .B0(n563), .Y(n564) );
  INVX1 U327 ( .A(n830), .Y(n546) );
  INVX1 U328 ( .A(n840), .Y(n555) );
  INVX1 U329 ( .A(n544), .Y(n541) );
  INVX1 U330 ( .A(n829), .Y(n544) );
  AOI22X1 U331 ( .A0(n533), .A1(n646), .B0(n645), .B1(n897), .Y(n654) );
  OAI222X1 U332 ( .A0(n545), .A1(n782), .B0(n551), .B1(n660), .C0(n894), .C1(
        n543), .Y(n646) );
  OAI221XL U333 ( .A0(n892), .A1(n536), .B0(n551), .B1(n819), .C0(n644), .Y(
        n645) );
  AOI2BB2X1 U334 ( .B0(n835), .B1(n539), .A0N(n545), .A1N(n726), .Y(n644) );
  NAND2X1 U335 ( .A(n699), .B(n622), .Y(n775) );
  NOR2BX1 U336 ( .AN(n660), .B(n862), .Y(n602) );
  AOI21X1 U337 ( .A0(n690), .A1(n758), .B0(n903), .Y(n661) );
  AOI22X1 U338 ( .A0(n556), .A1(n857), .B0(n539), .B1(n776), .Y(n777) );
  AOI22X1 U339 ( .A0(n549), .A1(n838), .B0(n882), .B1(n539), .Y(n839) );
  NAND2X1 U340 ( .A(n699), .B(n805), .Y(n715) );
  NAND2X1 U341 ( .A(n660), .B(n586), .Y(n756) );
  AOI21X1 U342 ( .A0(n660), .A1(n741), .B0(n545), .Y(n618) );
  AOI21X1 U343 ( .A0(n812), .A1(n538), .B0(n543), .Y(n720) );
  NAND2X1 U344 ( .A(n906), .B(n531), .Y(n717) );
  XNOR2X1 U345 ( .A(n903), .B(n531), .Y(n738) );
  NAND2X1 U346 ( .A(n539), .B(n537), .Y(n793) );
  XNOR2X1 U347 ( .A(n850), .B(n531), .Y(n762) );
  AOI21X1 U348 ( .A0(n833), .A1(n850), .B0(n556), .Y(n837) );
  AOI221X1 U349 ( .A0(n877), .A1(n540), .B0(n555), .B1(n735), .C0(n734), .Y(
        n750) );
  AOI21X1 U350 ( .A0(n536), .A1(n733), .B0(n799), .Y(n734) );
  OAI21XL U351 ( .A0(n861), .A1(n853), .B0(n850), .Y(n733) );
  AOI222X1 U352 ( .A0(n549), .A1(n713), .B0(n712), .B1(n711), .C0(n556), .C1(
        n537), .Y(n732) );
  OAI21XL U353 ( .A0(n850), .A1(n709), .B0(n550), .Y(n712) );
  AOI31X1 U354 ( .A0(n761), .A1(n624), .A2(n623), .B0(n767), .Y(n625) );
  AOI22X1 U355 ( .A0(n775), .A1(n850), .B0(n894), .B1(n554), .Y(n623) );
  AOI31X1 U356 ( .A0(n703), .A1(n793), .A2(n702), .B0(n815), .Y(n704) );
  OAI2BB1X1 U357 ( .A0N(n700), .A1N(n699), .B0(n554), .Y(n703) );
  AOI22X1 U358 ( .A0(n894), .A1(n556), .B0(n701), .B1(n547), .Y(n702) );
  INVX1 U359 ( .A(n830), .Y(n547) );
  INVX1 U360 ( .A(n830), .Y(n549) );
  INVX1 U361 ( .A(n830), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n565) );
  INVX1 U363 ( .A(n840), .Y(n553) );
  INVX1 U364 ( .A(n840), .Y(n554) );
  INVX1 U365 ( .A(n840), .Y(n552) );
  NOR2BX1 U366 ( .AN(n830), .B(n553), .Y(n614) );
  AOI22X1 U367 ( .A0(n581), .A1(a[0]), .B0(n580), .B1(n579), .Y(n582) );
  AOI31X1 U368 ( .A0(n717), .A1(n848), .A2(n571), .B0(n570), .Y(n583) );
  AOI22X1 U369 ( .A0(n576), .A1(n897), .B0(n556), .B1(n833), .Y(n580) );
  AOI22X1 U370 ( .A0(n673), .A1(n902), .B0(n534), .B1(n672), .Y(n674) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n654), .B0(n653), .B1(n848), .Y(n673) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n671), .B0(n670), .B1(n848), .Y(n672) );
  OAI22X1 U373 ( .A0(n698), .A1(n767), .B0(n697), .B1(n769), .Y(n705) );
  AOI221X1 U374 ( .A0(n548), .A1(n693), .B0(n556), .B1(n797), .C0(n692), .Y(
        n698) );
  AOI222X1 U375 ( .A0(n759), .A1(n547), .B0(a[2]), .B1(n696), .C0(n556), .C1(
        n695), .Y(n697) );
  OAI22X1 U376 ( .A0(n888), .A1(n542), .B0(n550), .B1(n537), .Y(n692) );
  NOR2X1 U377 ( .A(n863), .B(n861), .Y(n804) );
  BUFX3 U378 ( .A(n710), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n852), .Y(n710) );
  AOI221X1 U380 ( .A0(n916), .A1(n785), .B0(n851), .B1(n666), .C0(n665), .Y(
        n667) );
  NOR3X1 U381 ( .A(n851), .B(a[7]), .C(n860), .Y(n665) );
  INVX1 U382 ( .A(n762), .Y(n851) );
  OAI21XL U383 ( .A0(n857), .A1(n550), .B0(n664), .Y(n666) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI33X1 U385 ( .A0(n532), .A1(n540), .A2(n904), .B0(n738), .B1(n742), .B2(
        a[2]), .Y(n739) );
  AOI22X1 U386 ( .A0(n882), .A1(n850), .B0(a[2]), .B1(n612), .Y(n613) );
  CLKINVX3 U387 ( .A(a[0]), .Y(n848) );
  AOI211X1 U388 ( .A0(n724), .A1(n578), .B0(n577), .C0(a[0]), .Y(n579) );
  NAND2X1 U389 ( .A(n781), .B(n805), .Y(n578) );
  AOI21X1 U390 ( .A0(n803), .A1(n624), .B0(n897), .Y(n577) );
  BUFX3 U391 ( .A(a[5]), .Y(n533) );
  OAI221XL U392 ( .A0(n536), .A1(n808), .B0(n802), .B1(n545), .C0(n801), .Y(
        n818) );
  AOI22X1 U393 ( .A0(n539), .A1(n800), .B0(n799), .B1(a[2]), .Y(n801) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_9 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916;

  OAI221X4 U4 ( .A0(n857), .A1(n536), .B0(n862), .B1(n551), .C0(n839), .Y(n842) );
  OAI221X4 U6 ( .A0(n837), .A1(n836), .B0(n835), .B1(n551), .C0(n834), .Y(n843) );
  OAI221X4 U28 ( .A0(n883), .A1(n551), .B0(n865), .B1(n545), .C0(n786), .Y(
        n787) );
  OAI221X4 U35 ( .A0(n778), .A1(n545), .B0(n895), .B1(n551), .C0(n777), .Y(
        n779) );
  OAI221X4 U70 ( .A0(n877), .A1(n551), .B0(n860), .B1(n545), .C0(n723), .Y(
        n729) );
  OAI221X4 U103 ( .A0(n551), .A1(n836), .B0(n829), .B1(n819), .C0(n677), .Y(
        n688) );
  OAI221X4 U151 ( .A0(n856), .A1(n551), .B0(n542), .B1(n538), .C0(n629), .Y(
        n641) );
  OAI221X4 U166 ( .A0(n615), .A1(n551), .B0(n545), .B1(n758), .C0(n761), .Y(
        n616) );
  OAI32X4 U280 ( .A0(n551), .A1(n867), .A2(n870), .B0(n542), .B1(n820), .Y(
        n557) );
  AOI221X1 U1 ( .A0(n858), .A1(a[2]), .B0(n826), .B1(n565), .C0(n916), .Y(n566) );
  INVX1 U2 ( .A(a[7]), .Y(n903) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n820) );
  NAND2X2 U5 ( .A(n531), .B(n532), .Y(n808) );
  NAND2X1 U7 ( .A(n867), .B(n531), .Y(n694) );
  NAND2X2 U8 ( .A(n532), .B(n857), .Y(n742) );
  NAND2X1 U9 ( .A(n531), .B(n539), .Y(n803) );
  NAND2X1 U10 ( .A(n884), .B(n531), .Y(n781) );
  NAND2X2 U11 ( .A(n537), .B(n742), .Y(n810) );
  NAND2X2 U12 ( .A(n857), .B(n535), .Y(n807) );
  NAND2X2 U13 ( .A(n857), .B(n852), .Y(n785) );
  NAND2X1 U14 ( .A(n531), .B(n742), .Y(n821) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n850) );
  NAND2X1 U16 ( .A(n533), .B(n848), .Y(n813) );
  CLKINVX3 U17 ( .A(n533), .Y(n897) );
  NAND2X2 U18 ( .A(n848), .B(n897), .Y(n769) );
  NAND2X2 U19 ( .A(a[0]), .B(n897), .Y(n767) );
  OAI22X2 U20 ( .A0(n534), .A1(n643), .B0(n642), .B1(n902), .Y(d[2]) );
  OAI21X2 U21 ( .A0(n847), .A1(n902), .B0(n846), .Y(d[7]) );
  AOI221X1 U22 ( .A0(n899), .A1(n913), .B0(n898), .B1(n818), .C0(n817), .Y(
        n847) );
  OAI22X2 U23 ( .A0(n534), .A1(n708), .B0(n707), .B1(n902), .Y(d[4]) );
  NAND2X1 U24 ( .A(a[2]), .B(n903), .Y(n840) );
  NAND2X1 U25 ( .A(a[7]), .B(n850), .Y(n830) );
  AOI21XL U26 ( .A0(n916), .A1(a[4]), .B0(n907), .Y(n603) );
  OAI222X4 U27 ( .A0(n541), .A1(n805), .B0(n804), .B1(n545), .C0(a[4]), .C1(
        n803), .Y(n806) );
  NAND2X1 U29 ( .A(n531), .B(a[4]), .Y(n699) );
  NAND2X1 U30 ( .A(a[4]), .B(n535), .Y(n660) );
  NAND2X2 U31 ( .A(n532), .B(a[4]), .Y(n812) );
  CLKINVX3 U32 ( .A(a[4]), .Y(n857) );
  NAND2X1 U33 ( .A(n870), .B(n906), .Y(n635) );
  CLKINVX3 U34 ( .A(n541), .Y(n540) );
  INVX1 U36 ( .A(n598), .Y(n889) );
  NAND2X1 U37 ( .A(n810), .B(n535), .Y(n709) );
  NAND2X1 U38 ( .A(n867), .B(n535), .Y(n690) );
  NAND2X1 U39 ( .A(n877), .B(n535), .Y(n714) );
  NAND2X1 U40 ( .A(n873), .B(n535), .Y(n622) );
  NAND2X1 U41 ( .A(n538), .B(n655), .Y(n711) );
  NAND2X1 U42 ( .A(n776), .B(n709), .Y(n716) );
  NAND2X1 U43 ( .A(n808), .B(n714), .Y(n713) );
  INVX1 U44 ( .A(n755), .Y(n861) );
  INVX1 U45 ( .A(n538), .Y(n870) );
  INVX1 U46 ( .A(n741), .Y(n866) );
  NOR2X1 U47 ( .A(n535), .B(n884), .Y(n598) );
  CLKINVX3 U48 ( .A(n555), .Y(n550) );
  NAND2X1 U49 ( .A(n535), .B(n852), .Y(n805) );
  NAND2X1 U50 ( .A(n785), .B(n535), .Y(n700) );
  NAND2X1 U51 ( .A(n884), .B(n535), .Y(n675) );
  NAND2X1 U52 ( .A(n742), .B(n535), .Y(n757) );
  NAND2X1 U53 ( .A(n694), .B(n675), .Y(n836) );
  CLKINVX3 U54 ( .A(n813), .Y(n900) );
  INVX1 U55 ( .A(n821), .Y(n862) );
  NAND2X1 U56 ( .A(n808), .B(n700), .Y(n617) );
  INVX1 U57 ( .A(n693), .Y(n854) );
  INVX1 U58 ( .A(n807), .Y(n859) );
  INVX1 U59 ( .A(n820), .Y(n855) );
  BUFX3 U60 ( .A(n849), .Y(n535) );
  NAND2X1 U61 ( .A(n873), .B(n531), .Y(n776) );
  NAND2X1 U62 ( .A(n812), .B(n535), .Y(n655) );
  NAND2X1 U63 ( .A(n531), .B(n810), .Y(n758) );
  NAND2X1 U64 ( .A(n531), .B(n785), .Y(n741) );
  INVX1 U65 ( .A(n537), .Y(n877) );
  NAND2X1 U66 ( .A(n906), .B(n532), .Y(n664) );
  NAND2X1 U67 ( .A(n812), .B(n776), .Y(n827) );
  NOR2X1 U68 ( .A(n537), .B(n535), .Y(n799) );
  CLKINVX3 U69 ( .A(n812), .Y(n884) );
  NAND2X1 U71 ( .A(n531), .B(n852), .Y(n693) );
  NAND2X1 U72 ( .A(n531), .B(n857), .Y(n586) );
  NAND2BX1 U73 ( .AN(n799), .B(n660), .Y(n727) );
  INVX1 U74 ( .A(n767), .Y(n899) );
  NAND2X1 U75 ( .A(n699), .B(n655), .Y(n782) );
  NAND2BX1 U76 ( .AN(n830), .B(n537), .Y(n624) );
  NAND2X1 U77 ( .A(n699), .B(n690), .Y(n819) );
  NAND2X1 U78 ( .A(n660), .B(n781), .Y(n823) );
  CLKINVX3 U79 ( .A(n534), .Y(n902) );
  CLKINVX3 U80 ( .A(n815), .Y(n901) );
  INVX1 U81 ( .A(n674), .Y(d[3]) );
  BUFX3 U82 ( .A(a[1]), .Y(n531) );
  NAND2X1 U83 ( .A(a[7]), .B(a[2]), .Y(n829) );
  NAND2X1 U84 ( .A(n533), .B(a[0]), .Y(n815) );
  INVX1 U85 ( .A(n685), .Y(n907) );
  NAND2X1 U86 ( .A(n864), .B(n540), .Y(n809) );
  NAND2X1 U87 ( .A(n872), .B(n556), .Y(n685) );
  INVX1 U88 ( .A(n635), .Y(n908) );
  NOR2X1 U89 ( .A(n550), .B(n598), .Y(n724) );
  NOR2X1 U90 ( .A(n874), .B(n861), .Y(n676) );
  NAND2X1 U91 ( .A(n701), .B(n540), .Y(n761) );
  INVX1 U92 ( .A(n622), .Y(n874) );
  INVX1 U93 ( .A(n675), .Y(n886) );
  INVX1 U94 ( .A(n757), .Y(n863) );
  INVX1 U95 ( .A(n716), .Y(n875) );
  INVX1 U96 ( .A(n695), .Y(n872) );
  INVX4 U97 ( .A(n536), .Y(n556) );
  NOR2BX1 U98 ( .AN(n709), .B(n854), .Y(n835) );
  NOR2X1 U99 ( .A(n870), .B(n853), .Y(n597) );
  AOI22X1 U100 ( .A0(n900), .A1(n788), .B0(n898), .B1(n787), .Y(n789) );
  OAI221XL U101 ( .A0(n887), .A1(n550), .B0(n802), .B1(n543), .C0(n783), .Y(
        n788) );
  INVX1 U102 ( .A(n838), .Y(n887) );
  NOR2X1 U104 ( .A(n873), .B(n862), .Y(n637) );
  NAND2X1 U105 ( .A(n889), .B(n700), .Y(n740) );
  INVX1 U106 ( .A(n805), .Y(n853) );
  NAND2X1 U107 ( .A(n889), .B(n675), .Y(n800) );
  INVX1 U108 ( .A(n690), .Y(n868) );
  INVX1 U109 ( .A(n700), .Y(n864) );
  NOR2X1 U110 ( .A(n866), .B(n868), .Y(n726) );
  OAI221XL U111 ( .A0(n865), .A1(n545), .B0(n825), .B1(n829), .C0(n905), .Y(
        n576) );
  INVX1 U112 ( .A(n724), .Y(n905) );
  INVX1 U113 ( .A(n796), .Y(n888) );
  NOR2X1 U114 ( .A(n864), .B(n854), .Y(n825) );
  INVX1 U115 ( .A(n711), .Y(n882) );
  INVX1 U116 ( .A(n617), .Y(n865) );
  INVX1 U117 ( .A(n765), .Y(n881) );
  INVX1 U118 ( .A(n836), .Y(n885) );
  INVX1 U119 ( .A(n713), .Y(n879) );
  NAND2X1 U120 ( .A(n860), .B(n535), .Y(n680) );
  OAI22X1 U121 ( .A0(n683), .A1(n813), .B0(n682), .B1(n769), .Y(n687) );
  AOI222X1 U122 ( .A0(n862), .A1(n548), .B0(n556), .B1(n679), .C0(n678), .C1(
        n711), .Y(n683) );
  AOI211X1 U123 ( .A0(n556), .A1(n689), .B0(n681), .C0(n724), .Y(n682) );
  NAND2X1 U124 ( .A(n807), .B(n694), .Y(n679) );
  NOR2X1 U125 ( .A(n877), .B(n866), .Y(n701) );
  OAI22X1 U126 ( .A0(n829), .A1(n716), .B0(n545), .B1(n538), .Y(n681) );
  CLKINVX3 U127 ( .A(n810), .Y(n873) );
  CLKINVX3 U128 ( .A(n742), .Y(n860) );
  AOI22X1 U129 ( .A0(n899), .A1(n832), .B0(n900), .B1(n831), .Y(n845) );
  OAI221XL U130 ( .A0(n825), .A1(n545), .B0(n893), .B1(n543), .C0(n824), .Y(
        n832) );
  OAI221XL U131 ( .A0(n881), .A1(n545), .B0(n872), .B1(n543), .C0(n828), .Y(
        n831) );
  INVX1 U132 ( .A(n819), .Y(n893) );
  NAND2X1 U133 ( .A(n556), .B(n827), .Y(n736) );
  NAND2X1 U134 ( .A(n808), .B(n709), .Y(n695) );
  AOI22X1 U135 ( .A0(n900), .A1(n729), .B0(n901), .B1(n728), .Y(n730) );
  OAI221XL U136 ( .A0(n536), .A1(n727), .B0(n726), .B1(n545), .C0(n725), .Y(
        n728) );
  AOI211X1 U137 ( .A0(n722), .A1(n556), .B0(n721), .C0(n720), .Y(n723) );
  AOI22X1 U138 ( .A0(n900), .A1(n592), .B0(n901), .B1(n591), .Y(n593) );
  OAI221XL U139 ( .A0(n888), .A1(n545), .B0(n879), .B1(n543), .C0(n590), .Y(
        n591) );
  OAI211X1 U140 ( .A0(n597), .A1(n550), .B0(n635), .C0(n589), .Y(n592) );
  AOI22X1 U141 ( .A0(n888), .A1(n556), .B0(n884), .B1(n552), .Y(n590) );
  AOI22X1 U142 ( .A0(n548), .A1(n860), .B0(n676), .B1(n539), .Y(n589) );
  AOI21X1 U143 ( .A0(n808), .A1(n680), .B0(n550), .Y(n563) );
  INVX1 U144 ( .A(n803), .Y(n916) );
  AND2X2 U145 ( .A(n758), .B(n757), .Y(n794) );
  OAI21XL U146 ( .A0(n758), .A1(n550), .B0(n736), .Y(n657) );
  INVX1 U147 ( .A(n639), .Y(n911) );
  OAI31X1 U148 ( .A0(n721), .A1(n908), .A2(n638), .B0(n898), .Y(n639) );
  OAI21XL U149 ( .A0(n541), .A1(n637), .B0(n636), .Y(n638) );
  INVX1 U150 ( .A(n776), .Y(n876) );
  OAI22X1 U152 ( .A0(n621), .A1(n769), .B0(n620), .B1(n813), .Y(n626) );
  AOI211X1 U153 ( .A0(n556), .A1(n821), .B0(n619), .C0(n618), .Y(n620) );
  AOI221X1 U154 ( .A0(n910), .A1(n535), .B0(n896), .B1(n556), .C0(n616), .Y(
        n621) );
  OAI22X1 U155 ( .A0(n859), .A1(n543), .B0(n550), .B1(n617), .Y(n619) );
  AOI222X1 U156 ( .A0(n867), .A1(n540), .B0(n863), .B1(n554), .C0(n547), .C1(
        n852), .Y(n567) );
  AOI21X1 U157 ( .A0(n873), .A1(n556), .B0(n557), .Y(n558) );
  AOI2BB2X1 U158 ( .B0(n910), .B1(n535), .A0N(n536), .A1N(n676), .Y(n677) );
  CLKINVX8 U159 ( .A(n546), .Y(n545) );
  CLKINVX3 U160 ( .A(n541), .Y(n539) );
  NOR2X1 U161 ( .A(n545), .B(n535), .Y(n721) );
  AOI222X1 U162 ( .A0(n916), .A1(n810), .B0(n724), .B1(n873), .C0(n886), .C1(
        n540), .Y(n725) );
  AOI221X1 U163 ( .A0(n602), .A1(n553), .B0(n540), .B1(n612), .C0(n596), .Y(
        n608) );
  OAI221XL U164 ( .A0(n536), .A1(n714), .B0(n545), .B1(n820), .C0(n635), .Y(
        n596) );
  AOI221X1 U165 ( .A0(n916), .A1(n852), .B0(n553), .B1(n810), .C0(n737), .Y(
        n749) );
  OAI2BB1X1 U167 ( .A0N(n781), .A1N(n548), .B0(n736), .Y(n737) );
  NOR2X1 U168 ( .A(n854), .B(n855), .Y(n615) );
  OAI221XL U169 ( .A0(n869), .A1(n545), .B0(n890), .B1(n543), .C0(n691), .Y(
        n706) );
  INVX1 U170 ( .A(n689), .Y(n869) );
  AOI32X1 U171 ( .A0(n889), .A1(n742), .A2(n556), .B0(n553), .B1(n690), .Y(
        n691) );
  INVX1 U172 ( .A(n808), .Y(n856) );
  AOI211X1 U173 ( .A0(n875), .A1(n556), .B0(n914), .C0(n628), .Y(n629) );
  INVX1 U174 ( .A(n809), .Y(n914) );
  AOI211X1 U175 ( .A0(n863), .A1(n540), .B0(n909), .C0(n559), .Y(n560) );
  NOR3X1 U176 ( .A(n545), .B(n884), .C(n862), .Y(n559) );
  INVX1 U177 ( .A(n664), .Y(n909) );
  OAI221XL U178 ( .A0(n536), .A1(n755), .B0(n759), .B1(n551), .C0(n754), .Y(
        n773) );
  AOI22X1 U179 ( .A0(n549), .A1(n889), .B0(n875), .B1(n539), .Y(n754) );
  AOI211X1 U180 ( .A0(n554), .A1(n827), .B0(n908), .C0(n826), .Y(n828) );
  AOI211X1 U181 ( .A0(n878), .A1(n540), .B0(n719), .C0(n718), .Y(n731) );
  INVX1 U182 ( .A(n714), .Y(n878) );
  NAND2BX1 U183 ( .AN(n826), .B(n717), .Y(n718) );
  OAI222X1 U184 ( .A0(n551), .A1(n716), .B0(n742), .B1(n803), .C0(n545), .C1(
        n715), .Y(n719) );
  CLKINVX3 U185 ( .A(n555), .Y(n551) );
  INVX1 U186 ( .A(n798), .Y(n913) );
  AOI221X1 U187 ( .A0(n797), .A1(n552), .B0(n796), .B1(n549), .C0(n795), .Y(
        n798) );
  OAI21XL U188 ( .A0(n536), .A1(n794), .B0(n793), .Y(n795) );
  INVX1 U189 ( .A(n536), .Y(n906) );
  NOR2X1 U190 ( .A(n884), .B(n866), .Y(n744) );
  NAND3X1 U191 ( .A(n538), .B(n810), .C(n540), .Y(n834) );
  NAND2X1 U192 ( .A(n709), .B(n781), .Y(n833) );
  NAND2X1 U193 ( .A(n807), .B(n781), .Y(n838) );
  NAND2X1 U194 ( .A(n808), .B(n655), .Y(n765) );
  NAND2X1 U195 ( .A(n538), .B(n757), .Y(n612) );
  NOR2BX1 U196 ( .AN(n694), .B(n855), .Y(n759) );
  AOI21X1 U197 ( .A0(n742), .A1(n741), .B0(n536), .Y(n743) );
  AOI22X1 U198 ( .A0(n874), .A1(n548), .B0(n556), .B1(n782), .Y(n783) );
  AOI22X1 U199 ( .A0(n866), .A1(n546), .B0(n555), .B1(n810), .Y(n684) );
  AOI22X1 U200 ( .A0(n547), .A1(n612), .B0(n873), .B1(n539), .Y(n573) );
  NOR2X1 U201 ( .A(n785), .B(n536), .Y(n826) );
  NAND2X1 U202 ( .A(n680), .B(n781), .Y(n796) );
  INVX1 U203 ( .A(n769), .Y(n898) );
  NAND2X1 U204 ( .A(n694), .B(n680), .Y(n689) );
  CLKINVX3 U205 ( .A(n785), .Y(n867) );
  NAND2X1 U206 ( .A(n694), .B(n714), .Y(n663) );
  NOR2X1 U207 ( .A(n859), .B(n799), .Y(n802) );
  AOI211X1 U208 ( .A0(n556), .A1(n617), .B0(n588), .C0(n587), .Y(n594) );
  OAI2BB2X1 U209 ( .B0(n545), .B1(n740), .A0N(n735), .A1N(n540), .Y(n588) );
  AOI21X1 U210 ( .A0(n622), .A1(n586), .B0(n550), .Y(n587) );
  NAND2X1 U211 ( .A(n538), .B(n709), .Y(n797) );
  NAND2X1 U212 ( .A(n785), .B(n821), .Y(n696) );
  NAND2X1 U213 ( .A(n820), .B(n758), .Y(n735) );
  AOI21X1 U214 ( .A0(n556), .A1(n823), .B0(n822), .Y(n824) );
  AOI21X1 U215 ( .A0(n821), .A1(n820), .B0(n550), .Y(n822) );
  OAI221XL U216 ( .A0(n858), .A1(n551), .B0(n892), .B1(n536), .C0(n774), .Y(
        n780) );
  AOI2BB2X1 U217 ( .B0(n539), .B1(n836), .A0N(n545), .A1N(n802), .Y(n774) );
  INVX1 U218 ( .A(n586), .Y(n858) );
  INVX1 U219 ( .A(n715), .Y(n894) );
  INVX1 U220 ( .A(n624), .Y(n910) );
  INVX1 U221 ( .A(n823), .Y(n890) );
  AOI221XL U222 ( .A0(n556), .A1(n871), .B0(n548), .B1(n800), .C0(n599), .Y(
        n607) );
  INVX1 U223 ( .A(n597), .Y(n871) );
  OAI32X1 U224 ( .A0(n542), .A1(n860), .A2(n598), .B0(n886), .B1(n551), .Y(
        n599) );
  INVX1 U225 ( .A(n727), .Y(n892) );
  OAI221XL U226 ( .A0(n867), .A1(n545), .B0(n891), .B1(n542), .C0(n760), .Y(
        n772) );
  INVX1 U227 ( .A(n756), .Y(n891) );
  AOI22X1 U228 ( .A0(n759), .A1(n556), .B0(n794), .B1(n552), .Y(n760) );
  INVX1 U229 ( .A(n782), .Y(n896) );
  INVX1 U230 ( .A(n827), .Y(n883) );
  AOI31X1 U231 ( .A0(n821), .A1(n785), .A2(n556), .B0(n912), .Y(n786) );
  INVX1 U232 ( .A(n834), .Y(n912) );
  INVX1 U233 ( .A(n738), .Y(n904) );
  INVX1 U234 ( .A(n540), .Y(n542) );
  INVX1 U235 ( .A(n540), .Y(n543) );
  AOI211X1 U236 ( .A0(n901), .A1(n627), .B0(n626), .C0(n625), .Y(n643) );
  AOI211X1 U237 ( .A0(n901), .A1(n641), .B0(n640), .C0(n911), .Y(n642) );
  OAI2BB2X1 U238 ( .B0(n614), .B1(n613), .A0N(n744), .A1N(n614), .Y(n627) );
  AOI211X1 U239 ( .A0(n901), .A1(n688), .B0(n687), .C0(n686), .Y(n708) );
  AOI211X1 U240 ( .A0(n900), .A1(n706), .B0(n705), .C0(n704), .Y(n707) );
  AOI31X1 U241 ( .A0(n685), .A1(n793), .A2(n684), .B0(n767), .Y(n686) );
  OAI21X2 U242 ( .A0(n534), .A1(n792), .B0(n791), .Y(d[6]) );
  OAI2BB1X1 U243 ( .A0N(n790), .A1N(n789), .B0(n534), .Y(n791) );
  AOI221X1 U244 ( .A0(n900), .A1(n773), .B0(n901), .B1(n772), .C0(n771), .Y(
        n792) );
  AOI22X1 U245 ( .A0(n899), .A1(n780), .B0(n901), .B1(n779), .Y(n790) );
  OAI2BB1X1 U246 ( .A0N(n845), .A1N(n844), .B0(n902), .Y(n846) );
  AOI22X1 U247 ( .A0(n901), .A1(n843), .B0(n898), .B1(n842), .Y(n844) );
  AOI22X1 U248 ( .A0(n533), .A1(n669), .B0(n668), .B1(n897), .Y(n670) );
  OAI221XL U249 ( .A0(n862), .A1(n551), .B0(n545), .B1(n663), .C0(n662), .Y(
        n669) );
  OAI221XL U250 ( .A0(n882), .A1(n545), .B0(n543), .B1(n742), .C0(n667), .Y(
        n668) );
  AOI21X1 U251 ( .A0(n890), .A1(n906), .B0(n661), .Y(n662) );
  AOI22X1 U252 ( .A0(n575), .A1(n897), .B0(n533), .B1(n574), .Y(n581) );
  OAI221XL U253 ( .A0(n536), .A1(n757), .B0(n637), .B1(n545), .C0(n572), .Y(
        n575) );
  OAI211X1 U254 ( .A0(n835), .A1(n550), .B0(n736), .C0(n573), .Y(n574) );
  AOI2BB2X1 U255 ( .B0(n539), .B1(n727), .A0N(n550), .A1N(n744), .Y(n572) );
  OAI22X1 U256 ( .A0(n634), .A1(n813), .B0(n633), .B1(n767), .Y(n640) );
  AOI221XL U257 ( .A0(n549), .A1(n740), .B0(n799), .B1(n850), .C0(n632), .Y(
        n633) );
  AOI221XL U258 ( .A0(n867), .A1(n916), .B0(n547), .B1(n713), .C0(n630), .Y(
        n634) );
  OAI32X1 U259 ( .A0(n738), .A1(n860), .A2(n850), .B0(n631), .B1(n904), .Y(
        n632) );
  OAI22X1 U260 ( .A0(n770), .A1(n769), .B0(n768), .B1(n767), .Y(n771) );
  AOI211X1 U261 ( .A0(n881), .A1(n850), .B0(n766), .C0(n907), .Y(n768) );
  AOI221XL U262 ( .A0(n862), .A1(n554), .B0(n547), .B1(n776), .C0(n764), .Y(
        n770) );
  OAI22X1 U263 ( .A0(n542), .A1(n852), .B0(n886), .B1(n550), .Y(n766) );
  OAI22X1 U264 ( .A0(n816), .A1(n815), .B0(n814), .B1(n813), .Y(n817) );
  AOI221XL U265 ( .A0(n549), .A1(n812), .B0(n876), .B1(n540), .C0(n811), .Y(
        n814) );
  AOI221X1 U266 ( .A0(n556), .A1(n808), .B0(n553), .B1(n807), .C0(n806), .Y(
        n816) );
  OAI221XL U267 ( .A0(n536), .A1(n810), .B0(n879), .B1(n551), .C0(n809), .Y(
        n811) );
  AOI211X1 U268 ( .A0(n868), .A1(n556), .B0(n652), .C0(n651), .Y(n653) );
  AOI31X1 U269 ( .A0(n809), .A1(n717), .A2(n650), .B0(n533), .Y(n651) );
  OAI22X1 U270 ( .A0(n857), .A1(n803), .B0(n649), .B1(n897), .Y(n652) );
  AOI2BB2X1 U271 ( .B0(n853), .B1(n554), .A0N(n833), .A1N(n545), .Y(n650) );
  AOI2BB2X1 U272 ( .B0(n659), .B1(n897), .A0N(n897), .A1N(n658), .Y(n671) );
  OAI221XL U273 ( .A0(n877), .A1(n551), .B0(n545), .B1(n807), .C0(n656), .Y(
        n659) );
  AOI221XL U274 ( .A0(n548), .A1(n676), .B0(n711), .B1(n540), .C0(n657), .Y(
        n658) );
  AOI22X1 U275 ( .A0(n539), .A1(n765), .B0(n873), .B1(n903), .Y(n656) );
  AOI22X1 U276 ( .A0(n554), .A1(n532), .B0(n539), .B1(n857), .Y(n631) );
  AOI22X1 U277 ( .A0(n900), .A1(n747), .B0(n899), .B1(n746), .Y(n748) );
  OAI221XL U278 ( .A0(n860), .A1(n545), .B0(n542), .B1(n807), .C0(n745), .Y(
        n746) );
  OAI221XL U279 ( .A0(n885), .A1(n536), .B0(n545), .B1(n740), .C0(n739), .Y(
        n747) );
  AOI21X1 U281 ( .A0(n744), .A1(n552), .B0(n743), .Y(n745) );
  AOI22X1 U282 ( .A0(n533), .A1(n562), .B0(n561), .B1(n897), .Y(n571) );
  OAI221XL U283 ( .A0(n880), .A1(n545), .B0(n541), .B1(n889), .C0(n558), .Y(
        n562) );
  OAI221XL U284 ( .A0(n532), .A1(n803), .B0(n722), .B1(n551), .C0(n560), .Y(
        n561) );
  INVX1 U285 ( .A(n663), .Y(n880) );
  AOI22X1 U286 ( .A0(n901), .A1(n605), .B0(n900), .B1(n604), .Y(n606) );
  OAI21XL U287 ( .A0(n602), .A1(n536), .B0(n601), .Y(n605) );
  OAI221XL U288 ( .A0(n551), .A1(n810), .B0(n835), .B1(n545), .C0(n603), .Y(
        n604) );
  AOI31X1 U289 ( .A0(n538), .A1(n742), .A2(n600), .B0(n910), .Y(n601) );
  INVX1 U290 ( .A(n611), .Y(d[1]) );
  AOI22X1 U291 ( .A0(n534), .A1(n610), .B0(n609), .B1(n902), .Y(n611) );
  OAI221XL U292 ( .A0(n595), .A1(n767), .B0(n594), .B1(n769), .C0(n593), .Y(
        n610) );
  OAI221XL U293 ( .A0(n608), .A1(n767), .B0(n607), .B1(n769), .C0(n606), .Y(
        n609) );
  INVX1 U294 ( .A(n753), .Y(d[5]) );
  AOI22X1 U295 ( .A0(n752), .A1(n902), .B0(n534), .B1(n751), .Y(n753) );
  OAI221XL U296 ( .A0(n750), .A1(n815), .B0(n749), .B1(n769), .C0(n748), .Y(
        n751) );
  OAI221XL U297 ( .A0(n732), .A1(n769), .B0(n731), .B1(n767), .C0(n730), .Y(
        n752) );
  CLKINVX3 U298 ( .A(n532), .Y(n852) );
  OAI21XL U299 ( .A0(n545), .A1(n537), .B0(n803), .Y(n647) );
  NAND2X1 U300 ( .A(n860), .B(n531), .Y(n755) );
  AOI21X1 U301 ( .A0(n699), .A1(n680), .B0(n545), .Y(n628) );
  INVX1 U302 ( .A(n531), .Y(n849) );
  OAI21XL U303 ( .A0(n850), .A1(n622), .B0(n550), .Y(n600) );
  OAI21XL U304 ( .A0(n536), .A1(n805), .B0(n763), .Y(n764) );
  AOI31X1 U305 ( .A0(n812), .A1(n903), .A2(n762), .B0(n915), .Y(n763) );
  INVX1 U306 ( .A(n761), .Y(n915) );
  AOI211X1 U307 ( .A0(n884), .A1(n540), .B0(n648), .C0(n647), .Y(n649) );
  OAI222X1 U308 ( .A0(n551), .A1(n807), .B0(n850), .B1(n693), .C0(n545), .C1(
        n821), .Y(n648) );
  NAND2X1 U309 ( .A(n861), .B(n552), .Y(n636) );
  NOR2BX1 U310 ( .AN(n660), .B(n876), .Y(n722) );
  BUFX3 U311 ( .A(n841), .Y(n536) );
  NAND2X1 U312 ( .A(n850), .B(n903), .Y(n841) );
  OAI221XL U313 ( .A0(n531), .A1(n664), .B0(n829), .B1(n709), .C0(n636), .Y(
        n630) );
  BUFX3 U314 ( .A(n784), .Y(n538) );
  NAND2X1 U315 ( .A(n531), .B(n537), .Y(n784) );
  AOI211X1 U316 ( .A0(n540), .A1(n852), .B0(n585), .C0(n647), .Y(n595) );
  OAI222X1 U317 ( .A0(n551), .A1(n756), .B0(n584), .B1(n536), .C0(n545), .C1(
        n889), .Y(n585) );
  AOI21X1 U318 ( .A0(n537), .A1(n535), .B0(n858), .Y(n584) );
  AOI211X1 U319 ( .A0(n533), .A1(n569), .B0(n848), .C0(n568), .Y(n570) );
  OAI221XL U320 ( .A0(n545), .A1(n807), .B0(n602), .B1(n829), .C0(n564), .Y(
        n569) );
  AOI21X1 U321 ( .A0(n567), .A1(n566), .B0(n533), .Y(n568) );
  AOI31X1 U322 ( .A0(n556), .A1(n565), .A2(n884), .B0(n563), .Y(n564) );
  INVX1 U323 ( .A(n830), .Y(n546) );
  INVX1 U324 ( .A(n840), .Y(n554) );
  INVX1 U325 ( .A(n840), .Y(n555) );
  INVX1 U326 ( .A(n544), .Y(n541) );
  INVX1 U327 ( .A(n829), .Y(n544) );
  AOI22X1 U328 ( .A0(n533), .A1(n646), .B0(n645), .B1(n897), .Y(n654) );
  OAI222X1 U329 ( .A0(n545), .A1(n782), .B0(n551), .B1(n660), .C0(n894), .C1(
        n542), .Y(n646) );
  OAI221XL U330 ( .A0(n892), .A1(n536), .B0(n551), .B1(n819), .C0(n644), .Y(
        n645) );
  AOI2BB2X1 U331 ( .B0(n835), .B1(n539), .A0N(n545), .A1N(n726), .Y(n644) );
  NAND2X1 U332 ( .A(n699), .B(n622), .Y(n775) );
  NOR2BX1 U333 ( .AN(n660), .B(n862), .Y(n602) );
  AOI21X1 U334 ( .A0(n690), .A1(n758), .B0(n903), .Y(n661) );
  AOI22X1 U335 ( .A0(n549), .A1(n838), .B0(n882), .B1(n539), .Y(n839) );
  AOI31X1 U336 ( .A0(n703), .A1(n793), .A2(n702), .B0(n815), .Y(n704) );
  OAI2BB1X1 U337 ( .A0N(n700), .A1N(n699), .B0(n553), .Y(n703) );
  AOI22X1 U338 ( .A0(n894), .A1(n556), .B0(n701), .B1(n547), .Y(n702) );
  NAND2X1 U339 ( .A(n699), .B(n805), .Y(n715) );
  NAND2X1 U340 ( .A(n660), .B(n586), .Y(n756) );
  AOI21X1 U341 ( .A0(n660), .A1(n741), .B0(n545), .Y(n618) );
  AOI21X1 U342 ( .A0(n812), .A1(n538), .B0(n829), .Y(n720) );
  NAND2X1 U343 ( .A(n906), .B(n531), .Y(n717) );
  OAI21XL U344 ( .A0(n850), .A1(n680), .B0(n550), .Y(n678) );
  XNOR2X1 U345 ( .A(n903), .B(n531), .Y(n738) );
  NAND2X1 U346 ( .A(n539), .B(n537), .Y(n793) );
  XNOR2X1 U347 ( .A(n850), .B(n531), .Y(n762) );
  AOI21X1 U348 ( .A0(n833), .A1(n850), .B0(n556), .Y(n837) );
  AOI221X1 U349 ( .A0(n877), .A1(n540), .B0(n552), .B1(n735), .C0(n734), .Y(
        n750) );
  AOI21X1 U350 ( .A0(n536), .A1(n733), .B0(n799), .Y(n734) );
  OAI21XL U351 ( .A0(n861), .A1(n853), .B0(n850), .Y(n733) );
  AOI222X1 U352 ( .A0(n549), .A1(n713), .B0(n712), .B1(n711), .C0(n556), .C1(
        n537), .Y(n732) );
  OAI21XL U353 ( .A0(n850), .A1(n709), .B0(n550), .Y(n712) );
  NOR2X1 U354 ( .A(n861), .B(n868), .Y(n778) );
  AOI22X1 U355 ( .A0(n906), .A1(n857), .B0(n539), .B1(n776), .Y(n777) );
  INVX1 U356 ( .A(n775), .Y(n895) );
  AOI31X1 U357 ( .A0(n761), .A1(n624), .A2(n623), .B0(n767), .Y(n625) );
  AOI22X1 U358 ( .A0(n775), .A1(n850), .B0(n894), .B1(n553), .Y(n623) );
  INVX1 U359 ( .A(n830), .Y(n547) );
  INVX1 U360 ( .A(n830), .Y(n549) );
  INVX1 U361 ( .A(n830), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n565) );
  INVX1 U363 ( .A(n840), .Y(n552) );
  INVX1 U364 ( .A(n840), .Y(n553) );
  NOR2BX1 U365 ( .AN(n830), .B(n554), .Y(n614) );
  OAI22X2 U366 ( .A0(n583), .A1(n902), .B0(n534), .B1(n582), .Y(d[0]) );
  AOI22X1 U367 ( .A0(n581), .A1(a[0]), .B0(n580), .B1(n579), .Y(n582) );
  AOI31X1 U368 ( .A0(n717), .A1(n848), .A2(n571), .B0(n570), .Y(n583) );
  AOI22X1 U369 ( .A0(n576), .A1(n897), .B0(n556), .B1(n833), .Y(n580) );
  AOI22X1 U370 ( .A0(n673), .A1(n902), .B0(n534), .B1(n672), .Y(n674) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n654), .B0(n653), .B1(n848), .Y(n673) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n671), .B0(n670), .B1(n848), .Y(n672) );
  OAI22X1 U373 ( .A0(n698), .A1(n767), .B0(n697), .B1(n769), .Y(n705) );
  AOI221X1 U374 ( .A0(n548), .A1(n693), .B0(n556), .B1(n797), .C0(n692), .Y(
        n698) );
  AOI222X1 U375 ( .A0(n759), .A1(n547), .B0(a[2]), .B1(n696), .C0(n556), .C1(
        n695), .Y(n697) );
  OAI22X1 U376 ( .A0(n888), .A1(n543), .B0(n550), .B1(n537), .Y(n692) );
  NOR2X1 U377 ( .A(n863), .B(n861), .Y(n804) );
  BUFX3 U378 ( .A(n710), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n852), .Y(n710) );
  AOI221X1 U380 ( .A0(n916), .A1(n785), .B0(n851), .B1(n666), .C0(n665), .Y(
        n667) );
  NOR3X1 U381 ( .A(n851), .B(a[7]), .C(n860), .Y(n665) );
  INVX1 U382 ( .A(n762), .Y(n851) );
  OAI21XL U383 ( .A0(n857), .A1(n550), .B0(n664), .Y(n666) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI33X1 U385 ( .A0(n532), .A1(n540), .A2(n904), .B0(n738), .B1(n742), .B2(
        a[2]), .Y(n739) );
  AOI22X1 U386 ( .A0(n882), .A1(n850), .B0(a[2]), .B1(n612), .Y(n613) );
  CLKINVX3 U387 ( .A(a[0]), .Y(n848) );
  AOI211X1 U388 ( .A0(n724), .A1(n578), .B0(n577), .C0(a[0]), .Y(n579) );
  NAND2X1 U389 ( .A(n781), .B(n805), .Y(n578) );
  AOI21X1 U390 ( .A0(n803), .A1(n624), .B0(n897), .Y(n577) );
  BUFX3 U391 ( .A(a[5]), .Y(n533) );
  OAI221XL U392 ( .A0(n536), .A1(n808), .B0(n802), .B1(n545), .C0(n801), .Y(
        n818) );
  AOI22X1 U393 ( .A0(n539), .A1(n800), .B0(n799), .B1(a[2]), .Y(n801) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_11 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916;

  OAI221X4 U4 ( .A0(n857), .A1(n536), .B0(n862), .B1(n551), .C0(n839), .Y(n842) );
  OAI221X4 U6 ( .A0(n837), .A1(n836), .B0(n835), .B1(n551), .C0(n834), .Y(n843) );
  OAI221X4 U28 ( .A0(n883), .A1(n551), .B0(n865), .B1(n545), .C0(n786), .Y(
        n787) );
  OAI221X4 U35 ( .A0(n778), .A1(n545), .B0(n895), .B1(n551), .C0(n777), .Y(
        n779) );
  OAI221X4 U70 ( .A0(n877), .A1(n551), .B0(n860), .B1(n545), .C0(n723), .Y(
        n729) );
  OAI221X4 U103 ( .A0(n551), .A1(n836), .B0(n829), .B1(n819), .C0(n677), .Y(
        n688) );
  OAI221X4 U151 ( .A0(n856), .A1(n551), .B0(n542), .B1(n538), .C0(n629), .Y(
        n641) );
  OAI221X4 U166 ( .A0(n615), .A1(n551), .B0(n545), .B1(n758), .C0(n761), .Y(
        n616) );
  OAI32X4 U280 ( .A0(n551), .A1(n867), .A2(n870), .B0(n542), .B1(n820), .Y(
        n557) );
  AOI221X1 U1 ( .A0(n858), .A1(a[2]), .B0(n826), .B1(n565), .C0(n916), .Y(n566) );
  INVX1 U2 ( .A(a[7]), .Y(n903) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n820) );
  NAND2X2 U5 ( .A(n531), .B(n532), .Y(n808) );
  NAND2X1 U7 ( .A(n867), .B(n531), .Y(n694) );
  NAND2X2 U8 ( .A(n532), .B(n857), .Y(n742) );
  NAND2X1 U9 ( .A(n531), .B(n539), .Y(n803) );
  NAND2X1 U10 ( .A(n884), .B(n531), .Y(n781) );
  NAND2X2 U11 ( .A(n537), .B(n742), .Y(n810) );
  NAND2X2 U12 ( .A(n857), .B(n535), .Y(n807) );
  NAND2X2 U13 ( .A(n857), .B(n852), .Y(n785) );
  NAND2X1 U14 ( .A(n531), .B(n742), .Y(n821) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n850) );
  NAND2X1 U16 ( .A(n533), .B(n848), .Y(n813) );
  CLKINVX3 U17 ( .A(n533), .Y(n897) );
  NAND2X2 U18 ( .A(n848), .B(n897), .Y(n769) );
  NAND2X2 U19 ( .A(a[0]), .B(n897), .Y(n767) );
  OAI22X2 U20 ( .A0(n534), .A1(n643), .B0(n642), .B1(n902), .Y(d[2]) );
  OAI21X2 U21 ( .A0(n847), .A1(n902), .B0(n846), .Y(d[7]) );
  AOI221X1 U22 ( .A0(n899), .A1(n913), .B0(n898), .B1(n818), .C0(n817), .Y(
        n847) );
  OAI22X2 U23 ( .A0(n534), .A1(n708), .B0(n707), .B1(n902), .Y(d[4]) );
  NAND2X1 U24 ( .A(a[2]), .B(n903), .Y(n840) );
  NAND2X1 U25 ( .A(a[7]), .B(n850), .Y(n830) );
  AOI21XL U26 ( .A0(n916), .A1(a[4]), .B0(n907), .Y(n603) );
  OAI222X4 U27 ( .A0(n541), .A1(n805), .B0(n804), .B1(n545), .C0(a[4]), .C1(
        n803), .Y(n806) );
  NAND2X1 U29 ( .A(n531), .B(a[4]), .Y(n699) );
  NAND2X1 U30 ( .A(a[4]), .B(n535), .Y(n660) );
  NAND2X2 U31 ( .A(n532), .B(a[4]), .Y(n812) );
  CLKINVX3 U32 ( .A(a[4]), .Y(n857) );
  NAND2X1 U33 ( .A(n870), .B(n906), .Y(n635) );
  CLKINVX3 U34 ( .A(n541), .Y(n540) );
  INVX1 U36 ( .A(n598), .Y(n889) );
  NAND2X1 U37 ( .A(n810), .B(n535), .Y(n709) );
  NAND2X1 U38 ( .A(n867), .B(n535), .Y(n690) );
  NAND2X1 U39 ( .A(n877), .B(n535), .Y(n714) );
  NAND2X1 U40 ( .A(n873), .B(n535), .Y(n622) );
  NAND2X1 U41 ( .A(n538), .B(n655), .Y(n711) );
  NAND2X1 U42 ( .A(n776), .B(n709), .Y(n716) );
  NAND2X1 U43 ( .A(n808), .B(n714), .Y(n713) );
  INVX1 U44 ( .A(n755), .Y(n861) );
  INVX1 U45 ( .A(n538), .Y(n870) );
  INVX1 U46 ( .A(n741), .Y(n866) );
  NOR2X1 U47 ( .A(n535), .B(n884), .Y(n598) );
  CLKINVX3 U48 ( .A(n555), .Y(n550) );
  NAND2X1 U49 ( .A(n535), .B(n852), .Y(n805) );
  NAND2X1 U50 ( .A(n785), .B(n535), .Y(n700) );
  NAND2X1 U51 ( .A(n884), .B(n535), .Y(n675) );
  NAND2X1 U52 ( .A(n742), .B(n535), .Y(n757) );
  NAND2X1 U53 ( .A(n694), .B(n675), .Y(n836) );
  CLKINVX3 U54 ( .A(n813), .Y(n900) );
  INVX1 U55 ( .A(n821), .Y(n862) );
  NAND2X1 U56 ( .A(n808), .B(n700), .Y(n617) );
  INVX1 U57 ( .A(n693), .Y(n854) );
  INVX1 U58 ( .A(n807), .Y(n859) );
  INVX1 U59 ( .A(n820), .Y(n855) );
  BUFX3 U60 ( .A(n849), .Y(n535) );
  NAND2X1 U61 ( .A(n873), .B(n531), .Y(n776) );
  NAND2X1 U62 ( .A(n812), .B(n535), .Y(n655) );
  NAND2X1 U63 ( .A(n531), .B(n810), .Y(n758) );
  NAND2X1 U64 ( .A(n531), .B(n785), .Y(n741) );
  INVX1 U65 ( .A(n537), .Y(n877) );
  NAND2X1 U66 ( .A(n906), .B(n532), .Y(n664) );
  NAND2X1 U67 ( .A(n812), .B(n776), .Y(n827) );
  NOR2X1 U68 ( .A(n537), .B(n535), .Y(n799) );
  CLKINVX3 U69 ( .A(n812), .Y(n884) );
  NAND2X1 U71 ( .A(n531), .B(n852), .Y(n693) );
  NAND2X1 U72 ( .A(n531), .B(n857), .Y(n586) );
  NAND2BX1 U73 ( .AN(n799), .B(n660), .Y(n727) );
  INVX1 U74 ( .A(n767), .Y(n899) );
  NAND2X1 U75 ( .A(n699), .B(n655), .Y(n782) );
  NAND2BX1 U76 ( .AN(n830), .B(n537), .Y(n624) );
  NAND2X1 U77 ( .A(n699), .B(n690), .Y(n819) );
  NAND2X1 U78 ( .A(n660), .B(n781), .Y(n823) );
  CLKINVX3 U79 ( .A(n534), .Y(n902) );
  CLKINVX3 U80 ( .A(n815), .Y(n901) );
  INVX1 U81 ( .A(n674), .Y(d[3]) );
  BUFX3 U82 ( .A(a[1]), .Y(n531) );
  NAND2X1 U83 ( .A(a[7]), .B(a[2]), .Y(n829) );
  NAND2X1 U84 ( .A(n533), .B(a[0]), .Y(n815) );
  INVX1 U85 ( .A(n685), .Y(n907) );
  NAND2X1 U86 ( .A(n864), .B(n540), .Y(n809) );
  NAND2X1 U87 ( .A(n872), .B(n556), .Y(n685) );
  INVX1 U88 ( .A(n635), .Y(n908) );
  NOR2X1 U89 ( .A(n550), .B(n598), .Y(n724) );
  NOR2X1 U90 ( .A(n874), .B(n861), .Y(n676) );
  NAND2X1 U91 ( .A(n701), .B(n540), .Y(n761) );
  INVX1 U92 ( .A(n622), .Y(n874) );
  INVX1 U93 ( .A(n675), .Y(n886) );
  INVX1 U94 ( .A(n757), .Y(n863) );
  INVX1 U95 ( .A(n716), .Y(n875) );
  INVX1 U96 ( .A(n695), .Y(n872) );
  INVX4 U97 ( .A(n536), .Y(n556) );
  NOR2BX1 U98 ( .AN(n709), .B(n854), .Y(n835) );
  NOR2X1 U99 ( .A(n870), .B(n853), .Y(n597) );
  AOI22X1 U100 ( .A0(n900), .A1(n788), .B0(n898), .B1(n787), .Y(n789) );
  OAI221XL U101 ( .A0(n887), .A1(n550), .B0(n802), .B1(n543), .C0(n783), .Y(
        n788) );
  INVX1 U102 ( .A(n838), .Y(n887) );
  NOR2X1 U104 ( .A(n873), .B(n862), .Y(n637) );
  NAND2X1 U105 ( .A(n889), .B(n700), .Y(n740) );
  INVX1 U106 ( .A(n805), .Y(n853) );
  NAND2X1 U107 ( .A(n889), .B(n675), .Y(n800) );
  INVX1 U108 ( .A(n690), .Y(n868) );
  INVX1 U109 ( .A(n700), .Y(n864) );
  NOR2X1 U110 ( .A(n866), .B(n868), .Y(n726) );
  OAI221XL U111 ( .A0(n865), .A1(n545), .B0(n825), .B1(n829), .C0(n905), .Y(
        n576) );
  INVX1 U112 ( .A(n724), .Y(n905) );
  INVX1 U113 ( .A(n796), .Y(n888) );
  NOR2X1 U114 ( .A(n864), .B(n854), .Y(n825) );
  INVX1 U115 ( .A(n711), .Y(n882) );
  INVX1 U116 ( .A(n617), .Y(n865) );
  INVX1 U117 ( .A(n765), .Y(n881) );
  INVX1 U118 ( .A(n836), .Y(n885) );
  INVX1 U119 ( .A(n713), .Y(n879) );
  NAND2X1 U120 ( .A(n860), .B(n535), .Y(n680) );
  OAI22X1 U121 ( .A0(n683), .A1(n813), .B0(n682), .B1(n769), .Y(n687) );
  AOI222X1 U122 ( .A0(n862), .A1(n548), .B0(n556), .B1(n679), .C0(n678), .C1(
        n711), .Y(n683) );
  AOI211X1 U123 ( .A0(n556), .A1(n689), .B0(n681), .C0(n724), .Y(n682) );
  NAND2X1 U124 ( .A(n807), .B(n694), .Y(n679) );
  NOR2X1 U125 ( .A(n877), .B(n866), .Y(n701) );
  OAI22X1 U126 ( .A0(n829), .A1(n716), .B0(n545), .B1(n538), .Y(n681) );
  CLKINVX3 U127 ( .A(n810), .Y(n873) );
  CLKINVX3 U128 ( .A(n742), .Y(n860) );
  AOI22X1 U129 ( .A0(n899), .A1(n832), .B0(n900), .B1(n831), .Y(n845) );
  OAI221XL U130 ( .A0(n825), .A1(n545), .B0(n893), .B1(n543), .C0(n824), .Y(
        n832) );
  OAI221XL U131 ( .A0(n881), .A1(n545), .B0(n872), .B1(n543), .C0(n828), .Y(
        n831) );
  INVX1 U132 ( .A(n819), .Y(n893) );
  NAND2X1 U133 ( .A(n556), .B(n827), .Y(n736) );
  NAND2X1 U134 ( .A(n808), .B(n709), .Y(n695) );
  AOI22X1 U135 ( .A0(n900), .A1(n729), .B0(n901), .B1(n728), .Y(n730) );
  OAI221XL U136 ( .A0(n536), .A1(n727), .B0(n726), .B1(n545), .C0(n725), .Y(
        n728) );
  AOI211X1 U137 ( .A0(n722), .A1(n556), .B0(n721), .C0(n720), .Y(n723) );
  AOI22X1 U138 ( .A0(n900), .A1(n592), .B0(n901), .B1(n591), .Y(n593) );
  OAI221XL U139 ( .A0(n888), .A1(n545), .B0(n879), .B1(n543), .C0(n590), .Y(
        n591) );
  OAI211X1 U140 ( .A0(n597), .A1(n550), .B0(n635), .C0(n589), .Y(n592) );
  AOI22X1 U141 ( .A0(n888), .A1(n556), .B0(n884), .B1(n552), .Y(n590) );
  AOI22X1 U142 ( .A0(n548), .A1(n860), .B0(n676), .B1(n539), .Y(n589) );
  AOI21X1 U143 ( .A0(n808), .A1(n680), .B0(n550), .Y(n563) );
  INVX1 U144 ( .A(n803), .Y(n916) );
  AND2X2 U145 ( .A(n758), .B(n757), .Y(n794) );
  OAI21XL U146 ( .A0(n758), .A1(n550), .B0(n736), .Y(n657) );
  INVX1 U147 ( .A(n639), .Y(n911) );
  OAI31X1 U148 ( .A0(n721), .A1(n908), .A2(n638), .B0(n898), .Y(n639) );
  OAI21XL U149 ( .A0(n541), .A1(n637), .B0(n636), .Y(n638) );
  INVX1 U150 ( .A(n776), .Y(n876) );
  OAI22X1 U152 ( .A0(n621), .A1(n769), .B0(n620), .B1(n813), .Y(n626) );
  AOI211X1 U153 ( .A0(n556), .A1(n821), .B0(n619), .C0(n618), .Y(n620) );
  AOI221X1 U154 ( .A0(n910), .A1(n535), .B0(n896), .B1(n556), .C0(n616), .Y(
        n621) );
  OAI22X1 U155 ( .A0(n859), .A1(n543), .B0(n550), .B1(n617), .Y(n619) );
  AOI222X1 U156 ( .A0(n867), .A1(n540), .B0(n863), .B1(n554), .C0(n547), .C1(
        n852), .Y(n567) );
  AOI21X1 U157 ( .A0(n873), .A1(n556), .B0(n557), .Y(n558) );
  AOI2BB2X1 U158 ( .B0(n910), .B1(n535), .A0N(n536), .A1N(n676), .Y(n677) );
  CLKINVX8 U159 ( .A(n546), .Y(n545) );
  CLKINVX3 U160 ( .A(n541), .Y(n539) );
  NOR2X1 U161 ( .A(n545), .B(n535), .Y(n721) );
  AOI222X1 U162 ( .A0(n916), .A1(n810), .B0(n724), .B1(n873), .C0(n886), .C1(
        n540), .Y(n725) );
  AOI221X1 U163 ( .A0(n602), .A1(n553), .B0(n540), .B1(n612), .C0(n596), .Y(
        n608) );
  OAI221XL U164 ( .A0(n536), .A1(n714), .B0(n545), .B1(n820), .C0(n635), .Y(
        n596) );
  AOI221X1 U165 ( .A0(n916), .A1(n852), .B0(n553), .B1(n810), .C0(n737), .Y(
        n749) );
  OAI2BB1X1 U167 ( .A0N(n781), .A1N(n548), .B0(n736), .Y(n737) );
  NOR2X1 U168 ( .A(n854), .B(n855), .Y(n615) );
  OAI221XL U169 ( .A0(n869), .A1(n545), .B0(n890), .B1(n543), .C0(n691), .Y(
        n706) );
  INVX1 U170 ( .A(n689), .Y(n869) );
  AOI32X1 U171 ( .A0(n889), .A1(n742), .A2(n556), .B0(n553), .B1(n690), .Y(
        n691) );
  INVX1 U172 ( .A(n808), .Y(n856) );
  AOI211X1 U173 ( .A0(n875), .A1(n556), .B0(n914), .C0(n628), .Y(n629) );
  INVX1 U174 ( .A(n809), .Y(n914) );
  AOI211X1 U175 ( .A0(n863), .A1(n540), .B0(n909), .C0(n559), .Y(n560) );
  NOR3X1 U176 ( .A(n545), .B(n884), .C(n862), .Y(n559) );
  INVX1 U177 ( .A(n664), .Y(n909) );
  OAI221XL U178 ( .A0(n536), .A1(n755), .B0(n759), .B1(n551), .C0(n754), .Y(
        n773) );
  AOI22X1 U179 ( .A0(n549), .A1(n889), .B0(n875), .B1(n539), .Y(n754) );
  AOI211X1 U180 ( .A0(n554), .A1(n827), .B0(n908), .C0(n826), .Y(n828) );
  AOI211X1 U181 ( .A0(n878), .A1(n540), .B0(n719), .C0(n718), .Y(n731) );
  INVX1 U182 ( .A(n714), .Y(n878) );
  NAND2BX1 U183 ( .AN(n826), .B(n717), .Y(n718) );
  OAI222X1 U184 ( .A0(n551), .A1(n716), .B0(n742), .B1(n803), .C0(n545), .C1(
        n715), .Y(n719) );
  CLKINVX3 U185 ( .A(n555), .Y(n551) );
  INVX1 U186 ( .A(n798), .Y(n913) );
  AOI221X1 U187 ( .A0(n797), .A1(n552), .B0(n796), .B1(n549), .C0(n795), .Y(
        n798) );
  OAI21XL U188 ( .A0(n536), .A1(n794), .B0(n793), .Y(n795) );
  INVX1 U189 ( .A(n536), .Y(n906) );
  NOR2X1 U190 ( .A(n884), .B(n866), .Y(n744) );
  NAND3X1 U191 ( .A(n538), .B(n810), .C(n540), .Y(n834) );
  NAND2X1 U192 ( .A(n709), .B(n781), .Y(n833) );
  NAND2X1 U193 ( .A(n807), .B(n781), .Y(n838) );
  NAND2X1 U194 ( .A(n808), .B(n655), .Y(n765) );
  NAND2X1 U195 ( .A(n538), .B(n757), .Y(n612) );
  NOR2BX1 U196 ( .AN(n694), .B(n855), .Y(n759) );
  AOI21X1 U197 ( .A0(n742), .A1(n741), .B0(n536), .Y(n743) );
  AOI22X1 U198 ( .A0(n874), .A1(n548), .B0(n556), .B1(n782), .Y(n783) );
  AOI22X1 U199 ( .A0(n866), .A1(n546), .B0(n555), .B1(n810), .Y(n684) );
  AOI22X1 U200 ( .A0(n547), .A1(n612), .B0(n873), .B1(n539), .Y(n573) );
  NOR2X1 U201 ( .A(n785), .B(n536), .Y(n826) );
  NAND2X1 U202 ( .A(n680), .B(n781), .Y(n796) );
  INVX1 U203 ( .A(n769), .Y(n898) );
  NAND2X1 U204 ( .A(n694), .B(n680), .Y(n689) );
  CLKINVX3 U205 ( .A(n785), .Y(n867) );
  NAND2X1 U206 ( .A(n694), .B(n714), .Y(n663) );
  NOR2X1 U207 ( .A(n859), .B(n799), .Y(n802) );
  AOI211X1 U208 ( .A0(n556), .A1(n617), .B0(n588), .C0(n587), .Y(n594) );
  OAI2BB2X1 U209 ( .B0(n545), .B1(n740), .A0N(n735), .A1N(n540), .Y(n588) );
  AOI21X1 U210 ( .A0(n622), .A1(n586), .B0(n550), .Y(n587) );
  NAND2X1 U211 ( .A(n538), .B(n709), .Y(n797) );
  NAND2X1 U212 ( .A(n785), .B(n821), .Y(n696) );
  NAND2X1 U213 ( .A(n820), .B(n758), .Y(n735) );
  AOI21X1 U214 ( .A0(n556), .A1(n823), .B0(n822), .Y(n824) );
  AOI21X1 U215 ( .A0(n821), .A1(n820), .B0(n550), .Y(n822) );
  OAI221XL U216 ( .A0(n858), .A1(n551), .B0(n892), .B1(n536), .C0(n774), .Y(
        n780) );
  AOI2BB2X1 U217 ( .B0(n539), .B1(n836), .A0N(n545), .A1N(n802), .Y(n774) );
  INVX1 U218 ( .A(n586), .Y(n858) );
  INVX1 U219 ( .A(n715), .Y(n894) );
  INVX1 U220 ( .A(n624), .Y(n910) );
  INVX1 U221 ( .A(n823), .Y(n890) );
  AOI221XL U222 ( .A0(n556), .A1(n871), .B0(n548), .B1(n800), .C0(n599), .Y(
        n607) );
  INVX1 U223 ( .A(n597), .Y(n871) );
  OAI32X1 U224 ( .A0(n542), .A1(n860), .A2(n598), .B0(n886), .B1(n551), .Y(
        n599) );
  INVX1 U225 ( .A(n727), .Y(n892) );
  OAI221XL U226 ( .A0(n867), .A1(n545), .B0(n891), .B1(n542), .C0(n760), .Y(
        n772) );
  INVX1 U227 ( .A(n756), .Y(n891) );
  AOI22X1 U228 ( .A0(n759), .A1(n556), .B0(n794), .B1(n552), .Y(n760) );
  INVX1 U229 ( .A(n782), .Y(n896) );
  INVX1 U230 ( .A(n827), .Y(n883) );
  AOI31X1 U231 ( .A0(n821), .A1(n785), .A2(n556), .B0(n912), .Y(n786) );
  INVX1 U232 ( .A(n834), .Y(n912) );
  INVX1 U233 ( .A(n738), .Y(n904) );
  INVX1 U234 ( .A(n540), .Y(n542) );
  INVX1 U235 ( .A(n540), .Y(n543) );
  AOI211X1 U236 ( .A0(n901), .A1(n627), .B0(n626), .C0(n625), .Y(n643) );
  AOI211X1 U237 ( .A0(n901), .A1(n641), .B0(n640), .C0(n911), .Y(n642) );
  OAI2BB2X1 U238 ( .B0(n614), .B1(n613), .A0N(n744), .A1N(n614), .Y(n627) );
  AOI211X1 U239 ( .A0(n901), .A1(n688), .B0(n687), .C0(n686), .Y(n708) );
  AOI211X1 U240 ( .A0(n900), .A1(n706), .B0(n705), .C0(n704), .Y(n707) );
  AOI31X1 U241 ( .A0(n685), .A1(n793), .A2(n684), .B0(n767), .Y(n686) );
  OAI21X2 U242 ( .A0(n534), .A1(n792), .B0(n791), .Y(d[6]) );
  OAI2BB1X1 U243 ( .A0N(n790), .A1N(n789), .B0(n534), .Y(n791) );
  AOI221X1 U244 ( .A0(n900), .A1(n773), .B0(n901), .B1(n772), .C0(n771), .Y(
        n792) );
  AOI22X1 U245 ( .A0(n899), .A1(n780), .B0(n901), .B1(n779), .Y(n790) );
  OAI2BB1X1 U246 ( .A0N(n845), .A1N(n844), .B0(n902), .Y(n846) );
  AOI22X1 U247 ( .A0(n901), .A1(n843), .B0(n898), .B1(n842), .Y(n844) );
  AOI22X1 U248 ( .A0(n533), .A1(n669), .B0(n668), .B1(n897), .Y(n670) );
  OAI221XL U249 ( .A0(n862), .A1(n551), .B0(n545), .B1(n663), .C0(n662), .Y(
        n669) );
  OAI221XL U250 ( .A0(n882), .A1(n545), .B0(n543), .B1(n742), .C0(n667), .Y(
        n668) );
  AOI21X1 U251 ( .A0(n890), .A1(n906), .B0(n661), .Y(n662) );
  AOI22X1 U252 ( .A0(n575), .A1(n897), .B0(n533), .B1(n574), .Y(n581) );
  OAI221XL U253 ( .A0(n536), .A1(n757), .B0(n637), .B1(n545), .C0(n572), .Y(
        n575) );
  OAI211X1 U254 ( .A0(n835), .A1(n550), .B0(n736), .C0(n573), .Y(n574) );
  AOI2BB2X1 U255 ( .B0(n539), .B1(n727), .A0N(n550), .A1N(n744), .Y(n572) );
  OAI22X1 U256 ( .A0(n634), .A1(n813), .B0(n633), .B1(n767), .Y(n640) );
  AOI221XL U257 ( .A0(n549), .A1(n740), .B0(n799), .B1(n850), .C0(n632), .Y(
        n633) );
  AOI221XL U258 ( .A0(n867), .A1(n916), .B0(n547), .B1(n713), .C0(n630), .Y(
        n634) );
  OAI32X1 U259 ( .A0(n738), .A1(n860), .A2(n850), .B0(n631), .B1(n904), .Y(
        n632) );
  OAI22X1 U260 ( .A0(n770), .A1(n769), .B0(n768), .B1(n767), .Y(n771) );
  AOI211X1 U261 ( .A0(n881), .A1(n850), .B0(n766), .C0(n907), .Y(n768) );
  AOI221XL U262 ( .A0(n862), .A1(n554), .B0(n547), .B1(n776), .C0(n764), .Y(
        n770) );
  OAI22X1 U263 ( .A0(n542), .A1(n852), .B0(n886), .B1(n550), .Y(n766) );
  OAI22X1 U264 ( .A0(n816), .A1(n815), .B0(n814), .B1(n813), .Y(n817) );
  AOI221XL U265 ( .A0(n549), .A1(n812), .B0(n876), .B1(n540), .C0(n811), .Y(
        n814) );
  AOI221X1 U266 ( .A0(n556), .A1(n808), .B0(n553), .B1(n807), .C0(n806), .Y(
        n816) );
  OAI221XL U267 ( .A0(n536), .A1(n810), .B0(n879), .B1(n551), .C0(n809), .Y(
        n811) );
  AOI211X1 U268 ( .A0(n868), .A1(n556), .B0(n652), .C0(n651), .Y(n653) );
  AOI31X1 U269 ( .A0(n809), .A1(n717), .A2(n650), .B0(n533), .Y(n651) );
  OAI22X1 U270 ( .A0(n857), .A1(n803), .B0(n649), .B1(n897), .Y(n652) );
  AOI2BB2X1 U271 ( .B0(n853), .B1(n554), .A0N(n833), .A1N(n545), .Y(n650) );
  AOI2BB2X1 U272 ( .B0(n659), .B1(n897), .A0N(n897), .A1N(n658), .Y(n671) );
  OAI221XL U273 ( .A0(n877), .A1(n551), .B0(n545), .B1(n807), .C0(n656), .Y(
        n659) );
  AOI221XL U274 ( .A0(n548), .A1(n676), .B0(n711), .B1(n540), .C0(n657), .Y(
        n658) );
  AOI22X1 U275 ( .A0(n539), .A1(n765), .B0(n873), .B1(n903), .Y(n656) );
  AOI22X1 U276 ( .A0(n554), .A1(n532), .B0(n539), .B1(n857), .Y(n631) );
  AOI22X1 U277 ( .A0(n900), .A1(n747), .B0(n899), .B1(n746), .Y(n748) );
  OAI221XL U278 ( .A0(n860), .A1(n545), .B0(n542), .B1(n807), .C0(n745), .Y(
        n746) );
  OAI221XL U279 ( .A0(n885), .A1(n536), .B0(n545), .B1(n740), .C0(n739), .Y(
        n747) );
  AOI21X1 U281 ( .A0(n744), .A1(n552), .B0(n743), .Y(n745) );
  AOI22X1 U282 ( .A0(n533), .A1(n562), .B0(n561), .B1(n897), .Y(n571) );
  OAI221XL U283 ( .A0(n880), .A1(n545), .B0(n541), .B1(n889), .C0(n558), .Y(
        n562) );
  OAI221XL U284 ( .A0(n532), .A1(n803), .B0(n722), .B1(n551), .C0(n560), .Y(
        n561) );
  INVX1 U285 ( .A(n663), .Y(n880) );
  AOI22X1 U286 ( .A0(n901), .A1(n605), .B0(n900), .B1(n604), .Y(n606) );
  OAI21XL U287 ( .A0(n602), .A1(n536), .B0(n601), .Y(n605) );
  OAI221XL U288 ( .A0(n551), .A1(n810), .B0(n835), .B1(n545), .C0(n603), .Y(
        n604) );
  AOI31X1 U289 ( .A0(n538), .A1(n742), .A2(n600), .B0(n910), .Y(n601) );
  INVX1 U290 ( .A(n611), .Y(d[1]) );
  AOI22X1 U291 ( .A0(n534), .A1(n610), .B0(n609), .B1(n902), .Y(n611) );
  OAI221XL U292 ( .A0(n595), .A1(n767), .B0(n594), .B1(n769), .C0(n593), .Y(
        n610) );
  OAI221XL U293 ( .A0(n608), .A1(n767), .B0(n607), .B1(n769), .C0(n606), .Y(
        n609) );
  INVX1 U294 ( .A(n753), .Y(d[5]) );
  AOI22X1 U295 ( .A0(n752), .A1(n902), .B0(n534), .B1(n751), .Y(n753) );
  OAI221XL U296 ( .A0(n750), .A1(n815), .B0(n749), .B1(n769), .C0(n748), .Y(
        n751) );
  OAI221XL U297 ( .A0(n732), .A1(n769), .B0(n731), .B1(n767), .C0(n730), .Y(
        n752) );
  CLKINVX3 U298 ( .A(n532), .Y(n852) );
  OAI21XL U299 ( .A0(n545), .A1(n537), .B0(n803), .Y(n647) );
  NAND2X1 U300 ( .A(n860), .B(n531), .Y(n755) );
  AOI21X1 U301 ( .A0(n699), .A1(n680), .B0(n545), .Y(n628) );
  INVX1 U302 ( .A(n531), .Y(n849) );
  OAI21XL U303 ( .A0(n850), .A1(n622), .B0(n550), .Y(n600) );
  OAI21XL U304 ( .A0(n536), .A1(n805), .B0(n763), .Y(n764) );
  AOI31X1 U305 ( .A0(n812), .A1(n903), .A2(n762), .B0(n915), .Y(n763) );
  INVX1 U306 ( .A(n761), .Y(n915) );
  AOI211X1 U307 ( .A0(n884), .A1(n540), .B0(n648), .C0(n647), .Y(n649) );
  OAI222X1 U308 ( .A0(n551), .A1(n807), .B0(n850), .B1(n693), .C0(n545), .C1(
        n821), .Y(n648) );
  NAND2X1 U309 ( .A(n861), .B(n552), .Y(n636) );
  NOR2BX1 U310 ( .AN(n660), .B(n876), .Y(n722) );
  BUFX3 U311 ( .A(n841), .Y(n536) );
  NAND2X1 U312 ( .A(n850), .B(n903), .Y(n841) );
  OAI221XL U313 ( .A0(n531), .A1(n664), .B0(n829), .B1(n709), .C0(n636), .Y(
        n630) );
  BUFX3 U314 ( .A(n784), .Y(n538) );
  NAND2X1 U315 ( .A(n531), .B(n537), .Y(n784) );
  AOI211X1 U316 ( .A0(n540), .A1(n852), .B0(n585), .C0(n647), .Y(n595) );
  OAI222X1 U317 ( .A0(n551), .A1(n756), .B0(n584), .B1(n536), .C0(n545), .C1(
        n889), .Y(n585) );
  AOI21X1 U318 ( .A0(n537), .A1(n535), .B0(n858), .Y(n584) );
  AOI211X1 U319 ( .A0(n533), .A1(n569), .B0(n848), .C0(n568), .Y(n570) );
  OAI221XL U320 ( .A0(n545), .A1(n807), .B0(n602), .B1(n829), .C0(n564), .Y(
        n569) );
  AOI21X1 U321 ( .A0(n567), .A1(n566), .B0(n533), .Y(n568) );
  AOI31X1 U322 ( .A0(n556), .A1(n565), .A2(n884), .B0(n563), .Y(n564) );
  INVX1 U323 ( .A(n830), .Y(n546) );
  INVX1 U324 ( .A(n840), .Y(n554) );
  INVX1 U325 ( .A(n840), .Y(n555) );
  INVX1 U326 ( .A(n544), .Y(n541) );
  INVX1 U327 ( .A(n829), .Y(n544) );
  AOI22X1 U328 ( .A0(n533), .A1(n646), .B0(n645), .B1(n897), .Y(n654) );
  OAI222X1 U329 ( .A0(n545), .A1(n782), .B0(n551), .B1(n660), .C0(n894), .C1(
        n542), .Y(n646) );
  OAI221XL U330 ( .A0(n892), .A1(n536), .B0(n551), .B1(n819), .C0(n644), .Y(
        n645) );
  AOI2BB2X1 U331 ( .B0(n835), .B1(n539), .A0N(n545), .A1N(n726), .Y(n644) );
  NAND2X1 U332 ( .A(n699), .B(n622), .Y(n775) );
  NOR2BX1 U333 ( .AN(n660), .B(n862), .Y(n602) );
  AOI21X1 U334 ( .A0(n690), .A1(n758), .B0(n903), .Y(n661) );
  AOI22X1 U335 ( .A0(n549), .A1(n838), .B0(n882), .B1(n539), .Y(n839) );
  AOI31X1 U336 ( .A0(n703), .A1(n793), .A2(n702), .B0(n815), .Y(n704) );
  OAI2BB1X1 U337 ( .A0N(n700), .A1N(n699), .B0(n553), .Y(n703) );
  AOI22X1 U338 ( .A0(n894), .A1(n556), .B0(n701), .B1(n547), .Y(n702) );
  NAND2X1 U339 ( .A(n699), .B(n805), .Y(n715) );
  NAND2X1 U340 ( .A(n660), .B(n586), .Y(n756) );
  AOI21X1 U341 ( .A0(n660), .A1(n741), .B0(n545), .Y(n618) );
  AOI21X1 U342 ( .A0(n812), .A1(n538), .B0(n829), .Y(n720) );
  NAND2X1 U343 ( .A(n906), .B(n531), .Y(n717) );
  OAI21XL U344 ( .A0(n850), .A1(n680), .B0(n550), .Y(n678) );
  XNOR2X1 U345 ( .A(n903), .B(n531), .Y(n738) );
  NAND2X1 U346 ( .A(n539), .B(n537), .Y(n793) );
  XNOR2X1 U347 ( .A(n850), .B(n531), .Y(n762) );
  AOI21X1 U348 ( .A0(n833), .A1(n850), .B0(n556), .Y(n837) );
  AOI221X1 U349 ( .A0(n877), .A1(n540), .B0(n552), .B1(n735), .C0(n734), .Y(
        n750) );
  AOI21X1 U350 ( .A0(n536), .A1(n733), .B0(n799), .Y(n734) );
  OAI21XL U351 ( .A0(n861), .A1(n853), .B0(n850), .Y(n733) );
  AOI222X1 U352 ( .A0(n549), .A1(n713), .B0(n712), .B1(n711), .C0(n556), .C1(
        n537), .Y(n732) );
  OAI21XL U353 ( .A0(n850), .A1(n709), .B0(n550), .Y(n712) );
  NOR2X1 U354 ( .A(n861), .B(n868), .Y(n778) );
  AOI22X1 U355 ( .A0(n906), .A1(n857), .B0(n539), .B1(n776), .Y(n777) );
  INVX1 U356 ( .A(n775), .Y(n895) );
  AOI31X1 U357 ( .A0(n761), .A1(n624), .A2(n623), .B0(n767), .Y(n625) );
  AOI22X1 U358 ( .A0(n775), .A1(n850), .B0(n894), .B1(n553), .Y(n623) );
  INVX1 U359 ( .A(n830), .Y(n547) );
  INVX1 U360 ( .A(n830), .Y(n549) );
  INVX1 U361 ( .A(n830), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n565) );
  INVX1 U363 ( .A(n840), .Y(n552) );
  INVX1 U364 ( .A(n840), .Y(n553) );
  NOR2BX1 U365 ( .AN(n830), .B(n554), .Y(n614) );
  OAI22X2 U366 ( .A0(n583), .A1(n902), .B0(n534), .B1(n582), .Y(d[0]) );
  AOI22X1 U367 ( .A0(n581), .A1(a[0]), .B0(n580), .B1(n579), .Y(n582) );
  AOI31X1 U368 ( .A0(n717), .A1(n848), .A2(n571), .B0(n570), .Y(n583) );
  AOI22X1 U369 ( .A0(n576), .A1(n897), .B0(n556), .B1(n833), .Y(n580) );
  AOI22X1 U370 ( .A0(n673), .A1(n902), .B0(n534), .B1(n672), .Y(n674) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n654), .B0(n653), .B1(n848), .Y(n673) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n671), .B0(n670), .B1(n848), .Y(n672) );
  OAI22X1 U373 ( .A0(n698), .A1(n767), .B0(n697), .B1(n769), .Y(n705) );
  AOI221X1 U374 ( .A0(n548), .A1(n693), .B0(n556), .B1(n797), .C0(n692), .Y(
        n698) );
  AOI222X1 U375 ( .A0(n759), .A1(n547), .B0(a[2]), .B1(n696), .C0(n556), .C1(
        n695), .Y(n697) );
  OAI22X1 U376 ( .A0(n888), .A1(n543), .B0(n550), .B1(n537), .Y(n692) );
  NOR2X1 U377 ( .A(n863), .B(n861), .Y(n804) );
  BUFX3 U378 ( .A(n710), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n852), .Y(n710) );
  AOI221X1 U380 ( .A0(n916), .A1(n785), .B0(n851), .B1(n666), .C0(n665), .Y(
        n667) );
  NOR3X1 U381 ( .A(n851), .B(a[7]), .C(n860), .Y(n665) );
  INVX1 U382 ( .A(n762), .Y(n851) );
  OAI21XL U383 ( .A0(n857), .A1(n550), .B0(n664), .Y(n666) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI33X1 U385 ( .A0(n532), .A1(n540), .A2(n904), .B0(n738), .B1(n742), .B2(
        a[2]), .Y(n739) );
  AOI22X1 U386 ( .A0(n882), .A1(n850), .B0(a[2]), .B1(n612), .Y(n613) );
  CLKINVX3 U387 ( .A(a[0]), .Y(n848) );
  AOI211X1 U388 ( .A0(n724), .A1(n578), .B0(n577), .C0(a[0]), .Y(n579) );
  NAND2X1 U389 ( .A(n781), .B(n805), .Y(n578) );
  AOI21X1 U390 ( .A0(n803), .A1(n624), .B0(n897), .Y(n577) );
  BUFX3 U391 ( .A(a[5]), .Y(n533) );
  OAI221XL U392 ( .A0(n536), .A1(n808), .B0(n802), .B1(n545), .C0(n801), .Y(
        n818) );
  AOI22X1 U393 ( .A0(n539), .A1(n800), .B0(n799), .B1(a[2]), .Y(n801) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_14 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916;

  OAI221X4 U4 ( .A0(n857), .A1(n536), .B0(n862), .B1(n551), .C0(n839), .Y(n842) );
  OAI221X4 U6 ( .A0(n837), .A1(n836), .B0(n835), .B1(n551), .C0(n834), .Y(n843) );
  OAI222X4 U75 ( .A0(n551), .A1(n716), .B0(n742), .B1(n803), .C0(n545), .C1(
        n715), .Y(n719) );
  OAI32X4 U280 ( .A0(n551), .A1(n867), .A2(n870), .B0(n829), .B1(n820), .Y(
        n557) );
  AOI221X1 U1 ( .A0(n858), .A1(a[2]), .B0(n826), .B1(n565), .C0(n916), .Y(n566) );
  INVX1 U2 ( .A(a[7]), .Y(n903) );
  NAND2X1 U3 ( .A(n532), .B(n535), .Y(n820) );
  OAI222X1 U5 ( .A0(n829), .A1(n805), .B0(n804), .B1(n545), .C0(a[4]), .C1(
        n803), .Y(n806) );
  NAND2X2 U7 ( .A(n531), .B(n532), .Y(n808) );
  NAND2X1 U8 ( .A(n867), .B(n531), .Y(n694) );
  NAND2X2 U9 ( .A(n532), .B(n857), .Y(n742) );
  NAND2X1 U10 ( .A(n884), .B(n531), .Y(n781) );
  NAND2X2 U11 ( .A(n537), .B(n742), .Y(n810) );
  NAND2X2 U12 ( .A(n857), .B(n535), .Y(n807) );
  NAND2X2 U13 ( .A(n857), .B(n852), .Y(n785) );
  NAND2X1 U14 ( .A(n531), .B(n742), .Y(n821) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n850) );
  NAND2X1 U16 ( .A(n533), .B(n848), .Y(n813) );
  CLKINVX3 U17 ( .A(n533), .Y(n897) );
  NAND2X2 U18 ( .A(n848), .B(n897), .Y(n769) );
  NAND2X2 U19 ( .A(a[0]), .B(n897), .Y(n767) );
  CLKINVX3 U20 ( .A(n534), .Y(n902) );
  OAI22X2 U21 ( .A0(n583), .A1(n902), .B0(n534), .B1(n582), .Y(d[0]) );
  OAI22X2 U22 ( .A0(n534), .A1(n643), .B0(n642), .B1(n902), .Y(d[2]) );
  INVX1 U23 ( .A(n674), .Y(d[3]) );
  OAI21X2 U24 ( .A0(n847), .A1(n902), .B0(n846), .Y(d[7]) );
  AOI221X1 U25 ( .A0(n899), .A1(n913), .B0(n898), .B1(n818), .C0(n817), .Y(
        n847) );
  OAI22X2 U26 ( .A0(n534), .A1(n708), .B0(n707), .B1(n902), .Y(d[4]) );
  OAI21X2 U27 ( .A0(n534), .A1(n792), .B0(n791), .Y(d[6]) );
  AOI221X1 U28 ( .A0(n900), .A1(n773), .B0(n901), .B1(n772), .C0(n771), .Y(
        n792) );
  NAND2X1 U29 ( .A(a[2]), .B(n903), .Y(n840) );
  NAND2X1 U30 ( .A(a[7]), .B(n850), .Y(n830) );
  AOI21XL U31 ( .A0(n916), .A1(a[4]), .B0(n907), .Y(n603) );
  NAND2X1 U32 ( .A(a[4]), .B(n535), .Y(n660) );
  NAND2X1 U33 ( .A(n531), .B(a[4]), .Y(n699) );
  NAND2X2 U34 ( .A(n532), .B(a[4]), .Y(n812) );
  CLKINVX3 U35 ( .A(a[4]), .Y(n857) );
  NAND2X1 U36 ( .A(n870), .B(n906), .Y(n635) );
  CLKINVX3 U37 ( .A(n542), .Y(n540) );
  INVX1 U38 ( .A(n598), .Y(n889) );
  NAND2X1 U39 ( .A(n810), .B(n535), .Y(n709) );
  NAND2X1 U40 ( .A(n867), .B(n535), .Y(n690) );
  NAND2X1 U41 ( .A(n877), .B(n535), .Y(n714) );
  NAND2X1 U42 ( .A(n873), .B(n535), .Y(n622) );
  NAND2X1 U43 ( .A(n538), .B(n655), .Y(n711) );
  NAND2X1 U44 ( .A(n776), .B(n709), .Y(n716) );
  NAND2X1 U45 ( .A(n808), .B(n714), .Y(n713) );
  INVX1 U46 ( .A(n755), .Y(n861) );
  INVX1 U47 ( .A(n538), .Y(n870) );
  INVX1 U48 ( .A(n741), .Y(n866) );
  NOR2X1 U49 ( .A(n535), .B(n884), .Y(n598) );
  CLKINVX3 U50 ( .A(n555), .Y(n550) );
  NAND2X1 U51 ( .A(n535), .B(n852), .Y(n805) );
  NAND2X1 U52 ( .A(n785), .B(n535), .Y(n700) );
  NAND2X1 U53 ( .A(n884), .B(n535), .Y(n675) );
  NAND2X1 U54 ( .A(n742), .B(n535), .Y(n757) );
  NAND2X1 U55 ( .A(n694), .B(n675), .Y(n836) );
  INVX1 U56 ( .A(n821), .Y(n862) );
  NAND2X1 U57 ( .A(n808), .B(n700), .Y(n617) );
  INVX1 U58 ( .A(n693), .Y(n854) );
  INVX1 U59 ( .A(n807), .Y(n859) );
  INVX1 U60 ( .A(n820), .Y(n855) );
  BUFX3 U61 ( .A(n849), .Y(n535) );
  NAND2X1 U62 ( .A(n873), .B(n531), .Y(n776) );
  NAND2X1 U63 ( .A(n531), .B(n539), .Y(n803) );
  NAND2X1 U64 ( .A(n812), .B(n535), .Y(n655) );
  NAND2X1 U65 ( .A(n531), .B(n810), .Y(n758) );
  NAND2X1 U66 ( .A(n531), .B(n785), .Y(n741) );
  INVX1 U67 ( .A(n611), .Y(d[1]) );
  INVX1 U68 ( .A(n753), .Y(d[5]) );
  INVX1 U69 ( .A(n537), .Y(n877) );
  NAND2X1 U70 ( .A(n906), .B(n532), .Y(n664) );
  NAND2X1 U71 ( .A(n812), .B(n776), .Y(n827) );
  NOR2X1 U72 ( .A(n537), .B(n535), .Y(n799) );
  CLKINVX3 U73 ( .A(n812), .Y(n884) );
  NAND2X1 U74 ( .A(n531), .B(n852), .Y(n693) );
  NAND2X1 U76 ( .A(n531), .B(n857), .Y(n586) );
  NAND2BX1 U77 ( .AN(n799), .B(n660), .Y(n727) );
  INVX1 U78 ( .A(n767), .Y(n899) );
  NAND2X1 U79 ( .A(n699), .B(n655), .Y(n782) );
  NAND2BX1 U80 ( .AN(n830), .B(n537), .Y(n624) );
  NAND2X1 U81 ( .A(n699), .B(n690), .Y(n819) );
  NAND2X1 U82 ( .A(n660), .B(n781), .Y(n823) );
  CLKINVX3 U83 ( .A(n815), .Y(n901) );
  BUFX3 U84 ( .A(a[1]), .Y(n531) );
  NAND2X1 U85 ( .A(a[7]), .B(a[2]), .Y(n829) );
  NAND2X1 U86 ( .A(n533), .B(a[0]), .Y(n815) );
  INVX1 U87 ( .A(n685), .Y(n907) );
  NAND2X1 U88 ( .A(n864), .B(n540), .Y(n809) );
  NAND2X1 U89 ( .A(n872), .B(n556), .Y(n685) );
  INVX1 U90 ( .A(n635), .Y(n908) );
  NOR2X1 U91 ( .A(n550), .B(n598), .Y(n724) );
  NOR2X1 U92 ( .A(n874), .B(n861), .Y(n676) );
  NAND2X1 U93 ( .A(n701), .B(n540), .Y(n761) );
  INVX1 U94 ( .A(n622), .Y(n874) );
  INVX1 U95 ( .A(n757), .Y(n863) );
  INVX1 U96 ( .A(n716), .Y(n875) );
  INVX1 U97 ( .A(n695), .Y(n872) );
  INVX4 U98 ( .A(n536), .Y(n556) );
  NOR2BX1 U99 ( .AN(n709), .B(n854), .Y(n835) );
  NOR2X1 U100 ( .A(n870), .B(n853), .Y(n597) );
  NOR2X1 U101 ( .A(n873), .B(n862), .Y(n637) );
  NAND2X1 U102 ( .A(n889), .B(n700), .Y(n740) );
  INVX1 U103 ( .A(n805), .Y(n853) );
  NAND2X1 U104 ( .A(n889), .B(n675), .Y(n800) );
  INVX1 U105 ( .A(n690), .Y(n868) );
  INVX1 U106 ( .A(n700), .Y(n864) );
  NOR2X1 U107 ( .A(n866), .B(n868), .Y(n726) );
  INVX1 U108 ( .A(n675), .Y(n886) );
  OAI221XL U109 ( .A0(n865), .A1(n545), .B0(n825), .B1(n542), .C0(n905), .Y(
        n576) );
  INVX1 U110 ( .A(n724), .Y(n905) );
  INVX1 U111 ( .A(n796), .Y(n888) );
  NOR2X1 U112 ( .A(n864), .B(n854), .Y(n825) );
  INVX1 U113 ( .A(n711), .Y(n882) );
  NOR2X1 U114 ( .A(n861), .B(n868), .Y(n778) );
  INVX1 U115 ( .A(n617), .Y(n865) );
  INVX1 U116 ( .A(n765), .Y(n881) );
  INVX1 U117 ( .A(n836), .Y(n885) );
  INVX1 U118 ( .A(n713), .Y(n879) );
  NAND2X1 U119 ( .A(n860), .B(n535), .Y(n680) );
  OAI22X1 U120 ( .A0(n683), .A1(n813), .B0(n682), .B1(n769), .Y(n687) );
  AOI222X1 U121 ( .A0(n862), .A1(n547), .B0(n556), .B1(n679), .C0(n678), .C1(
        n711), .Y(n683) );
  AOI211X1 U122 ( .A0(n556), .A1(n689), .B0(n681), .C0(n724), .Y(n682) );
  NAND2X1 U123 ( .A(n807), .B(n694), .Y(n679) );
  NOR2X1 U124 ( .A(n877), .B(n866), .Y(n701) );
  OAI22X1 U125 ( .A0(n542), .A1(n716), .B0(n545), .B1(n538), .Y(n681) );
  CLKINVX3 U126 ( .A(n810), .Y(n873) );
  CLKINVX3 U127 ( .A(n742), .Y(n860) );
  AOI22X1 U128 ( .A0(n899), .A1(n832), .B0(n900), .B1(n831), .Y(n845) );
  OAI221XL U129 ( .A0(n825), .A1(n545), .B0(n893), .B1(n543), .C0(n824), .Y(
        n832) );
  OAI221XL U130 ( .A0(n881), .A1(n545), .B0(n872), .B1(n543), .C0(n828), .Y(
        n831) );
  INVX1 U131 ( .A(n819), .Y(n893) );
  NAND2X1 U132 ( .A(n556), .B(n827), .Y(n736) );
  NAND2X1 U133 ( .A(n808), .B(n709), .Y(n695) );
  AOI22X1 U134 ( .A0(n900), .A1(n729), .B0(n901), .B1(n728), .Y(n730) );
  OAI221XL U135 ( .A0(n877), .A1(n551), .B0(n860), .B1(n545), .C0(n723), .Y(
        n729) );
  OAI221XL U136 ( .A0(n536), .A1(n727), .B0(n726), .B1(n545), .C0(n725), .Y(
        n728) );
  AOI211X1 U137 ( .A0(n722), .A1(n556), .B0(n721), .C0(n720), .Y(n723) );
  AOI22X1 U138 ( .A0(n900), .A1(n592), .B0(n901), .B1(n591), .Y(n593) );
  OAI221XL U139 ( .A0(n888), .A1(n545), .B0(n879), .B1(n543), .C0(n590), .Y(
        n591) );
  OAI211X1 U140 ( .A0(n597), .A1(n550), .B0(n635), .C0(n589), .Y(n592) );
  AOI22X1 U141 ( .A0(n888), .A1(n556), .B0(n884), .B1(n554), .Y(n590) );
  AOI22X1 U142 ( .A0(n548), .A1(n860), .B0(n676), .B1(n539), .Y(n589) );
  AOI21X1 U143 ( .A0(n808), .A1(n680), .B0(n550), .Y(n563) );
  INVX1 U144 ( .A(n803), .Y(n916) );
  AND2X2 U145 ( .A(n758), .B(n757), .Y(n794) );
  OAI21XL U146 ( .A0(n758), .A1(n550), .B0(n736), .Y(n657) );
  INVX1 U147 ( .A(n639), .Y(n911) );
  OAI31X1 U148 ( .A0(n721), .A1(n908), .A2(n638), .B0(n898), .Y(n639) );
  OAI21XL U149 ( .A0(n541), .A1(n637), .B0(n636), .Y(n638) );
  INVX1 U150 ( .A(n776), .Y(n876) );
  OAI22X1 U151 ( .A0(n621), .A1(n769), .B0(n620), .B1(n813), .Y(n626) );
  AOI211X1 U152 ( .A0(n556), .A1(n821), .B0(n619), .C0(n618), .Y(n620) );
  AOI221X1 U153 ( .A0(n910), .A1(n535), .B0(n896), .B1(n556), .C0(n616), .Y(
        n621) );
  OAI22X1 U154 ( .A0(n859), .A1(n543), .B0(n550), .B1(n617), .Y(n619) );
  AOI222X1 U155 ( .A0(n867), .A1(n540), .B0(n863), .B1(n554), .C0(n549), .C1(
        n852), .Y(n567) );
  AOI21X1 U156 ( .A0(n873), .A1(n556), .B0(n557), .Y(n558) );
  OAI221XL U157 ( .A0(n551), .A1(n836), .B0(n829), .B1(n819), .C0(n677), .Y(
        n688) );
  AOI2BB2X1 U158 ( .B0(n910), .B1(n535), .A0N(n536), .A1N(n676), .Y(n677) );
  CLKINVX8 U159 ( .A(n546), .Y(n545) );
  CLKINVX3 U160 ( .A(n541), .Y(n539) );
  NOR2X1 U161 ( .A(n545), .B(n535), .Y(n721) );
  AOI211X1 U162 ( .A0(n878), .A1(n540), .B0(n719), .C0(n718), .Y(n731) );
  INVX1 U163 ( .A(n714), .Y(n878) );
  NAND2BX1 U164 ( .AN(n826), .B(n717), .Y(n718) );
  AOI222X1 U165 ( .A0(n916), .A1(n810), .B0(n724), .B1(n873), .C0(n886), .C1(
        n540), .Y(n725) );
  AOI221X1 U166 ( .A0(n602), .A1(n553), .B0(n540), .B1(n612), .C0(n596), .Y(
        n608) );
  OAI221XL U167 ( .A0(n536), .A1(n714), .B0(n545), .B1(n820), .C0(n635), .Y(
        n596) );
  AOI221X1 U168 ( .A0(n916), .A1(n852), .B0(n553), .B1(n810), .C0(n737), .Y(
        n749) );
  OAI2BB1X1 U169 ( .A0N(n781), .A1N(n547), .B0(n736), .Y(n737) );
  OAI221XL U170 ( .A0(n615), .A1(n551), .B0(n545), .B1(n758), .C0(n761), .Y(
        n616) );
  NOR2X1 U171 ( .A(n854), .B(n855), .Y(n615) );
  OAI221XL U172 ( .A0(n869), .A1(n545), .B0(n890), .B1(n543), .C0(n691), .Y(
        n706) );
  INVX1 U173 ( .A(n689), .Y(n869) );
  AOI32X1 U174 ( .A0(n889), .A1(n742), .A2(n556), .B0(n553), .B1(n690), .Y(
        n691) );
  OAI221XL U175 ( .A0(n856), .A1(n551), .B0(n829), .B1(n538), .C0(n629), .Y(
        n641) );
  INVX1 U176 ( .A(n808), .Y(n856) );
  AOI211X1 U177 ( .A0(n875), .A1(n556), .B0(n914), .C0(n628), .Y(n629) );
  INVX1 U178 ( .A(n809), .Y(n914) );
  AOI211X1 U179 ( .A0(n863), .A1(n540), .B0(n909), .C0(n559), .Y(n560) );
  NOR3X1 U180 ( .A(n545), .B(n884), .C(n862), .Y(n559) );
  INVX1 U181 ( .A(n664), .Y(n909) );
  OAI221XL U182 ( .A0(n536), .A1(n755), .B0(n759), .B1(n551), .C0(n754), .Y(
        n773) );
  AOI22X1 U183 ( .A0(n549), .A1(n889), .B0(n875), .B1(n539), .Y(n754) );
  AOI211X1 U184 ( .A0(n554), .A1(n827), .B0(n908), .C0(n826), .Y(n828) );
  CLKINVX3 U185 ( .A(n555), .Y(n551) );
  INVX1 U186 ( .A(n544), .Y(n542) );
  INVX1 U187 ( .A(n798), .Y(n913) );
  AOI221X1 U188 ( .A0(n797), .A1(n552), .B0(n796), .B1(n548), .C0(n795), .Y(
        n798) );
  OAI21XL U189 ( .A0(n536), .A1(n794), .B0(n793), .Y(n795) );
  INVX1 U190 ( .A(n536), .Y(n906) );
  NOR2X1 U191 ( .A(n884), .B(n866), .Y(n744) );
  CLKINVX3 U192 ( .A(n813), .Y(n900) );
  NAND3X1 U193 ( .A(n538), .B(n810), .C(n540), .Y(n834) );
  NAND2X1 U194 ( .A(n709), .B(n781), .Y(n833) );
  NAND2X1 U195 ( .A(n807), .B(n781), .Y(n838) );
  NAND2X1 U196 ( .A(n808), .B(n655), .Y(n765) );
  NAND2X1 U197 ( .A(n538), .B(n757), .Y(n612) );
  NOR2BX1 U198 ( .AN(n694), .B(n855), .Y(n759) );
  AOI21X1 U199 ( .A0(n742), .A1(n741), .B0(n536), .Y(n743) );
  OAI221XL U200 ( .A0(n887), .A1(n550), .B0(n802), .B1(n541), .C0(n783), .Y(
        n788) );
  INVX1 U201 ( .A(n838), .Y(n887) );
  AOI22X1 U202 ( .A0(n874), .A1(n548), .B0(n556), .B1(n782), .Y(n783) );
  AOI22X1 U203 ( .A0(n866), .A1(n546), .B0(n555), .B1(n810), .Y(n684) );
  AOI22X1 U204 ( .A0(n547), .A1(n612), .B0(n873), .B1(n539), .Y(n573) );
  NOR2X1 U205 ( .A(n785), .B(n536), .Y(n826) );
  NAND2X1 U206 ( .A(n680), .B(n781), .Y(n796) );
  INVX1 U207 ( .A(n769), .Y(n898) );
  NAND2X1 U208 ( .A(n694), .B(n680), .Y(n689) );
  CLKINVX3 U209 ( .A(n785), .Y(n867) );
  NAND2X1 U210 ( .A(n694), .B(n714), .Y(n663) );
  NOR2X1 U211 ( .A(n859), .B(n799), .Y(n802) );
  AOI211X1 U212 ( .A0(n556), .A1(n617), .B0(n588), .C0(n587), .Y(n594) );
  OAI2BB2X1 U213 ( .B0(n545), .B1(n740), .A0N(n735), .A1N(n540), .Y(n588) );
  AOI21X1 U214 ( .A0(n622), .A1(n586), .B0(n550), .Y(n587) );
  NAND2X1 U215 ( .A(n538), .B(n709), .Y(n797) );
  NAND2X1 U216 ( .A(n785), .B(n821), .Y(n696) );
  NAND2X1 U217 ( .A(n820), .B(n758), .Y(n735) );
  AOI21X1 U218 ( .A0(n556), .A1(n823), .B0(n822), .Y(n824) );
  AOI21X1 U219 ( .A0(n821), .A1(n820), .B0(n550), .Y(n822) );
  INVX1 U220 ( .A(n586), .Y(n858) );
  AOI22X1 U221 ( .A0(n899), .A1(n780), .B0(n901), .B1(n779), .Y(n790) );
  OAI221XL U222 ( .A0(n858), .A1(n551), .B0(n892), .B1(n536), .C0(n774), .Y(
        n780) );
  OAI221XL U223 ( .A0(n778), .A1(n545), .B0(n895), .B1(n551), .C0(n777), .Y(
        n779) );
  AOI2BB2X1 U224 ( .B0(n539), .B1(n836), .A0N(n545), .A1N(n802), .Y(n774) );
  INVX1 U225 ( .A(n715), .Y(n894) );
  INVX1 U226 ( .A(n624), .Y(n910) );
  INVX1 U227 ( .A(n823), .Y(n890) );
  AOI221XL U228 ( .A0(n556), .A1(n871), .B0(n548), .B1(n800), .C0(n599), .Y(
        n607) );
  INVX1 U229 ( .A(n597), .Y(n871) );
  OAI32X1 U230 ( .A0(n829), .A1(n860), .A2(n598), .B0(n886), .B1(n551), .Y(
        n599) );
  INVX1 U231 ( .A(n727), .Y(n892) );
  OAI221XL U232 ( .A0(n867), .A1(n545), .B0(n891), .B1(n543), .C0(n760), .Y(
        n772) );
  INVX1 U233 ( .A(n756), .Y(n891) );
  AOI22X1 U234 ( .A0(n759), .A1(n906), .B0(n794), .B1(n552), .Y(n760) );
  INVX1 U235 ( .A(n782), .Y(n896) );
  INVX1 U236 ( .A(n775), .Y(n895) );
  OAI221XL U237 ( .A0(n883), .A1(n551), .B0(n865), .B1(n545), .C0(n786), .Y(
        n787) );
  INVX1 U238 ( .A(n827), .Y(n883) );
  AOI31X1 U239 ( .A0(n821), .A1(n785), .A2(n556), .B0(n912), .Y(n786) );
  INVX1 U240 ( .A(n834), .Y(n912) );
  INVX1 U241 ( .A(n738), .Y(n904) );
  INVX1 U242 ( .A(n539), .Y(n543) );
  AOI211X1 U243 ( .A0(n901), .A1(n627), .B0(n626), .C0(n625), .Y(n643) );
  AOI211X1 U244 ( .A0(n901), .A1(n641), .B0(n640), .C0(n911), .Y(n642) );
  OAI2BB2X1 U245 ( .B0(n614), .B1(n613), .A0N(n744), .A1N(n614), .Y(n627) );
  AOI211X1 U246 ( .A0(n901), .A1(n688), .B0(n687), .C0(n686), .Y(n708) );
  AOI211X1 U247 ( .A0(n900), .A1(n706), .B0(n705), .C0(n704), .Y(n707) );
  AOI31X1 U248 ( .A0(n685), .A1(n793), .A2(n684), .B0(n767), .Y(n686) );
  AOI22X1 U249 ( .A0(n533), .A1(n669), .B0(n668), .B1(n897), .Y(n670) );
  OAI221XL U250 ( .A0(n862), .A1(n551), .B0(n545), .B1(n663), .C0(n662), .Y(
        n669) );
  OAI221XL U251 ( .A0(n882), .A1(n545), .B0(n541), .B1(n742), .C0(n667), .Y(
        n668) );
  AOI21X1 U252 ( .A0(n890), .A1(n906), .B0(n661), .Y(n662) );
  AOI22X1 U253 ( .A0(n575), .A1(n897), .B0(n533), .B1(n574), .Y(n581) );
  OAI221XL U254 ( .A0(n536), .A1(n757), .B0(n637), .B1(n545), .C0(n572), .Y(
        n575) );
  OAI211X1 U255 ( .A0(n835), .A1(n550), .B0(n736), .C0(n573), .Y(n574) );
  AOI2BB2X1 U256 ( .B0(n539), .B1(n727), .A0N(n550), .A1N(n744), .Y(n572) );
  OAI22X1 U257 ( .A0(n634), .A1(n813), .B0(n633), .B1(n767), .Y(n640) );
  AOI221XL U258 ( .A0(n549), .A1(n740), .B0(n799), .B1(n850), .C0(n632), .Y(
        n633) );
  AOI221XL U259 ( .A0(n867), .A1(n916), .B0(n547), .B1(n713), .C0(n630), .Y(
        n634) );
  OAI32X1 U260 ( .A0(n738), .A1(n860), .A2(n850), .B0(n631), .B1(n904), .Y(
        n632) );
  OAI22X1 U261 ( .A0(n770), .A1(n769), .B0(n768), .B1(n767), .Y(n771) );
  AOI211X1 U262 ( .A0(n881), .A1(n850), .B0(n766), .C0(n907), .Y(n768) );
  AOI221XL U263 ( .A0(n862), .A1(n554), .B0(n547), .B1(n776), .C0(n764), .Y(
        n770) );
  OAI22X1 U264 ( .A0(n541), .A1(n852), .B0(n886), .B1(n550), .Y(n766) );
  OAI22X1 U265 ( .A0(n816), .A1(n815), .B0(n814), .B1(n813), .Y(n817) );
  AOI221XL U266 ( .A0(n549), .A1(n812), .B0(n876), .B1(n540), .C0(n811), .Y(
        n814) );
  AOI221X1 U267 ( .A0(n556), .A1(n808), .B0(n552), .B1(n807), .C0(n806), .Y(
        n816) );
  OAI221XL U268 ( .A0(n536), .A1(n810), .B0(n879), .B1(n551), .C0(n809), .Y(
        n811) );
  AOI211X1 U269 ( .A0(n868), .A1(n556), .B0(n652), .C0(n651), .Y(n653) );
  AOI31X1 U270 ( .A0(n809), .A1(n717), .A2(n650), .B0(n533), .Y(n651) );
  OAI22X1 U271 ( .A0(n857), .A1(n803), .B0(n649), .B1(n897), .Y(n652) );
  AOI2BB2X1 U272 ( .B0(n853), .B1(n552), .A0N(n833), .A1N(n545), .Y(n650) );
  AOI2BB2X1 U273 ( .B0(n659), .B1(n897), .A0N(n897), .A1N(n658), .Y(n671) );
  OAI221XL U274 ( .A0(n877), .A1(n551), .B0(n545), .B1(n807), .C0(n656), .Y(
        n659) );
  AOI221XL U275 ( .A0(n548), .A1(n676), .B0(n711), .B1(n540), .C0(n657), .Y(
        n658) );
  AOI22X1 U276 ( .A0(n539), .A1(n765), .B0(n873), .B1(n903), .Y(n656) );
  AOI22X1 U277 ( .A0(n534), .A1(n610), .B0(n609), .B1(n902), .Y(n611) );
  OAI221XL U278 ( .A0(n595), .A1(n767), .B0(n594), .B1(n769), .C0(n593), .Y(
        n610) );
  OAI221XL U279 ( .A0(n608), .A1(n767), .B0(n607), .B1(n769), .C0(n606), .Y(
        n609) );
  AOI22X1 U281 ( .A0(n752), .A1(n902), .B0(n534), .B1(n751), .Y(n753) );
  OAI221XL U282 ( .A0(n750), .A1(n815), .B0(n749), .B1(n769), .C0(n748), .Y(
        n751) );
  OAI221XL U283 ( .A0(n732), .A1(n769), .B0(n731), .B1(n767), .C0(n730), .Y(
        n752) );
  AOI22X1 U284 ( .A0(n554), .A1(n532), .B0(n539), .B1(n857), .Y(n631) );
  AOI22X1 U285 ( .A0(n533), .A1(n562), .B0(n561), .B1(n897), .Y(n571) );
  OAI221XL U286 ( .A0(n880), .A1(n545), .B0(n829), .B1(n889), .C0(n558), .Y(
        n562) );
  OAI221XL U287 ( .A0(n532), .A1(n803), .B0(n722), .B1(n551), .C0(n560), .Y(
        n561) );
  INVX1 U288 ( .A(n663), .Y(n880) );
  AOI22X1 U289 ( .A0(n901), .A1(n605), .B0(n900), .B1(n604), .Y(n606) );
  OAI21XL U290 ( .A0(n602), .A1(n536), .B0(n601), .Y(n605) );
  OAI221XL U291 ( .A0(n551), .A1(n810), .B0(n835), .B1(n545), .C0(n603), .Y(
        n604) );
  AOI31X1 U292 ( .A0(n538), .A1(n742), .A2(n600), .B0(n910), .Y(n601) );
  CLKINVX3 U293 ( .A(n532), .Y(n852) );
  OAI21XL U294 ( .A0(n545), .A1(n537), .B0(n803), .Y(n647) );
  NAND2X1 U295 ( .A(n860), .B(n531), .Y(n755) );
  AOI21X1 U296 ( .A0(n699), .A1(n680), .B0(n545), .Y(n628) );
  INVX1 U297 ( .A(n531), .Y(n849) );
  OAI21XL U298 ( .A0(n850), .A1(n622), .B0(n550), .Y(n600) );
  OAI21XL U299 ( .A0(n536), .A1(n805), .B0(n763), .Y(n764) );
  AOI31X1 U300 ( .A0(n812), .A1(n903), .A2(n762), .B0(n915), .Y(n763) );
  INVX1 U301 ( .A(n761), .Y(n915) );
  OAI2BB1X1 U302 ( .A0N(n845), .A1N(n844), .B0(n902), .Y(n846) );
  AOI22X1 U303 ( .A0(n901), .A1(n843), .B0(n898), .B1(n842), .Y(n844) );
  AOI211X1 U304 ( .A0(n884), .A1(n540), .B0(n648), .C0(n647), .Y(n649) );
  OAI222X1 U305 ( .A0(n551), .A1(n807), .B0(n850), .B1(n693), .C0(n545), .C1(
        n821), .Y(n648) );
  NAND2X1 U306 ( .A(n861), .B(n552), .Y(n636) );
  OAI2BB1X1 U307 ( .A0N(n790), .A1N(n789), .B0(n534), .Y(n791) );
  AOI22X1 U308 ( .A0(n900), .A1(n788), .B0(n898), .B1(n787), .Y(n789) );
  NOR2BX1 U309 ( .AN(n660), .B(n876), .Y(n722) );
  BUFX3 U310 ( .A(n841), .Y(n536) );
  NAND2X1 U311 ( .A(n850), .B(n903), .Y(n841) );
  OAI221XL U312 ( .A0(n531), .A1(n664), .B0(n542), .B1(n709), .C0(n636), .Y(
        n630) );
  BUFX3 U313 ( .A(n784), .Y(n538) );
  NAND2X1 U314 ( .A(n531), .B(n537), .Y(n784) );
  AOI211X1 U315 ( .A0(n540), .A1(n852), .B0(n585), .C0(n647), .Y(n595) );
  OAI222X1 U316 ( .A0(n551), .A1(n756), .B0(n584), .B1(n536), .C0(n545), .C1(
        n889), .Y(n585) );
  AOI21X1 U317 ( .A0(n537), .A1(n535), .B0(n858), .Y(n584) );
  AOI211X1 U318 ( .A0(n533), .A1(n569), .B0(n848), .C0(n568), .Y(n570) );
  OAI221XL U319 ( .A0(n545), .A1(n807), .B0(n602), .B1(n542), .C0(n564), .Y(
        n569) );
  AOI21X1 U320 ( .A0(n567), .A1(n566), .B0(n533), .Y(n568) );
  AOI31X1 U321 ( .A0(n556), .A1(n565), .A2(n884), .B0(n563), .Y(n564) );
  INVX1 U322 ( .A(n830), .Y(n546) );
  INVX1 U323 ( .A(n840), .Y(n554) );
  INVX1 U324 ( .A(n840), .Y(n555) );
  INVX1 U325 ( .A(n544), .Y(n541) );
  INVX1 U326 ( .A(n829), .Y(n544) );
  AOI22X1 U327 ( .A0(n533), .A1(n646), .B0(n645), .B1(n897), .Y(n654) );
  OAI222X1 U328 ( .A0(n545), .A1(n782), .B0(n551), .B1(n660), .C0(n894), .C1(
        n541), .Y(n646) );
  OAI221XL U329 ( .A0(n892), .A1(n536), .B0(n551), .B1(n819), .C0(n644), .Y(
        n645) );
  AOI2BB2X1 U330 ( .B0(n835), .B1(n539), .A0N(n545), .A1N(n726), .Y(n644) );
  NAND2X1 U331 ( .A(n699), .B(n622), .Y(n775) );
  NOR2BX1 U332 ( .AN(n660), .B(n862), .Y(n602) );
  AOI21X1 U333 ( .A0(n690), .A1(n758), .B0(n903), .Y(n661) );
  AOI22X1 U334 ( .A0(n900), .A1(n747), .B0(n899), .B1(n746), .Y(n748) );
  OAI221XL U335 ( .A0(n860), .A1(n545), .B0(n543), .B1(n807), .C0(n745), .Y(
        n746) );
  OAI221XL U336 ( .A0(n885), .A1(n536), .B0(n545), .B1(n740), .C0(n739), .Y(
        n747) );
  AOI21X1 U337 ( .A0(n744), .A1(n552), .B0(n743), .Y(n745) );
  AOI22X1 U338 ( .A0(n556), .A1(n857), .B0(n539), .B1(n776), .Y(n777) );
  AOI22X1 U339 ( .A0(n549), .A1(n838), .B0(n882), .B1(n539), .Y(n839) );
  AOI31X1 U340 ( .A0(n703), .A1(n793), .A2(n702), .B0(n815), .Y(n704) );
  OAI2BB1X1 U341 ( .A0N(n700), .A1N(n699), .B0(n553), .Y(n703) );
  AOI22X1 U342 ( .A0(n894), .A1(n556), .B0(n701), .B1(n547), .Y(n702) );
  NAND2X1 U343 ( .A(n699), .B(n805), .Y(n715) );
  NAND2X1 U344 ( .A(n660), .B(n586), .Y(n756) );
  AOI21X1 U345 ( .A0(n660), .A1(n741), .B0(n545), .Y(n618) );
  AOI21X1 U346 ( .A0(n812), .A1(n538), .B0(n542), .Y(n720) );
  NAND2X1 U347 ( .A(n906), .B(n531), .Y(n717) );
  OAI21XL U348 ( .A0(n850), .A1(n680), .B0(n550), .Y(n678) );
  XNOR2X1 U349 ( .A(n903), .B(n531), .Y(n738) );
  NAND2X1 U350 ( .A(n539), .B(n537), .Y(n793) );
  XNOR2X1 U351 ( .A(n850), .B(n531), .Y(n762) );
  AOI21X1 U352 ( .A0(n833), .A1(n850), .B0(n556), .Y(n837) );
  AOI221X1 U353 ( .A0(n877), .A1(n540), .B0(n553), .B1(n735), .C0(n734), .Y(
        n750) );
  AOI21X1 U354 ( .A0(n536), .A1(n733), .B0(n799), .Y(n734) );
  OAI21XL U355 ( .A0(n861), .A1(n853), .B0(n850), .Y(n733) );
  AOI222X1 U356 ( .A0(n549), .A1(n713), .B0(n712), .B1(n711), .C0(n556), .C1(
        n537), .Y(n732) );
  OAI21XL U357 ( .A0(n850), .A1(n709), .B0(n550), .Y(n712) );
  AOI31X1 U358 ( .A0(n761), .A1(n624), .A2(n623), .B0(n767), .Y(n625) );
  AOI22X1 U359 ( .A0(n775), .A1(n850), .B0(n894), .B1(n553), .Y(n623) );
  INVX1 U360 ( .A(n830), .Y(n547) );
  INVX1 U361 ( .A(n830), .Y(n549) );
  INVX1 U362 ( .A(n830), .Y(n548) );
  XOR2X1 U363 ( .A(n533), .B(n531), .Y(n565) );
  INVX1 U364 ( .A(n840), .Y(n552) );
  INVX1 U365 ( .A(n840), .Y(n553) );
  NOR2BX1 U366 ( .AN(n830), .B(n554), .Y(n614) );
  AOI22X1 U367 ( .A0(n581), .A1(a[0]), .B0(n580), .B1(n579), .Y(n582) );
  AOI31X1 U368 ( .A0(n717), .A1(n848), .A2(n571), .B0(n570), .Y(n583) );
  AOI22X1 U369 ( .A0(n576), .A1(n897), .B0(n556), .B1(n833), .Y(n580) );
  AOI22X1 U370 ( .A0(n673), .A1(n902), .B0(n534), .B1(n672), .Y(n674) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n654), .B0(n653), .B1(n848), .Y(n673) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n671), .B0(n670), .B1(n848), .Y(n672) );
  OAI22X1 U373 ( .A0(n698), .A1(n767), .B0(n697), .B1(n769), .Y(n705) );
  AOI221X1 U374 ( .A0(n548), .A1(n693), .B0(n556), .B1(n797), .C0(n692), .Y(
        n698) );
  AOI222X1 U375 ( .A0(n759), .A1(n547), .B0(a[2]), .B1(n696), .C0(n556), .C1(
        n695), .Y(n697) );
  OAI22X1 U376 ( .A0(n888), .A1(n543), .B0(n550), .B1(n537), .Y(n692) );
  NOR2X1 U377 ( .A(n863), .B(n861), .Y(n804) );
  BUFX3 U378 ( .A(n710), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n852), .Y(n710) );
  AOI221X1 U380 ( .A0(n916), .A1(n785), .B0(n851), .B1(n666), .C0(n665), .Y(
        n667) );
  NOR3X1 U381 ( .A(n851), .B(a[7]), .C(n860), .Y(n665) );
  INVX1 U382 ( .A(n762), .Y(n851) );
  OAI21XL U383 ( .A0(n857), .A1(n550), .B0(n664), .Y(n666) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI22X1 U385 ( .A0(n882), .A1(n850), .B0(a[2]), .B1(n612), .Y(n613) );
  CLKINVX3 U386 ( .A(a[0]), .Y(n848) );
  AOI211X1 U387 ( .A0(n724), .A1(n578), .B0(n577), .C0(a[0]), .Y(n579) );
  NAND2X1 U388 ( .A(n781), .B(n805), .Y(n578) );
  AOI21X1 U389 ( .A0(n803), .A1(n624), .B0(n897), .Y(n577) );
  BUFX3 U390 ( .A(a[5]), .Y(n533) );
  OAI221XL U391 ( .A0(n536), .A1(n808), .B0(n802), .B1(n545), .C0(n801), .Y(
        n818) );
  AOI22X1 U392 ( .A0(n539), .A1(n800), .B0(n799), .B1(a[2]), .Y(n801) );
  AOI33X1 U393 ( .A0(n532), .A1(n540), .A2(n904), .B0(n738), .B1(n742), .B2(
        a[2]), .Y(n739) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_sbox_17 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916;

  OAI221X4 U4 ( .A0(n857), .A1(n536), .B0(n862), .B1(n551), .C0(n839), .Y(n842) );
  OAI221X4 U6 ( .A0(n837), .A1(n836), .B0(n835), .B1(n551), .C0(n834), .Y(n843) );
  OAI222X4 U75 ( .A0(n551), .A1(n716), .B0(n742), .B1(n803), .C0(n545), .C1(
        n715), .Y(n719) );
  OAI32X4 U280 ( .A0(n551), .A1(n867), .A2(n870), .B0(n829), .B1(n820), .Y(
        n557) );
  AOI221X1 U1 ( .A0(n858), .A1(a[2]), .B0(n826), .B1(n565), .C0(n916), .Y(n566) );
  INVX1 U2 ( .A(a[7]), .Y(n903) );
  NAND2X1 U3 ( .A(n867), .B(n531), .Y(n694) );
  NAND2X2 U5 ( .A(n532), .B(n857), .Y(n742) );
  NAND2X1 U7 ( .A(n884), .B(n531), .Y(n781) );
  NAND2X2 U8 ( .A(n857), .B(n852), .Y(n785) );
  NAND2X1 U9 ( .A(n532), .B(n535), .Y(n820) );
  NAND2X1 U10 ( .A(n531), .B(n742), .Y(n821) );
  NAND2X2 U11 ( .A(n537), .B(n742), .Y(n810) );
  OAI222X1 U12 ( .A0(n829), .A1(n805), .B0(n804), .B1(n545), .C0(a[4]), .C1(
        n803), .Y(n806) );
  NAND2X2 U13 ( .A(n857), .B(n535), .Y(n807) );
  NAND2X2 U14 ( .A(n531), .B(n532), .Y(n808) );
  CLKINVX3 U15 ( .A(a[2]), .Y(n850) );
  NAND2X1 U16 ( .A(n533), .B(n848), .Y(n813) );
  CLKINVX3 U17 ( .A(n533), .Y(n897) );
  NAND2X2 U18 ( .A(a[0]), .B(n897), .Y(n767) );
  NAND2X2 U19 ( .A(n848), .B(n897), .Y(n769) );
  NAND2X1 U20 ( .A(a[2]), .B(n903), .Y(n840) );
  NAND2X1 U21 ( .A(a[7]), .B(n850), .Y(n830) );
  AOI21XL U22 ( .A0(n916), .A1(a[4]), .B0(n907), .Y(n603) );
  NAND2X1 U23 ( .A(a[4]), .B(n535), .Y(n660) );
  NAND2X1 U24 ( .A(n531), .B(a[4]), .Y(n699) );
  NAND2X2 U25 ( .A(n532), .B(a[4]), .Y(n812) );
  CLKINVX3 U26 ( .A(a[4]), .Y(n857) );
  NAND2X1 U27 ( .A(n870), .B(n556), .Y(n635) );
  CLKINVX3 U28 ( .A(n543), .Y(n540) );
  INVX1 U29 ( .A(n598), .Y(n889) );
  NAND2X1 U30 ( .A(n810), .B(n535), .Y(n709) );
  NAND2X1 U31 ( .A(n877), .B(n535), .Y(n714) );
  NAND2X1 U32 ( .A(n873), .B(n535), .Y(n622) );
  NAND2X1 U33 ( .A(n538), .B(n655), .Y(n711) );
  NAND2X1 U34 ( .A(n776), .B(n709), .Y(n716) );
  NAND2X1 U35 ( .A(n808), .B(n714), .Y(n713) );
  INVX1 U36 ( .A(n538), .Y(n870) );
  INVX1 U37 ( .A(n741), .Y(n866) );
  NOR2X1 U38 ( .A(n535), .B(n884), .Y(n598) );
  CLKINVX3 U39 ( .A(n555), .Y(n550) );
  NAND2X1 U40 ( .A(n535), .B(n852), .Y(n805) );
  NAND2X1 U41 ( .A(n867), .B(n535), .Y(n690) );
  NAND2X1 U42 ( .A(n785), .B(n535), .Y(n700) );
  NAND2X1 U43 ( .A(n884), .B(n535), .Y(n675) );
  NAND2X1 U44 ( .A(n742), .B(n535), .Y(n757) );
  NAND2X1 U45 ( .A(n694), .B(n675), .Y(n836) );
  INVX1 U46 ( .A(n821), .Y(n862) );
  NAND2X1 U47 ( .A(n808), .B(n700), .Y(n617) );
  INVX1 U48 ( .A(n755), .Y(n861) );
  INVX1 U49 ( .A(n693), .Y(n854) );
  INVX1 U50 ( .A(n807), .Y(n859) );
  INVX1 U51 ( .A(n820), .Y(n855) );
  BUFX3 U52 ( .A(n849), .Y(n535) );
  NAND2X1 U53 ( .A(n873), .B(n531), .Y(n776) );
  NAND2X1 U54 ( .A(n531), .B(n539), .Y(n803) );
  NAND2X1 U55 ( .A(n531), .B(n810), .Y(n758) );
  NAND2X1 U56 ( .A(n531), .B(n785), .Y(n741) );
  INVX1 U57 ( .A(n753), .Y(d[5]) );
  INVX1 U58 ( .A(n611), .Y(d[1]) );
  INVX1 U59 ( .A(n537), .Y(n877) );
  NAND2X1 U60 ( .A(n906), .B(n532), .Y(n664) );
  NAND2X1 U61 ( .A(n812), .B(n776), .Y(n827) );
  NOR2X1 U62 ( .A(n537), .B(n535), .Y(n799) );
  NAND2X1 U63 ( .A(n812), .B(n535), .Y(n655) );
  CLKINVX3 U64 ( .A(n812), .Y(n884) );
  NAND2X1 U65 ( .A(n531), .B(n852), .Y(n693) );
  NAND2X1 U66 ( .A(n531), .B(n857), .Y(n586) );
  NAND2BX1 U67 ( .AN(n799), .B(n660), .Y(n727) );
  INVX1 U68 ( .A(n767), .Y(n899) );
  NAND2X1 U69 ( .A(n699), .B(n655), .Y(n782) );
  NAND2BX1 U70 ( .AN(n830), .B(n537), .Y(n624) );
  NAND2X1 U71 ( .A(n699), .B(n690), .Y(n819) );
  NAND2X1 U72 ( .A(n660), .B(n781), .Y(n823) );
  CLKINVX3 U73 ( .A(n534), .Y(n902) );
  CLKINVX3 U74 ( .A(n815), .Y(n901) );
  INVX1 U76 ( .A(n674), .Y(d[3]) );
  BUFX3 U77 ( .A(a[1]), .Y(n531) );
  NAND2X1 U78 ( .A(a[7]), .B(a[2]), .Y(n829) );
  NAND2X1 U79 ( .A(n533), .B(a[0]), .Y(n815) );
  INVX1 U80 ( .A(n685), .Y(n907) );
  NAND2X1 U81 ( .A(n864), .B(n540), .Y(n809) );
  NAND2X1 U82 ( .A(n872), .B(n556), .Y(n685) );
  INVX1 U83 ( .A(n635), .Y(n908) );
  NOR2X1 U84 ( .A(n550), .B(n598), .Y(n724) );
  NOR2X1 U85 ( .A(n874), .B(n861), .Y(n676) );
  NAND2X1 U86 ( .A(n701), .B(n540), .Y(n761) );
  INVX1 U87 ( .A(n622), .Y(n874) );
  INVX1 U88 ( .A(n757), .Y(n863) );
  INVX1 U89 ( .A(n716), .Y(n875) );
  INVX1 U90 ( .A(n695), .Y(n872) );
  INVX4 U91 ( .A(n536), .Y(n556) );
  NOR2BX1 U92 ( .AN(n709), .B(n854), .Y(n835) );
  NOR2X1 U93 ( .A(n870), .B(n853), .Y(n597) );
  NOR2X1 U94 ( .A(n873), .B(n862), .Y(n637) );
  NAND2X1 U95 ( .A(n889), .B(n700), .Y(n740) );
  INVX1 U96 ( .A(n805), .Y(n853) );
  NAND2X1 U97 ( .A(n889), .B(n675), .Y(n800) );
  INVX1 U98 ( .A(n690), .Y(n868) );
  INVX1 U99 ( .A(n700), .Y(n864) );
  NOR2X1 U100 ( .A(n866), .B(n868), .Y(n726) );
  INVX1 U101 ( .A(n675), .Y(n886) );
  OAI221XL U102 ( .A0(n865), .A1(n545), .B0(n825), .B1(n829), .C0(n905), .Y(
        n576) );
  INVX1 U103 ( .A(n724), .Y(n905) );
  INVX1 U104 ( .A(n796), .Y(n888) );
  NOR2X1 U105 ( .A(n864), .B(n854), .Y(n825) );
  INVX1 U106 ( .A(n711), .Y(n882) );
  NOR2X1 U107 ( .A(n861), .B(n868), .Y(n778) );
  INVX1 U108 ( .A(n617), .Y(n865) );
  INVX1 U109 ( .A(n765), .Y(n881) );
  INVX1 U110 ( .A(n836), .Y(n885) );
  INVX1 U111 ( .A(n713), .Y(n879) );
  NAND2X1 U112 ( .A(n860), .B(n535), .Y(n680) );
  OAI22X1 U113 ( .A0(n683), .A1(n813), .B0(n682), .B1(n769), .Y(n687) );
  AOI222X1 U114 ( .A0(n862), .A1(n547), .B0(n556), .B1(n679), .C0(n678), .C1(
        n711), .Y(n683) );
  AOI211X1 U115 ( .A0(n556), .A1(n689), .B0(n681), .C0(n724), .Y(n682) );
  NAND2X1 U116 ( .A(n807), .B(n694), .Y(n679) );
  NOR2X1 U117 ( .A(n877), .B(n866), .Y(n701) );
  OAI22X1 U118 ( .A0(n542), .A1(n716), .B0(n545), .B1(n538), .Y(n681) );
  CLKINVX3 U119 ( .A(n810), .Y(n873) );
  NAND2X1 U120 ( .A(n709), .B(n781), .Y(n833) );
  CLKINVX3 U121 ( .A(n742), .Y(n860) );
  AOI22X1 U122 ( .A0(n899), .A1(n832), .B0(n900), .B1(n831), .Y(n845) );
  OAI221XL U123 ( .A0(n825), .A1(n545), .B0(n893), .B1(n542), .C0(n824), .Y(
        n832) );
  OAI221XL U124 ( .A0(n881), .A1(n545), .B0(n872), .B1(n542), .C0(n828), .Y(
        n831) );
  INVX1 U125 ( .A(n819), .Y(n893) );
  NAND2X1 U126 ( .A(n556), .B(n827), .Y(n736) );
  NAND2X1 U127 ( .A(n808), .B(n709), .Y(n695) );
  AOI22X1 U128 ( .A0(n900), .A1(n729), .B0(n901), .B1(n728), .Y(n730) );
  OAI221XL U129 ( .A0(n877), .A1(n551), .B0(n860), .B1(n545), .C0(n723), .Y(
        n729) );
  OAI221XL U130 ( .A0(n536), .A1(n727), .B0(n726), .B1(n545), .C0(n725), .Y(
        n728) );
  AOI211X1 U131 ( .A0(n722), .A1(n556), .B0(n721), .C0(n720), .Y(n723) );
  AOI22X1 U132 ( .A0(n900), .A1(n592), .B0(n901), .B1(n591), .Y(n593) );
  OAI221XL U133 ( .A0(n888), .A1(n545), .B0(n879), .B1(n543), .C0(n590), .Y(
        n591) );
  OAI211X1 U134 ( .A0(n597), .A1(n550), .B0(n635), .C0(n589), .Y(n592) );
  AOI22X1 U135 ( .A0(n888), .A1(n556), .B0(n884), .B1(n554), .Y(n590) );
  AOI22X1 U136 ( .A0(n548), .A1(n860), .B0(n676), .B1(n539), .Y(n589) );
  AOI21X1 U137 ( .A0(n808), .A1(n680), .B0(n550), .Y(n563) );
  INVX1 U138 ( .A(n803), .Y(n916) );
  AND2X2 U139 ( .A(n758), .B(n757), .Y(n794) );
  NAND2X1 U140 ( .A(n538), .B(n709), .Y(n797) );
  OAI21XL U141 ( .A0(n758), .A1(n550), .B0(n736), .Y(n657) );
  INVX1 U142 ( .A(n639), .Y(n911) );
  OAI31X1 U143 ( .A0(n721), .A1(n908), .A2(n638), .B0(n898), .Y(n639) );
  OAI21XL U144 ( .A0(n541), .A1(n637), .B0(n636), .Y(n638) );
  INVX1 U145 ( .A(n776), .Y(n876) );
  OAI22X1 U146 ( .A0(n621), .A1(n769), .B0(n620), .B1(n813), .Y(n626) );
  AOI211X1 U147 ( .A0(n556), .A1(n821), .B0(n619), .C0(n618), .Y(n620) );
  AOI221X1 U148 ( .A0(n910), .A1(n535), .B0(n896), .B1(n556), .C0(n616), .Y(
        n621) );
  OAI22X1 U149 ( .A0(n859), .A1(n542), .B0(n550), .B1(n617), .Y(n619) );
  AOI222X1 U150 ( .A0(n867), .A1(n540), .B0(n863), .B1(n554), .C0(n548), .C1(
        n852), .Y(n567) );
  AOI21X1 U151 ( .A0(n873), .A1(n906), .B0(n557), .Y(n558) );
  OAI221XL U152 ( .A0(n551), .A1(n836), .B0(n829), .B1(n819), .C0(n677), .Y(
        n688) );
  AOI2BB2X1 U153 ( .B0(n910), .B1(n535), .A0N(n536), .A1N(n676), .Y(n677) );
  CLKINVX8 U154 ( .A(n546), .Y(n545) );
  CLKINVX3 U155 ( .A(n541), .Y(n539) );
  NOR2X1 U156 ( .A(n545), .B(n535), .Y(n721) );
  AOI211X1 U157 ( .A0(n878), .A1(n540), .B0(n719), .C0(n718), .Y(n731) );
  INVX1 U158 ( .A(n714), .Y(n878) );
  NAND2BX1 U159 ( .AN(n826), .B(n717), .Y(n718) );
  AOI222X1 U160 ( .A0(n916), .A1(n810), .B0(n724), .B1(n873), .C0(n886), .C1(
        n540), .Y(n725) );
  AOI221X1 U161 ( .A0(n602), .A1(n553), .B0(n540), .B1(n612), .C0(n596), .Y(
        n608) );
  OAI221XL U162 ( .A0(n536), .A1(n714), .B0(n545), .B1(n820), .C0(n635), .Y(
        n596) );
  AOI221X1 U163 ( .A0(n916), .A1(n852), .B0(n553), .B1(n810), .C0(n737), .Y(
        n749) );
  OAI2BB1X1 U164 ( .A0N(n781), .A1N(n547), .B0(n736), .Y(n737) );
  OAI221XL U165 ( .A0(n615), .A1(n551), .B0(n545), .B1(n758), .C0(n761), .Y(
        n616) );
  NOR2X1 U166 ( .A(n854), .B(n855), .Y(n615) );
  OAI221XL U167 ( .A0(n869), .A1(n545), .B0(n890), .B1(n542), .C0(n691), .Y(
        n706) );
  INVX1 U168 ( .A(n689), .Y(n869) );
  AOI32X1 U169 ( .A0(n889), .A1(n742), .A2(n556), .B0(n553), .B1(n690), .Y(
        n691) );
  OAI221XL U170 ( .A0(n856), .A1(n551), .B0(n829), .B1(n538), .C0(n629), .Y(
        n641) );
  INVX1 U171 ( .A(n808), .Y(n856) );
  AOI211X1 U172 ( .A0(n875), .A1(n556), .B0(n914), .C0(n628), .Y(n629) );
  INVX1 U173 ( .A(n809), .Y(n914) );
  AOI211X1 U174 ( .A0(n863), .A1(n540), .B0(n909), .C0(n559), .Y(n560) );
  NOR3X1 U175 ( .A(n545), .B(n884), .C(n862), .Y(n559) );
  INVX1 U176 ( .A(n664), .Y(n909) );
  OAI221XL U177 ( .A0(n536), .A1(n755), .B0(n759), .B1(n551), .C0(n754), .Y(
        n773) );
  AOI22X1 U178 ( .A0(n549), .A1(n889), .B0(n875), .B1(n539), .Y(n754) );
  AOI211X1 U179 ( .A0(n554), .A1(n827), .B0(n908), .C0(n826), .Y(n828) );
  CLKINVX3 U180 ( .A(n555), .Y(n551) );
  INVX1 U181 ( .A(n798), .Y(n913) );
  AOI221X1 U182 ( .A0(n797), .A1(n552), .B0(n796), .B1(n549), .C0(n795), .Y(
        n798) );
  OAI21XL U183 ( .A0(n536), .A1(n794), .B0(n793), .Y(n795) );
  INVX1 U184 ( .A(n536), .Y(n906) );
  NOR2X1 U185 ( .A(n884), .B(n866), .Y(n744) );
  CLKINVX3 U186 ( .A(n813), .Y(n900) );
  NAND3X1 U187 ( .A(n538), .B(n810), .C(n540), .Y(n834) );
  NAND2X1 U188 ( .A(n807), .B(n781), .Y(n838) );
  NAND2X1 U189 ( .A(n808), .B(n655), .Y(n765) );
  NAND2X1 U190 ( .A(n538), .B(n757), .Y(n612) );
  NOR2BX1 U191 ( .AN(n694), .B(n855), .Y(n759) );
  AOI21X1 U192 ( .A0(n742), .A1(n741), .B0(n536), .Y(n743) );
  OAI221XL U193 ( .A0(n887), .A1(n550), .B0(n802), .B1(n543), .C0(n783), .Y(
        n788) );
  INVX1 U194 ( .A(n838), .Y(n887) );
  AOI22X1 U195 ( .A0(n874), .A1(n549), .B0(n556), .B1(n782), .Y(n783) );
  AOI22X1 U196 ( .A0(n866), .A1(n546), .B0(n555), .B1(n810), .Y(n684) );
  AOI22X1 U197 ( .A0(n547), .A1(n612), .B0(n873), .B1(n539), .Y(n573) );
  NOR2X1 U198 ( .A(n785), .B(n536), .Y(n826) );
  NAND2X1 U199 ( .A(n680), .B(n781), .Y(n796) );
  INVX1 U200 ( .A(n769), .Y(n898) );
  NAND2X1 U201 ( .A(n694), .B(n680), .Y(n689) );
  CLKINVX3 U202 ( .A(n785), .Y(n867) );
  NAND2X1 U203 ( .A(n694), .B(n714), .Y(n663) );
  NOR2X1 U204 ( .A(n859), .B(n799), .Y(n802) );
  AOI211X1 U205 ( .A0(n556), .A1(n617), .B0(n588), .C0(n587), .Y(n594) );
  OAI2BB2X1 U206 ( .B0(n545), .B1(n740), .A0N(n735), .A1N(n540), .Y(n588) );
  AOI21X1 U207 ( .A0(n622), .A1(n586), .B0(n550), .Y(n587) );
  NAND2X1 U208 ( .A(n785), .B(n821), .Y(n696) );
  NAND2X1 U209 ( .A(n820), .B(n758), .Y(n735) );
  AOI21X1 U210 ( .A0(n906), .A1(n823), .B0(n822), .Y(n824) );
  AOI21X1 U211 ( .A0(n821), .A1(n820), .B0(n550), .Y(n822) );
  INVX1 U212 ( .A(n586), .Y(n858) );
  AOI22X1 U213 ( .A0(n899), .A1(n780), .B0(n901), .B1(n779), .Y(n790) );
  OAI221XL U214 ( .A0(n858), .A1(n551), .B0(n892), .B1(n536), .C0(n774), .Y(
        n780) );
  OAI221XL U215 ( .A0(n778), .A1(n545), .B0(n895), .B1(n551), .C0(n777), .Y(
        n779) );
  AOI2BB2X1 U216 ( .B0(n539), .B1(n836), .A0N(n545), .A1N(n802), .Y(n774) );
  INVX1 U217 ( .A(n715), .Y(n894) );
  INVX1 U218 ( .A(n624), .Y(n910) );
  INVX1 U219 ( .A(n823), .Y(n890) );
  AOI221XL U220 ( .A0(n556), .A1(n871), .B0(n548), .B1(n800), .C0(n599), .Y(
        n607) );
  INVX1 U221 ( .A(n597), .Y(n871) );
  OAI32X1 U222 ( .A0(n829), .A1(n860), .A2(n598), .B0(n886), .B1(n551), .Y(
        n599) );
  INVX1 U223 ( .A(n727), .Y(n892) );
  OAI221XL U224 ( .A0(n867), .A1(n545), .B0(n891), .B1(n543), .C0(n760), .Y(
        n772) );
  INVX1 U225 ( .A(n756), .Y(n891) );
  AOI22X1 U226 ( .A0(n759), .A1(n906), .B0(n794), .B1(n554), .Y(n760) );
  INVX1 U227 ( .A(n782), .Y(n896) );
  INVX1 U228 ( .A(n775), .Y(n895) );
  OAI221XL U229 ( .A0(n883), .A1(n551), .B0(n865), .B1(n545), .C0(n786), .Y(
        n787) );
  INVX1 U230 ( .A(n827), .Y(n883) );
  AOI31X1 U231 ( .A0(n821), .A1(n785), .A2(n556), .B0(n912), .Y(n786) );
  INVX1 U232 ( .A(n834), .Y(n912) );
  INVX1 U233 ( .A(n738), .Y(n904) );
  INVX1 U234 ( .A(n544), .Y(n543) );
  INVX1 U235 ( .A(n539), .Y(n542) );
  OAI22X2 U236 ( .A0(n534), .A1(n643), .B0(n642), .B1(n902), .Y(d[2]) );
  AOI211X1 U237 ( .A0(n901), .A1(n627), .B0(n626), .C0(n625), .Y(n643) );
  AOI211X1 U238 ( .A0(n901), .A1(n641), .B0(n640), .C0(n911), .Y(n642) );
  OAI2BB2X1 U239 ( .B0(n614), .B1(n613), .A0N(n744), .A1N(n614), .Y(n627) );
  OAI22X2 U240 ( .A0(n534), .A1(n708), .B0(n707), .B1(n902), .Y(d[4]) );
  AOI211X1 U241 ( .A0(n901), .A1(n688), .B0(n687), .C0(n686), .Y(n708) );
  AOI211X1 U242 ( .A0(n900), .A1(n706), .B0(n705), .C0(n704), .Y(n707) );
  AOI31X1 U243 ( .A0(n685), .A1(n793), .A2(n684), .B0(n767), .Y(n686) );
  OAI21X2 U244 ( .A0(n847), .A1(n902), .B0(n846), .Y(d[7]) );
  OAI2BB1X1 U245 ( .A0N(n845), .A1N(n844), .B0(n902), .Y(n846) );
  AOI221X1 U246 ( .A0(n899), .A1(n913), .B0(n898), .B1(n818), .C0(n817), .Y(
        n847) );
  AOI22X1 U247 ( .A0(n901), .A1(n843), .B0(n898), .B1(n842), .Y(n844) );
  AOI22X1 U248 ( .A0(n533), .A1(n669), .B0(n668), .B1(n897), .Y(n670) );
  OAI221XL U249 ( .A0(n862), .A1(n551), .B0(n545), .B1(n663), .C0(n662), .Y(
        n669) );
  OAI221XL U250 ( .A0(n882), .A1(n545), .B0(n542), .B1(n742), .C0(n667), .Y(
        n668) );
  AOI21X1 U251 ( .A0(n890), .A1(n556), .B0(n661), .Y(n662) );
  AOI22X1 U252 ( .A0(n575), .A1(n897), .B0(n533), .B1(n574), .Y(n581) );
  OAI221XL U253 ( .A0(n536), .A1(n757), .B0(n637), .B1(n545), .C0(n572), .Y(
        n575) );
  OAI211X1 U254 ( .A0(n835), .A1(n550), .B0(n736), .C0(n573), .Y(n574) );
  AOI2BB2X1 U255 ( .B0(n539), .B1(n727), .A0N(n550), .A1N(n744), .Y(n572) );
  OAI22X1 U256 ( .A0(n634), .A1(n813), .B0(n633), .B1(n767), .Y(n640) );
  AOI221XL U257 ( .A0(n549), .A1(n740), .B0(n799), .B1(n850), .C0(n632), .Y(
        n633) );
  AOI221XL U258 ( .A0(n867), .A1(n916), .B0(n547), .B1(n713), .C0(n630), .Y(
        n634) );
  OAI32X1 U259 ( .A0(n738), .A1(n860), .A2(n850), .B0(n631), .B1(n904), .Y(
        n632) );
  OAI22X1 U260 ( .A0(n770), .A1(n769), .B0(n768), .B1(n767), .Y(n771) );
  AOI211X1 U261 ( .A0(n881), .A1(n850), .B0(n766), .C0(n907), .Y(n768) );
  AOI221XL U262 ( .A0(n862), .A1(n552), .B0(n547), .B1(n776), .C0(n764), .Y(
        n770) );
  OAI22X1 U263 ( .A0(n541), .A1(n852), .B0(n886), .B1(n550), .Y(n766) );
  OAI22X1 U264 ( .A0(n816), .A1(n815), .B0(n814), .B1(n813), .Y(n817) );
  AOI221XL U265 ( .A0(n549), .A1(n812), .B0(n876), .B1(n540), .C0(n811), .Y(
        n814) );
  AOI221X1 U266 ( .A0(n556), .A1(n808), .B0(n552), .B1(n807), .C0(n806), .Y(
        n816) );
  OAI221XL U267 ( .A0(n536), .A1(n810), .B0(n879), .B1(n551), .C0(n809), .Y(
        n811) );
  AOI211X1 U268 ( .A0(n868), .A1(n556), .B0(n652), .C0(n651), .Y(n653) );
  AOI31X1 U269 ( .A0(n809), .A1(n717), .A2(n650), .B0(n533), .Y(n651) );
  OAI22X1 U270 ( .A0(n857), .A1(n803), .B0(n649), .B1(n897), .Y(n652) );
  AOI2BB2X1 U271 ( .B0(n853), .B1(n552), .A0N(n833), .A1N(n545), .Y(n650) );
  AOI2BB2X1 U272 ( .B0(n659), .B1(n897), .A0N(n897), .A1N(n658), .Y(n671) );
  OAI221XL U273 ( .A0(n877), .A1(n551), .B0(n545), .B1(n807), .C0(n656), .Y(
        n659) );
  AOI221XL U274 ( .A0(n548), .A1(n676), .B0(n711), .B1(n540), .C0(n657), .Y(
        n658) );
  AOI22X1 U275 ( .A0(n539), .A1(n765), .B0(n873), .B1(n903), .Y(n656) );
  AOI22X1 U276 ( .A0(n534), .A1(n610), .B0(n609), .B1(n902), .Y(n611) );
  OAI221XL U277 ( .A0(n595), .A1(n767), .B0(n594), .B1(n769), .C0(n593), .Y(
        n610) );
  OAI221XL U278 ( .A0(n608), .A1(n767), .B0(n607), .B1(n769), .C0(n606), .Y(
        n609) );
  AOI22X1 U279 ( .A0(n752), .A1(n902), .B0(n534), .B1(n751), .Y(n753) );
  OAI221XL U281 ( .A0(n750), .A1(n815), .B0(n749), .B1(n769), .C0(n748), .Y(
        n751) );
  OAI221XL U282 ( .A0(n732), .A1(n769), .B0(n731), .B1(n767), .C0(n730), .Y(
        n752) );
  AOI22X1 U283 ( .A0(n552), .A1(n532), .B0(n539), .B1(n857), .Y(n631) );
  AOI22X1 U284 ( .A0(n533), .A1(n562), .B0(n561), .B1(n897), .Y(n571) );
  OAI221XL U285 ( .A0(n880), .A1(n545), .B0(n542), .B1(n889), .C0(n558), .Y(
        n562) );
  OAI221XL U286 ( .A0(n532), .A1(n803), .B0(n722), .B1(n551), .C0(n560), .Y(
        n561) );
  INVX1 U287 ( .A(n663), .Y(n880) );
  AOI22X1 U288 ( .A0(n901), .A1(n605), .B0(n900), .B1(n604), .Y(n606) );
  OAI21XL U289 ( .A0(n602), .A1(n536), .B0(n601), .Y(n605) );
  OAI221XL U290 ( .A0(n551), .A1(n810), .B0(n835), .B1(n545), .C0(n603), .Y(
        n604) );
  AOI31X1 U291 ( .A0(n538), .A1(n742), .A2(n600), .B0(n910), .Y(n601) );
  CLKINVX3 U292 ( .A(n532), .Y(n852) );
  OAI21XL U293 ( .A0(n545), .A1(n537), .B0(n803), .Y(n647) );
  NAND2X1 U294 ( .A(n860), .B(n531), .Y(n755) );
  AOI21X1 U295 ( .A0(n699), .A1(n680), .B0(n545), .Y(n628) );
  INVX1 U296 ( .A(n531), .Y(n849) );
  OAI21XL U297 ( .A0(n850), .A1(n622), .B0(n550), .Y(n600) );
  OAI21XL U298 ( .A0(n850), .A1(n680), .B0(n550), .Y(n678) );
  OAI21XL U299 ( .A0(n536), .A1(n805), .B0(n763), .Y(n764) );
  AOI31X1 U300 ( .A0(n812), .A1(n903), .A2(n762), .B0(n915), .Y(n763) );
  INVX1 U301 ( .A(n761), .Y(n915) );
  AOI211X1 U302 ( .A0(n884), .A1(n540), .B0(n648), .C0(n647), .Y(n649) );
  OAI222X1 U303 ( .A0(n551), .A1(n807), .B0(n850), .B1(n693), .C0(n545), .C1(
        n821), .Y(n648) );
  NAND2X1 U304 ( .A(n861), .B(n554), .Y(n636) );
  OAI21X2 U305 ( .A0(n534), .A1(n792), .B0(n791), .Y(d[6]) );
  OAI2BB1X1 U306 ( .A0N(n790), .A1N(n789), .B0(n534), .Y(n791) );
  AOI221X1 U307 ( .A0(n900), .A1(n773), .B0(n901), .B1(n772), .C0(n771), .Y(
        n792) );
  AOI22X1 U308 ( .A0(n900), .A1(n788), .B0(n898), .B1(n787), .Y(n789) );
  NOR2BX1 U309 ( .AN(n660), .B(n876), .Y(n722) );
  BUFX3 U310 ( .A(n841), .Y(n536) );
  NAND2X1 U311 ( .A(n850), .B(n903), .Y(n841) );
  OAI221XL U312 ( .A0(n531), .A1(n664), .B0(n543), .B1(n709), .C0(n636), .Y(
        n630) );
  BUFX3 U313 ( .A(n784), .Y(n538) );
  NAND2X1 U314 ( .A(n531), .B(n537), .Y(n784) );
  AOI211X1 U315 ( .A0(n540), .A1(n852), .B0(n585), .C0(n647), .Y(n595) );
  OAI222X1 U316 ( .A0(n551), .A1(n756), .B0(n584), .B1(n536), .C0(n545), .C1(
        n889), .Y(n585) );
  AOI21X1 U317 ( .A0(n537), .A1(n535), .B0(n858), .Y(n584) );
  AOI211X1 U318 ( .A0(n533), .A1(n569), .B0(n848), .C0(n568), .Y(n570) );
  OAI221XL U319 ( .A0(n545), .A1(n807), .B0(n602), .B1(n541), .C0(n564), .Y(
        n569) );
  AOI21X1 U320 ( .A0(n567), .A1(n566), .B0(n533), .Y(n568) );
  AOI31X1 U321 ( .A0(n556), .A1(n565), .A2(n884), .B0(n563), .Y(n564) );
  INVX1 U322 ( .A(n830), .Y(n546) );
  INVX1 U323 ( .A(n840), .Y(n554) );
  INVX1 U324 ( .A(n840), .Y(n555) );
  INVX1 U325 ( .A(n544), .Y(n541) );
  INVX1 U326 ( .A(n829), .Y(n544) );
  AOI22X1 U327 ( .A0(n533), .A1(n646), .B0(n645), .B1(n897), .Y(n654) );
  OAI222X1 U328 ( .A0(n545), .A1(n782), .B0(n551), .B1(n660), .C0(n894), .C1(
        n541), .Y(n646) );
  OAI221XL U329 ( .A0(n892), .A1(n536), .B0(n551), .B1(n819), .C0(n644), .Y(
        n645) );
  AOI2BB2X1 U330 ( .B0(n835), .B1(n539), .A0N(n545), .A1N(n726), .Y(n644) );
  NAND2X1 U331 ( .A(n699), .B(n622), .Y(n775) );
  NOR2BX1 U332 ( .AN(n660), .B(n862), .Y(n602) );
  AOI21X1 U333 ( .A0(n690), .A1(n758), .B0(n903), .Y(n661) );
  AOI22X1 U334 ( .A0(n900), .A1(n747), .B0(n899), .B1(n746), .Y(n748) );
  OAI221XL U335 ( .A0(n860), .A1(n545), .B0(n542), .B1(n807), .C0(n745), .Y(
        n746) );
  OAI221XL U336 ( .A0(n885), .A1(n536), .B0(n545), .B1(n740), .C0(n739), .Y(
        n747) );
  AOI21X1 U337 ( .A0(n744), .A1(n552), .B0(n743), .Y(n745) );
  AOI22X1 U338 ( .A0(n556), .A1(n857), .B0(n539), .B1(n776), .Y(n777) );
  AOI22X1 U339 ( .A0(n548), .A1(n838), .B0(n882), .B1(n539), .Y(n839) );
  AOI31X1 U340 ( .A0(n703), .A1(n793), .A2(n702), .B0(n815), .Y(n704) );
  OAI2BB1X1 U341 ( .A0N(n700), .A1N(n699), .B0(n553), .Y(n703) );
  AOI22X1 U342 ( .A0(n894), .A1(n556), .B0(n701), .B1(n547), .Y(n702) );
  NAND2X1 U343 ( .A(n699), .B(n805), .Y(n715) );
  NAND2X1 U344 ( .A(n660), .B(n586), .Y(n756) );
  AOI21X1 U345 ( .A0(n660), .A1(n741), .B0(n545), .Y(n618) );
  AOI21X1 U346 ( .A0(n812), .A1(n538), .B0(n541), .Y(n720) );
  NAND2X1 U347 ( .A(n906), .B(n531), .Y(n717) );
  XNOR2X1 U348 ( .A(n903), .B(n531), .Y(n738) );
  NAND2X1 U349 ( .A(n539), .B(n537), .Y(n793) );
  XNOR2X1 U350 ( .A(n850), .B(n531), .Y(n762) );
  AOI21X1 U351 ( .A0(n833), .A1(n850), .B0(n556), .Y(n837) );
  AOI221X1 U352 ( .A0(n877), .A1(n540), .B0(n553), .B1(n735), .C0(n734), .Y(
        n750) );
  AOI21X1 U353 ( .A0(n536), .A1(n733), .B0(n799), .Y(n734) );
  OAI21XL U354 ( .A0(n861), .A1(n853), .B0(n850), .Y(n733) );
  AOI222X1 U355 ( .A0(n549), .A1(n713), .B0(n712), .B1(n711), .C0(n556), .C1(
        n537), .Y(n732) );
  OAI21XL U356 ( .A0(n850), .A1(n709), .B0(n550), .Y(n712) );
  AOI31X1 U357 ( .A0(n761), .A1(n624), .A2(n623), .B0(n767), .Y(n625) );
  AOI22X1 U358 ( .A0(n775), .A1(n850), .B0(n894), .B1(n553), .Y(n623) );
  INVX1 U359 ( .A(n830), .Y(n547) );
  INVX1 U360 ( .A(n830), .Y(n549) );
  INVX1 U361 ( .A(n830), .Y(n548) );
  XOR2X1 U362 ( .A(n533), .B(n531), .Y(n565) );
  INVX1 U363 ( .A(n840), .Y(n552) );
  INVX1 U364 ( .A(n840), .Y(n553) );
  NOR2BX1 U365 ( .AN(n830), .B(n554), .Y(n614) );
  OAI22X2 U366 ( .A0(n583), .A1(n902), .B0(n534), .B1(n582), .Y(d[0]) );
  AOI22X1 U367 ( .A0(n581), .A1(a[0]), .B0(n580), .B1(n579), .Y(n582) );
  AOI31X1 U368 ( .A0(n717), .A1(n848), .A2(n571), .B0(n570), .Y(n583) );
  AOI22X1 U369 ( .A0(n576), .A1(n897), .B0(n556), .B1(n833), .Y(n580) );
  AOI22X1 U370 ( .A0(n673), .A1(n902), .B0(n534), .B1(n672), .Y(n674) );
  OAI22X1 U371 ( .A0(a[0]), .A1(n654), .B0(n653), .B1(n848), .Y(n673) );
  OAI22X1 U372 ( .A0(a[0]), .A1(n671), .B0(n670), .B1(n848), .Y(n672) );
  OAI22X1 U373 ( .A0(n698), .A1(n767), .B0(n697), .B1(n769), .Y(n705) );
  AOI221X1 U374 ( .A0(n548), .A1(n693), .B0(n556), .B1(n797), .C0(n692), .Y(
        n698) );
  AOI222X1 U375 ( .A0(n759), .A1(n547), .B0(a[2]), .B1(n696), .C0(n556), .C1(
        n695), .Y(n697) );
  OAI22X1 U376 ( .A0(n888), .A1(n543), .B0(n550), .B1(n537), .Y(n692) );
  NOR2X1 U377 ( .A(n863), .B(n861), .Y(n804) );
  BUFX3 U378 ( .A(n710), .Y(n537) );
  NAND2X1 U379 ( .A(a[4]), .B(n852), .Y(n710) );
  AOI221X1 U380 ( .A0(n916), .A1(n785), .B0(n851), .B1(n666), .C0(n665), .Y(
        n667) );
  NOR3X1 U381 ( .A(n851), .B(a[7]), .C(n860), .Y(n665) );
  INVX1 U382 ( .A(n762), .Y(n851) );
  OAI21XL U383 ( .A0(n857), .A1(n550), .B0(n664), .Y(n666) );
  BUFX3 U384 ( .A(a[3]), .Y(n532) );
  AOI22X1 U385 ( .A0(n882), .A1(n850), .B0(a[2]), .B1(n612), .Y(n613) );
  CLKINVX3 U386 ( .A(a[0]), .Y(n848) );
  AOI211X1 U387 ( .A0(n724), .A1(n578), .B0(n577), .C0(a[0]), .Y(n579) );
  NAND2X1 U388 ( .A(n781), .B(n805), .Y(n578) );
  AOI21X1 U389 ( .A0(n803), .A1(n624), .B0(n897), .Y(n577) );
  BUFX3 U390 ( .A(a[5]), .Y(n533) );
  OAI221XL U391 ( .A0(n536), .A1(n808), .B0(n802), .B1(n545), .C0(n801), .Y(
        n818) );
  AOI22X1 U392 ( .A0(n539), .A1(n800), .B0(n799), .B1(a[2]), .Y(n801) );
  AOI33X1 U393 ( .A0(n532), .A1(n540), .A2(n904), .B0(n738), .B1(n742), .B2(
        a[2]), .Y(n739) );
  BUFX3 U394 ( .A(a[6]), .Y(n534) );
endmodule


module aes_cipher_top ( clk, rst, ld, done, key, text_in, text_out );
  input [127:0] key;
  input [127:0] text_in;
  output [127:0] text_out;
  input clk, rst, ld;
  output done;
  wire   N21, N32, N33, N34, N35, N36, N37, N38, N39, N48, N49, N50, N51, N52,
         N53, N54, N55, N64, N65, N66, N67, N68, N69, N70, N71, N80, N81, N82,
         N83, N84, N85, N86, N87, N96, N97, N98, N99, N100, N101, N102, N103,
         N112, N113, N114, N115, N116, N117, N118, N119, N128, N129, N130,
         N131, N132, N133, N134, N135, N144, N145, N146, N147, N148, N149,
         N150, N151, N160, N161, N162, N163, N164, N165, N166, N167, N176,
         N177, N178, N179, N180, N181, N182, N183, N192, N193, N194, N195,
         N196, N197, N198, N199, N208, N209, N210, N211, N212, N213, N214,
         N215, N224, N225, N226, N227, N228, N229, N230, N231, N240, N241,
         N242, N243, N244, N245, N246, N247, N256, N257, N258, N259, N260,
         N261, N262, N263, N272, N273, N274, N275, N276, N277, N278, N279,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463,
         N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474,
         N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, n6, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n727, n728, n729, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013;
  wire   [3:0] dcnt;
  wire   [31:0] w3;
  wire   [7:0] sa33;
  wire   [7:0] sa33_next;
  wire   [7:0] sa23;
  wire   [7:0] sa23_next;
  wire   [7:0] sa13;
  wire   [7:0] sa13_next;
  wire   [7:0] sa03;
  wire   [7:0] sa03_next;
  wire   [31:0] w2;
  wire   [7:0] sa32;
  wire   [7:0] sa32_next;
  wire   [7:0] sa22;
  wire   [7:0] sa22_next;
  wire   [7:0] sa12;
  wire   [7:0] sa12_next;
  wire   [7:0] sa02;
  wire   [7:0] sa02_next;
  wire   [31:0] w1;
  wire   [7:0] sa31;
  wire   [7:0] sa31_next;
  wire   [7:0] sa21;
  wire   [7:0] sa21_next;
  wire   [7:0] sa11;
  wire   [7:0] sa11_next;
  wire   [7:0] sa01;
  wire   [7:0] sa01_next;
  wire   [31:0] w0;
  wire   [7:0] sa30;
  wire   [7:0] sa30_next;
  wire   [7:0] sa20;
  wire   [7:0] sa20_next;
  wire   [7:0] sa10;
  wire   [7:0] sa10_next;
  wire   [7:0] sa00;
  wire   [7:0] sa00_next;
  wire   [7:0] sa00_sr;
  wire   [7:0] sa01_sr;
  wire   [7:0] sa02_sr;
  wire   [7:0] sa03_sr;
  wire   [7:0] sa10_sr;
  wire   [7:0] sa11_sr;
  wire   [7:0] sa12_sr;
  wire   [7:0] sa13_sr;
  wire   [7:0] sa20_sr;
  wire   [7:0] sa21_sr;
  wire   [7:0] sa22_sr;
  wire   [7:0] sa23_sr;
  wire   [7:0] sa30_sr;
  wire   [7:0] sa31_sr;
  wire   [7:0] sa32_sr;
  wire   [7:0] sa33_sr;

  aes_key_expand_128 u0 ( .clk(clk), .kld(n1009), .key(key), .wo_0(w0), .wo_1(
        w1), .wo_2(w2), .wo_3(w3) );
  aes_sbox_0 us00 ( .a(sa00), .d(sa00_sr) );
  aes_sbox_19 us01 ( .a(sa01), .d(sa01_sr) );
  aes_sbox_18 us02 ( .a(sa02), .d(sa02_sr) );
  aes_sbox_17 us03 ( .a(sa03), .d(sa03_sr) );
  aes_sbox_16 us10 ( .a(sa10), .d(sa13_sr) );
  aes_sbox_15 us11 ( .a(sa11), .d(sa10_sr) );
  aes_sbox_14 us12 ( .a(sa12), .d(sa11_sr) );
  aes_sbox_13 us13 ( .a(sa13), .d(sa12_sr) );
  aes_sbox_12 us20 ( .a(sa20), .d(sa22_sr) );
  aes_sbox_11 us21 ( .a(sa21), .d(sa23_sr) );
  aes_sbox_10 us22 ( .a(sa22), .d(sa20_sr) );
  aes_sbox_9 us23 ( .a(sa23), .d(sa21_sr) );
  aes_sbox_8 us30 ( .a(sa30), .d(sa31_sr) );
  aes_sbox_7 us31 ( .a(sa31), .d(sa32_sr) );
  aes_sbox_6 us32 ( .a(sa32), .d(sa33_sr) );
  aes_sbox_5 us33 ( .a(sa33), .d(sa30_sr) );
  EDFFX1 \text_in_r_reg[127]  ( .D(text_in[127]), .E(n1009), .CK(clk), .QN(
        n934) );
  EDFFX1 \text_in_r_reg[126]  ( .D(text_in[126]), .E(n1011), .CK(clk), .QN(
        n869) );
  EDFFX1 \text_in_r_reg[125]  ( .D(text_in[125]), .E(n1011), .CK(clk), .QN(
        n965) );
  EDFFX1 \text_in_r_reg[124]  ( .D(text_in[124]), .E(n1011), .CK(clk), .QN(
        n903) );
  EDFFX1 \text_in_r_reg[123]  ( .D(text_in[123]), .E(n1011), .CK(clk), .QN(
        n906) );
  EDFFX1 \text_in_r_reg[122]  ( .D(text_in[122]), .E(n1011), .CK(clk), .QN(
        n949) );
  EDFFX1 \text_in_r_reg[121]  ( .D(text_in[121]), .E(n1011), .CK(clk), .QN(
        n886) );
  EDFFX1 \text_in_r_reg[120]  ( .D(text_in[120]), .E(n1011), .CK(clk), .QN(
        n994) );
  EDFFX1 \text_in_r_reg[119]  ( .D(text_in[119]), .E(n1011), .CK(clk), .QN(
        n933) );
  EDFFX1 \text_in_r_reg[118]  ( .D(text_in[118]), .E(n1011), .CK(clk), .QN(
        n868) );
  EDFFX1 \text_in_r_reg[117]  ( .D(text_in[117]), .E(n1011), .CK(clk), .QN(
        n964) );
  EDFFX1 \text_in_r_reg[116]  ( .D(text_in[116]), .E(n1011), .CK(clk), .QN(
        n902) );
  EDFFX1 \text_in_r_reg[115]  ( .D(text_in[115]), .E(n1011), .CK(clk), .QN(
        n905) );
  EDFFX1 \text_in_r_reg[114]  ( .D(text_in[114]), .E(n1011), .CK(clk), .QN(
        n948) );
  EDFFX1 \text_in_r_reg[113]  ( .D(text_in[113]), .E(n1011), .CK(clk), .QN(
        n885) );
  EDFFX1 \text_in_r_reg[112]  ( .D(text_in[112]), .E(n1011), .CK(clk), .QN(
        n987) );
  EDFFX1 \text_in_r_reg[111]  ( .D(text_in[111]), .E(n1011), .CK(clk), .QN(
        n946) );
  EDFFX1 \text_in_r_reg[110]  ( .D(text_in[110]), .E(n1011), .CK(clk), .QN(
        n870) );
  EDFFX1 \text_in_r_reg[109]  ( .D(text_in[109]), .E(n1011), .CK(clk), .QN(
        n966) );
  EDFFX1 \text_in_r_reg[108]  ( .D(text_in[108]), .E(n1011), .CK(clk), .QN(
        n900) );
  EDFFX1 \text_in_r_reg[107]  ( .D(text_in[107]), .E(n1011), .CK(clk), .QN(
        n899) );
  EDFFX1 \text_in_r_reg[106]  ( .D(text_in[106]), .E(n1011), .CK(clk), .QN(
        n950) );
  EDFFX1 \text_in_r_reg[105]  ( .D(text_in[105]), .E(n1011), .CK(clk), .QN(
        n883) );
  EDFFX1 \text_in_r_reg[104]  ( .D(text_in[104]), .E(n1011), .CK(clk), .QN(
        n979) );
  EDFFX1 \text_in_r_reg[103]  ( .D(text_in[103]), .E(n1011), .CK(clk), .QN(
        n932) );
  EDFFX1 \text_in_r_reg[102]  ( .D(text_in[102]), .E(n1011), .CK(clk), .QN(
        n867) );
  EDFFX1 \text_in_r_reg[101]  ( .D(text_in[101]), .E(n1011), .CK(clk), .QN(
        n963) );
  EDFFX1 \text_in_r_reg[100]  ( .D(text_in[100]), .E(n1011), .CK(clk), .QN(
        n901) );
  EDFFX1 \text_in_r_reg[99]  ( .D(text_in[99]), .E(n1011), .CK(clk), .QN(n904)
         );
  EDFFX1 \text_in_r_reg[98]  ( .D(text_in[98]), .E(n1011), .CK(clk), .QN(n947)
         );
  EDFFX1 \text_in_r_reg[97]  ( .D(text_in[97]), .E(n1011), .CK(clk), .QN(n884)
         );
  EDFFX1 \text_in_r_reg[96]  ( .D(text_in[96]), .E(n1011), .CK(clk), .QN(n993)
         );
  EDFFX1 \text_in_r_reg[95]  ( .D(text_in[95]), .E(n1011), .CK(clk), .QN(n944)
         );
  EDFFX1 \text_in_r_reg[94]  ( .D(text_in[94]), .E(n1011), .CK(clk), .QN(n882)
         );
  EDFFX1 \text_in_r_reg[93]  ( .D(text_in[93]), .E(n1011), .CK(clk), .QN(n978)
         );
  EDFFX1 \text_in_r_reg[92]  ( .D(text_in[92]), .E(n1011), .CK(clk), .QN(n926)
         );
  EDFFX1 \text_in_r_reg[91]  ( .D(text_in[91]), .E(n1011), .CK(clk), .QN(n925)
         );
  EDFFX1 \text_in_r_reg[90]  ( .D(text_in[90]), .E(n1011), .CK(clk), .QN(n962)
         );
  EDFFX1 \text_in_r_reg[89]  ( .D(text_in[89]), .E(n1011), .CK(clk), .QN(n896)
         );
  EDFFX1 \text_in_r_reg[88]  ( .D(text_in[88]), .E(n1010), .CK(clk), .QN(n986)
         );
  EDFFX1 \text_in_r_reg[87]  ( .D(text_in[87]), .E(n1010), .CK(clk), .QN(n942)
         );
  EDFFX1 \text_in_r_reg[86]  ( .D(text_in[86]), .E(n1010), .CK(clk), .QN(n879)
         );
  EDFFX1 \text_in_r_reg[85]  ( .D(text_in[85]), .E(n1010), .CK(clk), .QN(n975)
         );
  EDFFX1 \text_in_r_reg[84]  ( .D(text_in[84]), .E(n1010), .CK(clk), .QN(n927)
         );
  EDFFX1 \text_in_r_reg[83]  ( .D(text_in[83]), .E(n1010), .CK(clk), .QN(n929)
         );
  EDFFX1 \text_in_r_reg[82]  ( .D(text_in[82]), .E(n1010), .CK(clk), .QN(n959)
         );
  EDFFX1 \text_in_r_reg[81]  ( .D(text_in[81]), .E(n1010), .CK(clk), .QN(n897)
         );
  EDFFX1 \text_in_r_reg[80]  ( .D(text_in[80]), .E(n1010), .CK(clk), .QN(n988)
         );
  EDFFX1 \text_in_r_reg[79]  ( .D(text_in[79]), .E(n1010), .CK(clk), .QN(n943)
         );
  EDFFX1 \text_in_r_reg[78]  ( .D(text_in[78]), .E(n1010), .CK(clk), .QN(n881)
         );
  EDFFX1 \text_in_r_reg[77]  ( .D(text_in[77]), .E(n1010), .CK(clk), .QN(n977)
         );
  EDFFX1 \text_in_r_reg[76]  ( .D(text_in[76]), .E(n1010), .CK(clk), .QN(n924)
         );
  EDFFX1 \text_in_r_reg[75]  ( .D(text_in[75]), .E(n1010), .CK(clk), .QN(n923)
         );
  EDFFX1 \text_in_r_reg[74]  ( .D(text_in[74]), .E(n1010), .CK(clk), .QN(n961)
         );
  EDFFX1 \text_in_r_reg[73]  ( .D(text_in[73]), .E(n1010), .CK(clk), .QN(n895)
         );
  EDFFX1 \text_in_r_reg[72]  ( .D(text_in[72]), .E(n1010), .CK(clk), .QN(n985)
         );
  EDFFX1 \text_in_r_reg[71]  ( .D(text_in[71]), .E(n1010), .CK(clk), .QN(n939)
         );
  EDFFX1 \text_in_r_reg[70]  ( .D(text_in[70]), .E(n1010), .CK(clk), .QN(n880)
         );
  EDFFX1 \text_in_r_reg[69]  ( .D(text_in[69]), .E(n1010), .CK(clk), .QN(n976)
         );
  EDFFX1 \text_in_r_reg[68]  ( .D(text_in[68]), .E(n1010), .CK(clk), .QN(n928)
         );
  EDFFX1 \text_in_r_reg[67]  ( .D(text_in[67]), .E(n1010), .CK(clk), .QN(n930)
         );
  EDFFX1 \text_in_r_reg[66]  ( .D(text_in[66]), .E(n1010), .CK(clk), .QN(n960)
         );
  EDFFX1 \text_in_r_reg[65]  ( .D(text_in[65]), .E(n1010), .CK(clk), .QN(n898)
         );
  EDFFX1 \text_in_r_reg[64]  ( .D(text_in[64]), .E(n1010), .CK(clk), .QN(n992)
         );
  EDFFX1 \text_in_r_reg[63]  ( .D(text_in[63]), .E(n1010), .CK(clk), .QN(n937)
         );
  EDFFX1 \text_in_r_reg[62]  ( .D(text_in[62]), .E(n1010), .CK(clk), .QN(n874)
         );
  EDFFX1 \text_in_r_reg[61]  ( .D(text_in[61]), .E(n1010), .CK(clk), .QN(n970)
         );
  EDFFX1 \text_in_r_reg[60]  ( .D(text_in[60]), .E(n1010), .CK(clk), .QN(n913)
         );
  EDFFX1 \text_in_r_reg[59]  ( .D(text_in[59]), .E(n1010), .CK(clk), .QN(n914)
         );
  EDFFX1 \text_in_r_reg[58]  ( .D(text_in[58]), .E(n1010), .CK(clk), .QN(n954)
         );
  EDFFX1 \text_in_r_reg[57]  ( .D(text_in[57]), .E(n1010), .CK(clk), .QN(n890)
         );
  EDFFX1 \text_in_r_reg[56]  ( .D(text_in[56]), .E(n1010), .CK(clk), .QN(n981)
         );
  EDFFX1 \text_in_r_reg[55]  ( .D(text_in[55]), .E(n1010), .CK(clk), .QN(n936)
         );
  EDFFX1 \text_in_r_reg[54]  ( .D(text_in[54]), .E(n1010), .CK(clk), .QN(n871)
         );
  EDFFX1 \text_in_r_reg[53]  ( .D(text_in[53]), .E(n1010), .CK(clk), .QN(n967)
         );
  EDFFX1 \text_in_r_reg[52]  ( .D(text_in[52]), .E(n1010), .CK(clk), .QN(n907)
         );
  EDFFX1 \text_in_r_reg[51]  ( .D(text_in[51]), .E(n1010), .CK(clk), .QN(n910)
         );
  EDFFX1 \text_in_r_reg[50]  ( .D(text_in[50]), .E(n1010), .CK(clk), .QN(n951)
         );
  EDFFX1 \text_in_r_reg[49]  ( .D(text_in[49]), .E(n1010), .CK(clk), .QN(n887)
         );
  EDFFX1 \text_in_r_reg[48]  ( .D(text_in[48]), .E(n1010), .CK(clk), .QN(n989)
         );
  EDFFX1 \text_in_r_reg[47]  ( .D(text_in[47]), .E(n1010), .CK(clk), .QN(n935)
         );
  EDFFX1 \text_in_r_reg[46]  ( .D(text_in[46]), .E(n1010), .CK(clk), .QN(n873)
         );
  EDFFX1 \text_in_r_reg[45]  ( .D(text_in[45]), .E(n1010), .CK(clk), .QN(n969)
         );
  EDFFX1 \text_in_r_reg[44]  ( .D(text_in[44]), .E(n1010), .CK(clk), .QN(n909)
         );
  EDFFX1 \text_in_r_reg[43]  ( .D(text_in[43]), .E(n1010), .CK(clk), .QN(n912)
         );
  EDFFX1 \text_in_r_reg[42]  ( .D(text_in[42]), .E(n1010), .CK(clk), .QN(n953)
         );
  EDFFX1 \text_in_r_reg[41]  ( .D(text_in[41]), .E(n1010), .CK(clk), .QN(n889)
         );
  EDFFX1 \text_in_r_reg[40]  ( .D(text_in[40]), .E(n1009), .CK(clk), .QN(n980)
         );
  EDFFX1 \text_in_r_reg[39]  ( .D(text_in[39]), .E(n1009), .CK(clk), .QN(n931)
         );
  EDFFX1 \text_in_r_reg[38]  ( .D(text_in[38]), .E(n1009), .CK(clk), .QN(n872)
         );
  EDFFX1 \text_in_r_reg[37]  ( .D(text_in[37]), .E(n1009), .CK(clk), .QN(n968)
         );
  EDFFX1 \text_in_r_reg[36]  ( .D(text_in[36]), .E(n1009), .CK(clk), .QN(n908)
         );
  EDFFX1 \text_in_r_reg[35]  ( .D(text_in[35]), .E(n1009), .CK(clk), .QN(n911)
         );
  EDFFX1 \text_in_r_reg[34]  ( .D(text_in[34]), .E(n1009), .CK(clk), .QN(n952)
         );
  EDFFX1 \text_in_r_reg[33]  ( .D(text_in[33]), .E(n1009), .CK(clk), .QN(n888)
         );
  EDFFX1 \text_in_r_reg[32]  ( .D(text_in[32]), .E(n1009), .CK(clk), .QN(n991)
         );
  EDFFX1 \text_in_r_reg[31]  ( .D(text_in[31]), .E(n1009), .CK(clk), .QN(n941)
         );
  EDFFX1 \text_in_r_reg[30]  ( .D(text_in[30]), .E(n1009), .CK(clk), .QN(n878)
         );
  EDFFX1 \text_in_r_reg[29]  ( .D(text_in[29]), .E(n1010), .CK(clk), .QN(n974)
         );
  EDFFX1 \text_in_r_reg[28]  ( .D(text_in[28]), .E(n1009), .CK(clk), .QN(n921)
         );
  EDFFX1 \text_in_r_reg[27]  ( .D(text_in[27]), .E(n1009), .CK(clk), .QN(n922)
         );
  EDFFX1 \text_in_r_reg[26]  ( .D(text_in[26]), .E(n1009), .CK(clk), .QN(n958)
         );
  EDFFX1 \text_in_r_reg[25]  ( .D(text_in[25]), .E(n1009), .CK(clk), .QN(n894)
         );
  EDFFX1 \text_in_r_reg[24]  ( .D(text_in[24]), .E(n1009), .CK(clk), .QN(n984)
         );
  EDFFX1 \text_in_r_reg[23]  ( .D(text_in[23]), .E(n1009), .CK(clk), .QN(n940)
         );
  EDFFX1 \text_in_r_reg[22]  ( .D(text_in[22]), .E(n1009), .CK(clk), .QN(n875)
         );
  EDFFX1 \text_in_r_reg[21]  ( .D(text_in[21]), .E(n1009), .CK(clk), .QN(n971)
         );
  EDFFX1 \text_in_r_reg[20]  ( .D(text_in[20]), .E(n1009), .CK(clk), .QN(n916)
         );
  EDFFX1 \text_in_r_reg[19]  ( .D(text_in[19]), .E(n1009), .CK(clk), .QN(n915)
         );
  EDFFX1 \text_in_r_reg[18]  ( .D(text_in[18]), .E(n1009), .CK(clk), .QN(n955)
         );
  EDFFX1 \text_in_r_reg[17]  ( .D(text_in[17]), .E(n1009), .CK(clk), .QN(n891)
         );
  EDFFX1 \text_in_r_reg[16]  ( .D(text_in[16]), .E(n1009), .CK(clk), .QN(n982)
         );
  EDFFX1 \text_in_r_reg[15]  ( .D(text_in[15]), .E(n1009), .CK(clk), .QN(n945)
         );
  EDFFX1 \text_in_r_reg[14]  ( .D(text_in[14]), .E(n1009), .CK(clk), .QN(n877)
         );
  EDFFX1 \text_in_r_reg[13]  ( .D(text_in[13]), .E(n1009), .CK(clk), .QN(n973)
         );
  EDFFX1 \text_in_r_reg[12]  ( .D(text_in[12]), .E(n1009), .CK(clk), .QN(n918)
         );
  EDFFX1 \text_in_r_reg[11]  ( .D(text_in[11]), .E(n1009), .CK(clk), .QN(n917)
         );
  EDFFX1 \text_in_r_reg[10]  ( .D(text_in[10]), .E(n1009), .CK(clk), .QN(n957)
         );
  EDFFX1 \text_in_r_reg[9]  ( .D(text_in[9]), .E(n1009), .CK(clk), .QN(n892)
         );
  EDFFX1 \text_in_r_reg[8]  ( .D(text_in[8]), .E(n1009), .CK(clk), .QN(n983)
         );
  EDFFX1 \text_in_r_reg[7]  ( .D(text_in[7]), .E(n1009), .CK(clk), .QN(n938)
         );
  EDFFX1 \text_in_r_reg[6]  ( .D(text_in[6]), .E(n1009), .CK(clk), .QN(n876)
         );
  EDFFX1 \text_in_r_reg[5]  ( .D(text_in[5]), .E(n1009), .CK(clk), .QN(n972)
         );
  EDFFX1 \text_in_r_reg[4]  ( .D(text_in[4]), .E(n1009), .CK(clk), .QN(n919)
         );
  EDFFX1 \text_in_r_reg[3]  ( .D(text_in[3]), .E(n1009), .CK(clk), .QN(n920)
         );
  EDFFX1 \text_in_r_reg[2]  ( .D(text_in[2]), .E(n1009), .CK(clk), .QN(n956)
         );
  EDFFX1 \text_in_r_reg[1]  ( .D(text_in[1]), .E(n1009), .CK(clk), .QN(n893)
         );
  EDFFX1 \text_in_r_reg[0]  ( .D(text_in[0]), .E(n1009), .CK(clk), .QN(n990)
         );
  DFFHQX1 \dcnt_reg[3]  ( .D(n995), .CK(clk), .Q(dcnt[3]) );
  DFFHQX1 \dcnt_reg[1]  ( .D(n146), .CK(clk), .Q(dcnt[1]) );
  DFFHQX1 \dcnt_reg[0]  ( .D(n147), .CK(clk), .Q(dcnt[0]) );
  DFFX1 ld_r_reg ( .D(n1011), .CK(clk), .Q(n996), .QN(n6) );
  DFFHQX1 \sa01_reg[6]  ( .D(N214), .CK(clk), .Q(sa01[6]) );
  DFFHQX1 \sa21_reg[6]  ( .D(N182), .CK(clk), .Q(sa21[6]) );
  DFFHQX1 \sa31_reg[6]  ( .D(N166), .CK(clk), .Q(sa31[6]) );
  DFFHQX1 \sa11_reg[6]  ( .D(N198), .CK(clk), .Q(sa11[6]) );
  DFFHQX1 \sa03_reg[6]  ( .D(N86), .CK(clk), .Q(sa03[6]) );
  DFFHQX1 \sa23_reg[6]  ( .D(N54), .CK(clk), .Q(sa23[6]) );
  DFFHQX1 \sa33_reg[6]  ( .D(N38), .CK(clk), .Q(sa33[6]) );
  DFFHQX1 \sa13_reg[6]  ( .D(N70), .CK(clk), .Q(sa13[6]) );
  DFFHQX1 \sa02_reg[6]  ( .D(N150), .CK(clk), .Q(sa02[6]) );
  DFFHQX1 \sa22_reg[6]  ( .D(N118), .CK(clk), .Q(sa22[6]) );
  DFFHQX1 \sa32_reg[6]  ( .D(N102), .CK(clk), .Q(sa32[6]) );
  DFFHQX1 \sa12_reg[6]  ( .D(N134), .CK(clk), .Q(sa12[6]) );
  DFFHQX1 \sa20_reg[6]  ( .D(N246), .CK(clk), .Q(sa20[6]) );
  DFFHQX1 \sa00_reg[6]  ( .D(N278), .CK(clk), .Q(sa00[6]) );
  DFFHQX1 \sa10_reg[6]  ( .D(N262), .CK(clk), .Q(sa10[6]) );
  DFFHQX1 \sa30_reg[6]  ( .D(N230), .CK(clk), .Q(sa30[6]) );
  DFFHQX1 \sa01_reg[5]  ( .D(N213), .CK(clk), .Q(sa01[5]) );
  DFFHQX1 \sa21_reg[5]  ( .D(N181), .CK(clk), .Q(sa21[5]) );
  DFFHQX1 \sa31_reg[5]  ( .D(N165), .CK(clk), .Q(sa31[5]) );
  DFFHQX1 \sa11_reg[5]  ( .D(N197), .CK(clk), .Q(sa11[5]) );
  DFFHQX1 \sa03_reg[5]  ( .D(N85), .CK(clk), .Q(sa03[5]) );
  DFFHQX1 \sa23_reg[5]  ( .D(N53), .CK(clk), .Q(sa23[5]) );
  DFFHQX1 \sa33_reg[5]  ( .D(N37), .CK(clk), .Q(sa33[5]) );
  DFFHQX1 \sa13_reg[5]  ( .D(N69), .CK(clk), .Q(sa13[5]) );
  DFFHQX1 \sa02_reg[5]  ( .D(N149), .CK(clk), .Q(sa02[5]) );
  DFFHQX1 \sa22_reg[5]  ( .D(N117), .CK(clk), .Q(sa22[5]) );
  DFFHQX1 \sa32_reg[5]  ( .D(N101), .CK(clk), .Q(sa32[5]) );
  DFFHQX1 \sa12_reg[5]  ( .D(N133), .CK(clk), .Q(sa12[5]) );
  DFFHQX1 \sa20_reg[5]  ( .D(N245), .CK(clk), .Q(sa20[5]) );
  DFFHQX1 \sa00_reg[5]  ( .D(N277), .CK(clk), .Q(sa00[5]) );
  DFFHQX1 \sa10_reg[5]  ( .D(N261), .CK(clk), .Q(sa10[5]) );
  DFFHQX1 \sa30_reg[5]  ( .D(N229), .CK(clk), .Q(sa30[5]) );
  DFFHQX1 \sa31_reg[3]  ( .D(N163), .CK(clk), .Q(sa31[3]) );
  DFFHQX1 \sa11_reg[3]  ( .D(N195), .CK(clk), .Q(sa11[3]) );
  DFFHQX1 \sa01_reg[3]  ( .D(N211), .CK(clk), .Q(sa01[3]) );
  DFFHQX1 \sa21_reg[3]  ( .D(N179), .CK(clk), .Q(sa21[3]) );
  DFFHQX1 \sa03_reg[3]  ( .D(N83), .CK(clk), .Q(sa03[3]) );
  DFFHQX1 \sa33_reg[3]  ( .D(N35), .CK(clk), .Q(sa33[3]) );
  DFFHQX1 \sa23_reg[3]  ( .D(N51), .CK(clk), .Q(sa23[3]) );
  DFFHQX1 \sa13_reg[3]  ( .D(N67), .CK(clk), .Q(sa13[3]) );
  DFFHQX1 \sa02_reg[3]  ( .D(N147), .CK(clk), .Q(sa02[3]) );
  DFFHQX1 \sa22_reg[3]  ( .D(N115), .CK(clk), .Q(sa22[3]) );
  DFFHQX1 \sa32_reg[3]  ( .D(N99), .CK(clk), .Q(sa32[3]) );
  DFFHQX1 \sa12_reg[3]  ( .D(N131), .CK(clk), .Q(sa12[3]) );
  DFFHQX1 \sa00_reg[3]  ( .D(N275), .CK(clk), .Q(sa00[3]) );
  DFFHQX1 \sa10_reg[3]  ( .D(N259), .CK(clk), .Q(sa10[3]) );
  DFFHQX1 \sa30_reg[3]  ( .D(N227), .CK(clk), .Q(sa30[3]) );
  DFFHQX1 \sa20_reg[3]  ( .D(N243), .CK(clk), .Q(sa20[3]) );
  DFFHQX1 \sa31_reg[1]  ( .D(N161), .CK(clk), .Q(sa31[1]) );
  DFFHQX1 \sa11_reg[1]  ( .D(N193), .CK(clk), .Q(sa11[1]) );
  DFFHQX1 \sa01_reg[1]  ( .D(N209), .CK(clk), .Q(sa01[1]) );
  DFFHQX1 \sa21_reg[1]  ( .D(N177), .CK(clk), .Q(sa21[1]) );
  DFFHQX1 \sa03_reg[1]  ( .D(N81), .CK(clk), .Q(sa03[1]) );
  DFFHQX1 \sa33_reg[1]  ( .D(N33), .CK(clk), .Q(sa33[1]) );
  DFFHQX1 \sa23_reg[1]  ( .D(N49), .CK(clk), .Q(sa23[1]) );
  DFFHQX1 \sa13_reg[1]  ( .D(N65), .CK(clk), .Q(sa13[1]) );
  DFFHQX1 \sa02_reg[1]  ( .D(N145), .CK(clk), .Q(sa02[1]) );
  DFFHQX1 \sa22_reg[1]  ( .D(N113), .CK(clk), .Q(sa22[1]) );
  DFFHQX1 \sa32_reg[1]  ( .D(N97), .CK(clk), .Q(sa32[1]) );
  DFFHQX1 \sa12_reg[1]  ( .D(N129), .CK(clk), .Q(sa12[1]) );
  DFFHQX1 \sa00_reg[1]  ( .D(N273), .CK(clk), .Q(sa00[1]) );
  DFFHQX1 \sa10_reg[1]  ( .D(N257), .CK(clk), .Q(sa10[1]) );
  DFFHQX1 \sa30_reg[1]  ( .D(N225), .CK(clk), .Q(sa30[1]) );
  DFFHQX1 \sa20_reg[1]  ( .D(N241), .CK(clk), .Q(sa20[1]) );
  DFFHQX1 \sa20_reg[7]  ( .D(N247), .CK(clk), .Q(sa20[7]) );
  DFFHQX1 \sa23_reg[7]  ( .D(N55), .CK(clk), .Q(sa23[7]) );
  DFFHQX1 \sa01_reg[7]  ( .D(N215), .CK(clk), .Q(sa01[7]) );
  DFFHQX1 \sa21_reg[7]  ( .D(N183), .CK(clk), .Q(sa21[7]) );
  DFFHQX1 \sa11_reg[7]  ( .D(N199), .CK(clk), .Q(sa11[7]) );
  DFFHQX1 \sa03_reg[7]  ( .D(N87), .CK(clk), .Q(sa03[7]) );
  DFFHQX1 \sa13_reg[7]  ( .D(N71), .CK(clk), .Q(sa13[7]) );
  DFFHQX1 \sa31_reg[7]  ( .D(N167), .CK(clk), .Q(sa31[7]) );
  DFFHQX1 \sa33_reg[7]  ( .D(N39), .CK(clk), .Q(sa33[7]) );
  DFFHQX1 \sa02_reg[7]  ( .D(N151), .CK(clk), .Q(sa02[7]) );
  DFFHQX1 \sa12_reg[7]  ( .D(N135), .CK(clk), .Q(sa12[7]) );
  DFFHQX1 \sa22_reg[7]  ( .D(N119), .CK(clk), .Q(sa22[7]) );
  DFFHQX1 \sa00_reg[7]  ( .D(N279), .CK(clk), .Q(sa00[7]) );
  DFFHQX1 \sa10_reg[7]  ( .D(N263), .CK(clk), .Q(sa10[7]) );
  DFFHQX1 \sa30_reg[7]  ( .D(N231), .CK(clk), .Q(sa30[7]) );
  DFFHQX1 \sa32_reg[7]  ( .D(N103), .CK(clk), .Q(sa32[7]) );
  XOR2XL U709 ( .A(sa21_sr[5]), .B(sa31_sr[4]), .Y(n309) );
  XOR2X1 U711 ( .A(n309), .B(n308), .Y(sa31_next[5]) );
  XOR2XL U569 ( .A(sa22_sr[5]), .B(sa32_sr[4]), .Y(n399) );
  XOR2X1 U571 ( .A(n399), .B(n398), .Y(sa32_next[5]) );
  XOR2XL U849 ( .A(sa20_sr[5]), .B(sa30_sr[4]), .Y(n219) );
  XOR2X1 U851 ( .A(n219), .B(n218), .Y(sa30_next[5]) );
  XOR2X1 U756 ( .A(sa11_sr[1]), .B(sa21_sr[1]), .Y(n275) );
  XOR2X1 U758 ( .A(n275), .B(n274), .Y(sa11_next[2]) );
  XOR2X1 U476 ( .A(sa13_sr[1]), .B(sa23_sr[1]), .Y(n455) );
  XOR2X1 U478 ( .A(n455), .B(n454), .Y(sa13_next[2]) );
  XOR2X1 U616 ( .A(sa12_sr[1]), .B(sa22_sr[1]), .Y(n365) );
  XOR2X1 U618 ( .A(n365), .B(n364), .Y(sa12_next[2]) );
  XOR2X1 U896 ( .A(sa10_sr[1]), .B(sa20_sr[1]), .Y(n185) );
  XOR2X1 U898 ( .A(n185), .B(n184), .Y(sa10_next[2]) );
  XOR2X1 U700 ( .A(n318), .B(n317), .Y(n315) );
  XOR2X1 U701 ( .A(n316), .B(n315), .Y(sa31_next[3]) );
  XOR2X1 U805 ( .A(n529), .B(n246), .Y(n244) );
  XOR2X1 U806 ( .A(n245), .B(n244), .Y(sa01_next[4]) );
  XOR2X1 U735 ( .A(n534), .B(n538), .Y(n290) );
  XOR2X1 U737 ( .A(n290), .B(n289), .Y(sa21_next[4]) );
  XOR2X1 U525 ( .A(n565), .B(n426), .Y(n424) );
  XOR2X1 U526 ( .A(n425), .B(n424), .Y(sa03_next[4]) );
  XOR2X1 U420 ( .A(n498), .B(n497), .Y(n495) );
  XOR2X1 U421 ( .A(n496), .B(n495), .Y(sa33_next[3]) );
  XOR2X1 U455 ( .A(n570), .B(n574), .Y(n470) );
  XOR2X1 U457 ( .A(n470), .B(n469), .Y(sa23_next[4]) );
  XOR2X1 U665 ( .A(n547), .B(n336), .Y(n334) );
  XOR2X1 U666 ( .A(n335), .B(n334), .Y(sa02_next[4]) );
  XOR2X1 U560 ( .A(n408), .B(n407), .Y(n405) );
  XOR2X1 U561 ( .A(n406), .B(n405), .Y(sa32_next[3]) );
  XOR2X1 U595 ( .A(n552), .B(n556), .Y(n380) );
  XOR2X1 U597 ( .A(n380), .B(n379), .Y(sa22_next[4]) );
  XOR2X1 U840 ( .A(n228), .B(n227), .Y(n225) );
  XOR2X1 U841 ( .A(n226), .B(n225), .Y(sa30_next[3]) );
  XOR2X1 U945 ( .A(n511), .B(n156), .Y(n154) );
  XOR2X1 U946 ( .A(n155), .B(n154), .Y(sa00_next[4]) );
  XOR2X1 U875 ( .A(n516), .B(n520), .Y(n200) );
  XOR2X1 U877 ( .A(n200), .B(n199), .Y(sa20_next[4]) );
  XOR2X1 U690 ( .A(n543), .B(n541), .Y(n323) );
  XOR2X1 U692 ( .A(n323), .B(n322), .Y(sa31_next[1]) );
  XOR2X1 U410 ( .A(n579), .B(n577), .Y(n503) );
  XOR2X1 U412 ( .A(n503), .B(n502), .Y(sa33_next[1]) );
  XOR2X1 U550 ( .A(n561), .B(n559), .Y(n413) );
  XOR2X1 U552 ( .A(n413), .B(n412), .Y(sa32_next[1]) );
  XOR2X1 U830 ( .A(n525), .B(n523), .Y(n233) );
  XOR2X1 U832 ( .A(n233), .B(n232), .Y(sa30_next[1]) );
  XOR2X1 U775 ( .A(sa11_sr[5]), .B(sa21_sr[5]), .Y(n261) );
  XOR2X1 U777 ( .A(n261), .B(n260), .Y(sa11_next[6]) );
  XOR2X1 U635 ( .A(sa12_sr[5]), .B(sa22_sr[5]), .Y(n351) );
  XOR2X1 U637 ( .A(n351), .B(n350), .Y(sa12_next[6]) );
  XOR2X1 U915 ( .A(sa10_sr[5]), .B(sa20_sr[5]), .Y(n171) );
  XOR2X1 U917 ( .A(n171), .B(n170), .Y(sa10_next[6]) );
  XOR2X1 U759 ( .A(w1[19]), .B(sa01_sr[3]), .Y(n273) );
  XOR2X1 U619 ( .A(w2[19]), .B(sa02_sr[3]), .Y(n363) );
  XOR2X1 U899 ( .A(w0[19]), .B(sa00_sr[3]), .Y(n183) );
  XOR2X1 U697 ( .A(w1[3]), .B(sa01_sr[2]), .Y(n318) );
  XOR2X1 U557 ( .A(w2[3]), .B(sa02_sr[2]), .Y(n408) );
  XOR2X1 U837 ( .A(w0[3]), .B(sa00_sr[2]), .Y(n228) );
  XOR2X1 U417 ( .A(w3[3]), .B(sa03_sr[2]), .Y(n498) );
  XOR2X1 U479 ( .A(w3[19]), .B(sa03_sr[3]), .Y(n453) );
  XOR2X1 U475 ( .A(w3[18]), .B(sa03_sr[2]), .Y(n456) );
  XOR2X1 U477 ( .A(n567), .B(n456), .Y(n454) );
  XOR2X1 U428 ( .A(w3[5]), .B(sa03_sr[4]), .Y(n490) );
  XOR2X1 U430 ( .A(n573), .B(n490), .Y(n488) );
  XOR2X1 U494 ( .A(w3[22]), .B(sa03_sr[6]), .Y(n442) );
  XOR2X1 U496 ( .A(n563), .B(n442), .Y(n440) );
  XOR2X1 U456 ( .A(n566), .B(n471), .Y(n469) );
  XOR2X1 U708 ( .A(w1[5]), .B(sa01_sr[4]), .Y(n310) );
  XOR2X1 U710 ( .A(n537), .B(n310), .Y(n308) );
  XOR2X1 U568 ( .A(w2[5]), .B(sa02_sr[4]), .Y(n400) );
  XOR2X1 U570 ( .A(n555), .B(n400), .Y(n398) );
  XOR2X1 U848 ( .A(w0[5]), .B(sa00_sr[4]), .Y(n220) );
  XOR2X1 U850 ( .A(n519), .B(n220), .Y(n218) );
  XOR2X1 U755 ( .A(w1[18]), .B(sa01_sr[2]), .Y(n276) );
  XOR2X1 U757 ( .A(n531), .B(n276), .Y(n274) );
  XOR2X1 U615 ( .A(w2[18]), .B(sa02_sr[2]), .Y(n366) );
  XOR2X1 U617 ( .A(n549), .B(n366), .Y(n364) );
  XOR2X1 U895 ( .A(w0[18]), .B(sa00_sr[2]), .Y(n186) );
  XOR2X1 U897 ( .A(n513), .B(n186), .Y(n184) );
  XOR2X1 U734 ( .A(w1[12]), .B(sa31_sr[4]), .Y(n291) );
  XOR2X1 U736 ( .A(n530), .B(n291), .Y(n289) );
  XOR2X1 U594 ( .A(w2[12]), .B(sa32_sr[4]), .Y(n381) );
  XOR2X1 U596 ( .A(n548), .B(n381), .Y(n379) );
  XOR2X1 U874 ( .A(w0[12]), .B(sa30_sr[4]), .Y(n201) );
  XOR2X1 U876 ( .A(n512), .B(n201), .Y(n199) );
  XOR2X1 U774 ( .A(w1[22]), .B(sa01_sr[6]), .Y(n262) );
  XOR2X1 U776 ( .A(n527), .B(n262), .Y(n260) );
  XOR2X1 U634 ( .A(w2[22]), .B(sa02_sr[6]), .Y(n352) );
  XOR2X1 U636 ( .A(n545), .B(n352), .Y(n350) );
  XOR2X1 U914 ( .A(w0[22]), .B(sa00_sr[6]), .Y(n172) );
  XOR2X1 U916 ( .A(n509), .B(n172), .Y(n170) );
  XOR2XL U689 ( .A(sa21_sr[1]), .B(sa31_sr[0]), .Y(n324) );
  XOR2X1 U688 ( .A(w1[1]), .B(sa01_sr[0]), .Y(n325) );
  XOR2X1 U691 ( .A(n325), .B(n324), .Y(n322) );
  XOR2XL U409 ( .A(sa23_sr[1]), .B(sa33_sr[0]), .Y(n504) );
  XOR2X1 U408 ( .A(w3[1]), .B(sa03_sr[0]), .Y(n505) );
  XOR2X1 U411 ( .A(n505), .B(n504), .Y(n502) );
  XOR2XL U549 ( .A(sa22_sr[1]), .B(sa32_sr[0]), .Y(n414) );
  XOR2X1 U548 ( .A(w2[1]), .B(sa02_sr[0]), .Y(n415) );
  XOR2X1 U551 ( .A(n415), .B(n414), .Y(n412) );
  XOR2XL U829 ( .A(sa20_sr[1]), .B(sa30_sr[0]), .Y(n234) );
  XOR2X1 U828 ( .A(w0[1]), .B(sa00_sr[0]), .Y(n235) );
  XOR2X1 U831 ( .A(n235), .B(n234), .Y(n232) );
  XOR2X1 U751 ( .A(sa11_sr[0]), .B(sa21_sr[0]), .Y(n279) );
  XOR2X1 U750 ( .A(w1[17]), .B(sa01_sr[1]), .Y(n280) );
  XOR2X1 U753 ( .A(n280), .B(n279), .Y(n277) );
  XOR2X1 U471 ( .A(sa13_sr[0]), .B(sa23_sr[0]), .Y(n459) );
  XOR2X1 U470 ( .A(w3[17]), .B(sa03_sr[1]), .Y(n460) );
  XOR2X1 U473 ( .A(n460), .B(n459), .Y(n457) );
  XOR2X1 U611 ( .A(sa12_sr[0]), .B(sa22_sr[0]), .Y(n369) );
  XOR2X1 U610 ( .A(w2[17]), .B(sa02_sr[1]), .Y(n370) );
  XOR2X1 U613 ( .A(n370), .B(n369), .Y(n367) );
  XOR2X1 U891 ( .A(sa10_sr[0]), .B(sa20_sr[0]), .Y(n189) );
  XOR2X1 U890 ( .A(w0[17]), .B(sa00_sr[1]), .Y(n190) );
  XOR2X1 U893 ( .A(n190), .B(n189), .Y(n187) );
  XOR2X1 U765 ( .A(sa11_sr[3]), .B(sa21_sr[3]), .Y(n268) );
  XOR2X1 U764 ( .A(w1[20]), .B(sa01_sr[4]), .Y(n269) );
  XOR2X1 U767 ( .A(n269), .B(n268), .Y(n266) );
  XOR2X1 U485 ( .A(sa13_sr[3]), .B(sa23_sr[3]), .Y(n448) );
  XOR2X1 U484 ( .A(w3[20]), .B(sa03_sr[4]), .Y(n449) );
  XOR2X1 U487 ( .A(n449), .B(n448), .Y(n446) );
  XOR2X1 U625 ( .A(sa12_sr[3]), .B(sa22_sr[3]), .Y(n358) );
  XOR2X1 U624 ( .A(w2[20]), .B(sa02_sr[4]), .Y(n359) );
  XOR2X1 U627 ( .A(n359), .B(n358), .Y(n356) );
  XOR2X1 U905 ( .A(sa10_sr[3]), .B(sa20_sr[3]), .Y(n178) );
  XOR2X1 U904 ( .A(w0[20]), .B(sa00_sr[4]), .Y(n179) );
  XOR2X1 U907 ( .A(n179), .B(n178), .Y(n176) );
  XOR2X1 U770 ( .A(w1[21]), .B(sa01_sr[5]), .Y(n265) );
  XOR2X1 U772 ( .A(n528), .B(n265), .Y(n263) );
  XOR2X1 U490 ( .A(w3[21]), .B(sa03_sr[5]), .Y(n445) );
  XOR2X1 U492 ( .A(n564), .B(n445), .Y(n443) );
  XOR2X1 U630 ( .A(w2[21]), .B(sa02_sr[5]), .Y(n355) );
  XOR2X1 U632 ( .A(n546), .B(n355), .Y(n353) );
  XOR2X1 U910 ( .A(w0[21]), .B(sa00_sr[5]), .Y(n175) );
  XOR2X1 U912 ( .A(n510), .B(n175), .Y(n173) );
  XOR2X1 U693 ( .A(w1[2]), .B(sa01_sr[1]), .Y(n321) );
  XOR2X1 U695 ( .A(n540), .B(n321), .Y(n319) );
  XOR2X1 U413 ( .A(w3[2]), .B(sa03_sr[1]), .Y(n501) );
  XOR2X1 U415 ( .A(n576), .B(n501), .Y(n499) );
  XOR2X1 U553 ( .A(w2[2]), .B(sa02_sr[1]), .Y(n411) );
  XOR2X1 U555 ( .A(n558), .B(n411), .Y(n409) );
  XOR2X1 U833 ( .A(w0[2]), .B(sa00_sr[1]), .Y(n231) );
  XOR2X1 U835 ( .A(n522), .B(n231), .Y(n229) );
  XOR2X1 U797 ( .A(w1[27]), .B(sa11_sr[3]), .Y(n249) );
  XOR2X1 U799 ( .A(n530), .B(n249), .Y(n247) );
  XOR2X1 U517 ( .A(w3[27]), .B(sa13_sr[3]), .Y(n429) );
  XOR2X1 U519 ( .A(n566), .B(n429), .Y(n427) );
  XOR2X1 U657 ( .A(w2[27]), .B(sa12_sr[3]), .Y(n339) );
  XOR2X1 U659 ( .A(n548), .B(n339), .Y(n337) );
  XOR2X1 U937 ( .A(w0[27]), .B(sa10_sr[3]), .Y(n159) );
  XOR2X1 U939 ( .A(n512), .B(n159), .Y(n157) );
  XOR2X1 U432 ( .A(w3[6]), .B(sa03_sr[5]), .Y(n487) );
  XOR2X1 U434 ( .A(n572), .B(n487), .Y(n485) );
  XOR2X1 U723 ( .A(w1[9]), .B(sa31_sr[1]), .Y(n299) );
  XOR2X1 U725 ( .A(n533), .B(n299), .Y(n297) );
  XOR2X1 U443 ( .A(w3[9]), .B(sa33_sr[1]), .Y(n479) );
  XOR2X1 U445 ( .A(n569), .B(n479), .Y(n477) );
  XOR2X1 U583 ( .A(w2[9]), .B(sa32_sr[1]), .Y(n389) );
  XOR2X1 U585 ( .A(n551), .B(n389), .Y(n387) );
  XOR2X1 U863 ( .A(w0[9]), .B(sa30_sr[1]), .Y(n209) );
  XOR2X1 U865 ( .A(n515), .B(n209), .Y(n207) );
  XOR2X1 U778 ( .A(w1[23]), .B(sa01_sr[7]), .Y(n259) );
  XOR2X1 U780 ( .A(n534), .B(n259), .Y(n257) );
  XOR2X1 U498 ( .A(w3[23]), .B(sa03_sr[7]), .Y(n439) );
  XOR2X1 U500 ( .A(n570), .B(n439), .Y(n437) );
  XOR2X1 U716 ( .A(w1[7]), .B(sa01_sr[6]), .Y(n304) );
  XOR2X1 U718 ( .A(n535), .B(n304), .Y(n302) );
  XOR2X1 U436 ( .A(w3[7]), .B(sa03_sr[6]), .Y(n484) );
  XOR2X1 U438 ( .A(n571), .B(n484), .Y(n482) );
  XOR2X1 U638 ( .A(w2[23]), .B(sa02_sr[7]), .Y(n349) );
  XOR2X1 U640 ( .A(n552), .B(n349), .Y(n347) );
  XOR2X1 U918 ( .A(w0[23]), .B(sa00_sr[7]), .Y(n169) );
  XOR2X1 U920 ( .A(n516), .B(n169), .Y(n167) );
  XOR2X1 U856 ( .A(w0[7]), .B(sa00_sr[6]), .Y(n214) );
  XOR2X1 U858 ( .A(n517), .B(n214), .Y(n212) );
  XOR2X1 U576 ( .A(w2[7]), .B(sa02_sr[6]), .Y(n394) );
  XOR2X1 U578 ( .A(n553), .B(n394), .Y(n392) );
  XOR2X1 U712 ( .A(w1[6]), .B(sa01_sr[5]), .Y(n307) );
  XOR2X1 U714 ( .A(n536), .B(n307), .Y(n305) );
  XOR2X1 U572 ( .A(w2[6]), .B(sa02_sr[5]), .Y(n397) );
  XOR2X1 U574 ( .A(n554), .B(n397), .Y(n395) );
  XOR2X1 U852 ( .A(w0[6]), .B(sa00_sr[5]), .Y(n217) );
  XOR2X1 U854 ( .A(n518), .B(n217), .Y(n215) );
  XOR2X1 U786 ( .A(w1[25]), .B(sa11_sr[1]), .Y(n254) );
  XOR2X1 U646 ( .A(w2[25]), .B(sa12_sr[1]), .Y(n344) );
  XOR2X1 U926 ( .A(w0[25]), .B(sa10_sr[1]), .Y(n164) );
  XOR2X1 U730 ( .A(w1[11]), .B(sa31_sr[3]), .Y(n294) );
  XOR2X1 U590 ( .A(w2[11]), .B(sa32_sr[3]), .Y(n384) );
  XOR2X1 U870 ( .A(w0[11]), .B(sa30_sr[3]), .Y(n204) );
  XOR2X1 U506 ( .A(w3[25]), .B(sa13_sr[1]), .Y(n434) );
  XOR2X1 U803 ( .A(w1[28]), .B(sa11_sr[4]), .Y(n246) );
  XOR2X1 U663 ( .A(w2[28]), .B(sa12_sr[4]), .Y(n336) );
  XOR2X1 U943 ( .A(w0[28]), .B(sa10_sr[4]), .Y(n156) );
  XOR2X1 U405 ( .A(w3[0]), .B(sa23_sr[0]), .Y(n507) );
  XOR2X1 U407 ( .A(n507), .B(n506), .Y(sa33_next[0]) );
  XOR2X1 U502 ( .A(w3[24]), .B(sa13_sr[0]), .Y(n436) );
  XOR2X1 U504 ( .A(n436), .B(n435), .Y(sa03_next[0]) );
  XOR2X1 U440 ( .A(w3[8]), .B(sa33_sr[0]), .Y(n481) );
  XOR2X1 U442 ( .A(n481), .B(n480), .Y(sa23_next[0]) );
  XOR2X1 U467 ( .A(w3[16]), .B(sa03_sr[0]), .Y(n462) );
  XOR2X1 U469 ( .A(n462), .B(n461), .Y(sa13_next[0]) );
  XOR2X1 U512 ( .A(w3[26]), .B(sa13_sr[2]), .Y(n431) );
  XOR2X1 U514 ( .A(n431), .B(n430), .Y(sa03_next[2]) );
  XOR2XL U447 ( .A(w3[10]), .B(sa33_sr[2]), .Y(n476) );
  XOR2X1 U449 ( .A(n476), .B(n475), .Y(sa23_next[2]) );
  XOR2X1 U414 ( .A(sa23_sr[2]), .B(sa33_sr[1]), .Y(n500) );
  XOR2X1 U416 ( .A(n500), .B(n499), .Y(sa33_next[2]) );
  XOR2X1 U518 ( .A(n571), .B(n576), .Y(n428) );
  XOR2X1 U520 ( .A(n428), .B(n427), .Y(sa03_next[3]) );
  XOR2X1 U424 ( .A(n579), .B(n574), .Y(n492) );
  XOR2X1 U426 ( .A(n492), .B(n491), .Y(sa33_next[4]) );
  XOR2X1 U452 ( .A(n567), .B(n474), .Y(n472) );
  XOR2X1 U453 ( .A(n473), .B(n472), .Y(sa23_next[3]) );
  XOR2X1 U486 ( .A(n562), .B(n565), .Y(n447) );
  XOR2X1 U488 ( .A(n447), .B(n446), .Y(sa13_next[4]) );
  XOR2X1 U482 ( .A(n453), .B(n452), .Y(n450) );
  XOR2X1 U483 ( .A(n451), .B(n450), .Y(sa13_next[3]) );
  XOR2X1 U464 ( .A(w3[15]), .B(sa33_sr[7]), .Y(n464) );
  XOR2X1 U466 ( .A(n464), .B(n463), .Y(sa23_next[7]) );
  XOR2X1 U540 ( .A(w3[31]), .B(sa13_sr[7]), .Y(n419) );
  XOR2X1 U542 ( .A(n419), .B(n418), .Y(sa03_next[7]) );
  XOR2X1 U499 ( .A(sa13_sr[6]), .B(sa23_sr[6]), .Y(n438) );
  XOR2X1 U501 ( .A(n438), .B(n437), .Y(sa13_next[7]) );
  XOR2X1 U437 ( .A(sa23_sr[7]), .B(sa33_sr[6]), .Y(n483) );
  XOR2X1 U439 ( .A(n483), .B(n482), .Y(sa33_next[7]) );
  XOR2X1 U530 ( .A(w3[29]), .B(sa13_sr[5]), .Y(n423) );
  XOR2X1 U532 ( .A(n423), .B(n422), .Y(sa03_next[5]) );
  XOR2X1 U458 ( .A(w3[13]), .B(sa33_sr[5]), .Y(n468) );
  XOR2X1 U460 ( .A(n468), .B(n467), .Y(sa23_next[5]) );
  XOR2X1 U429 ( .A(sa23_sr[5]), .B(sa33_sr[4]), .Y(n489) );
  XOR2X1 U431 ( .A(n489), .B(n488), .Y(sa33_next[5]) );
  XOR2X1 U491 ( .A(sa13_sr[4]), .B(sa23_sr[4]), .Y(n444) );
  XOR2X1 U493 ( .A(n444), .B(n443), .Y(sa13_next[5]) );
  XOR2X1 U508 ( .A(n568), .B(n434), .Y(n432) );
  XOR2X1 U509 ( .A(n433), .B(n432), .Y(sa03_next[1]) );
  XOR2X1 U444 ( .A(n570), .B(n577), .Y(n478) );
  XOR2X1 U446 ( .A(n478), .B(n477), .Y(sa23_next[1]) );
  XOR2X1 U472 ( .A(n562), .B(n568), .Y(n458) );
  XOR2X1 U474 ( .A(n458), .B(n457), .Y(sa13_next[1]) );
  XOR2X1 U535 ( .A(w3[30]), .B(sa13_sr[6]), .Y(n421) );
  XOR2X1 U537 ( .A(n421), .B(n420), .Y(sa03_next[6]) );
  XOR2X1 U461 ( .A(w3[14]), .B(sa33_sr[6]), .Y(n466) );
  XOR2X1 U463 ( .A(n466), .B(n465), .Y(sa23_next[6]) );
  XOR2X1 U433 ( .A(sa23_sr[6]), .B(sa33_sr[5]), .Y(n486) );
  XOR2X1 U435 ( .A(n486), .B(n485), .Y(sa33_next[6]) );
  XOR2X1 U495 ( .A(sa13_sr[5]), .B(sa23_sr[5]), .Y(n441) );
  XOR2X1 U497 ( .A(n441), .B(n440), .Y(sa13_next[6]) );
  XOR2X1 U922 ( .A(w0[24]), .B(sa10_sr[0]), .Y(n166) );
  XOR2X1 U924 ( .A(n166), .B(n165), .Y(sa00_next[0]) );
  XOR2X1 U825 ( .A(w0[0]), .B(sa20_sr[0]), .Y(n237) );
  XOR2X1 U827 ( .A(n237), .B(n236), .Y(sa30_next[0]) );
  XOR2X1 U685 ( .A(w1[0]), .B(sa21_sr[0]), .Y(n327) );
  XOR2X1 U687 ( .A(n327), .B(n326), .Y(sa31_next[0]) );
  XOR2X1 U545 ( .A(w2[0]), .B(sa22_sr[0]), .Y(n417) );
  XOR2X1 U547 ( .A(n417), .B(n416), .Y(sa32_next[0]) );
  XOR2X1 U607 ( .A(w2[16]), .B(sa02_sr[0]), .Y(n372) );
  XOR2X1 U609 ( .A(n372), .B(n371), .Y(sa12_next[0]) );
  XOR2X1 U747 ( .A(w1[16]), .B(sa01_sr[0]), .Y(n282) );
  XOR2X1 U749 ( .A(n282), .B(n281), .Y(sa11_next[0]) );
  XOR2X1 U887 ( .A(w0[16]), .B(sa00_sr[0]), .Y(n192) );
  XOR2X1 U889 ( .A(n192), .B(n191), .Y(sa10_next[0]) );
  XOR2X1 U782 ( .A(w1[24]), .B(sa11_sr[0]), .Y(n256) );
  XOR2X1 U784 ( .A(n256), .B(n255), .Y(sa01_next[0]) );
  XOR2X1 U720 ( .A(w1[8]), .B(sa31_sr[0]), .Y(n301) );
  XOR2X1 U722 ( .A(n301), .B(n300), .Y(sa21_next[0]) );
  XOR2X1 U642 ( .A(w2[24]), .B(sa12_sr[0]), .Y(n346) );
  XOR2X1 U644 ( .A(n346), .B(n345), .Y(sa02_next[0]) );
  XOR2X1 U580 ( .A(w2[8]), .B(sa32_sr[0]), .Y(n391) );
  XOR2X1 U582 ( .A(n391), .B(n390), .Y(sa22_next[0]) );
  XOR2X1 U860 ( .A(w0[8]), .B(sa30_sr[0]), .Y(n211) );
  XOR2X1 U862 ( .A(n211), .B(n210), .Y(sa20_next[0]) );
  XOR2X1 U810 ( .A(w1[29]), .B(sa11_sr[5]), .Y(n243) );
  XOR2X1 U812 ( .A(n243), .B(n242), .Y(sa01_next[5]) );
  XOR2X1 U738 ( .A(w1[13]), .B(sa31_sr[5]), .Y(n288) );
  XOR2X1 U740 ( .A(n288), .B(n287), .Y(sa21_next[5]) );
  XOR2X1 U771 ( .A(sa11_sr[4]), .B(sa21_sr[4]), .Y(n264) );
  XOR2X1 U773 ( .A(n264), .B(n263), .Y(sa11_next[5]) );
  XOR2X1 U670 ( .A(w2[29]), .B(sa12_sr[5]), .Y(n333) );
  XOR2X1 U672 ( .A(n333), .B(n332), .Y(sa02_next[5]) );
  XOR2X1 U598 ( .A(w2[13]), .B(sa32_sr[5]), .Y(n378) );
  XOR2X1 U600 ( .A(n378), .B(n377), .Y(sa22_next[5]) );
  XOR2X1 U631 ( .A(sa12_sr[4]), .B(sa22_sr[4]), .Y(n354) );
  XOR2X1 U633 ( .A(n354), .B(n353), .Y(sa12_next[5]) );
  XOR2X1 U878 ( .A(w0[13]), .B(sa30_sr[5]), .Y(n198) );
  XOR2X1 U880 ( .A(n198), .B(n197), .Y(sa20_next[5]) );
  XOR2X1 U950 ( .A(w0[29]), .B(sa10_sr[5]), .Y(n153) );
  XOR2X1 U952 ( .A(n153), .B(n152), .Y(sa00_next[5]) );
  XOR2X1 U911 ( .A(sa10_sr[4]), .B(sa20_sr[4]), .Y(n174) );
  XOR2X1 U913 ( .A(n174), .B(n173), .Y(sa10_next[5]) );
  XOR2X1 U792 ( .A(w1[26]), .B(sa11_sr[2]), .Y(n251) );
  XOR2X1 U794 ( .A(n251), .B(n250), .Y(sa01_next[2]) );
  XOR2XL U727 ( .A(w1[10]), .B(sa31_sr[2]), .Y(n296) );
  XOR2X1 U729 ( .A(n296), .B(n295), .Y(sa21_next[2]) );
  XOR2X1 U694 ( .A(sa21_sr[2]), .B(sa31_sr[1]), .Y(n320) );
  XOR2X1 U696 ( .A(n320), .B(n319), .Y(sa31_next[2]) );
  XOR2X1 U652 ( .A(w2[26]), .B(sa12_sr[2]), .Y(n341) );
  XOR2X1 U654 ( .A(n341), .B(n340), .Y(sa02_next[2]) );
  XOR2XL U587 ( .A(w2[10]), .B(sa32_sr[2]), .Y(n386) );
  XOR2X1 U589 ( .A(n386), .B(n385), .Y(sa22_next[2]) );
  XOR2X1 U554 ( .A(sa22_sr[2]), .B(sa32_sr[1]), .Y(n410) );
  XOR2X1 U556 ( .A(n410), .B(n409), .Y(sa32_next[2]) );
  XOR2XL U867 ( .A(w0[10]), .B(sa30_sr[2]), .Y(n206) );
  XOR2X1 U869 ( .A(n206), .B(n205), .Y(sa20_next[2]) );
  XOR2X1 U932 ( .A(w0[26]), .B(sa10_sr[2]), .Y(n161) );
  XOR2X1 U934 ( .A(n161), .B(n160), .Y(sa00_next[2]) );
  XOR2X1 U834 ( .A(sa20_sr[2]), .B(sa30_sr[1]), .Y(n230) );
  XOR2X1 U836 ( .A(n230), .B(n229), .Y(sa30_next[2]) );
  XOR2X1 U884 ( .A(w0[15]), .B(sa30_sr[7]), .Y(n194) );
  XOR2X1 U886 ( .A(n194), .B(n193), .Y(sa20_next[7]) );
  XOR2X1 U820 ( .A(w1[31]), .B(sa11_sr[7]), .Y(n239) );
  XOR2X1 U822 ( .A(n239), .B(n238), .Y(sa01_next[7]) );
  XOR2X1 U744 ( .A(w1[15]), .B(sa31_sr[7]), .Y(n284) );
  XOR2X1 U746 ( .A(n284), .B(n283), .Y(sa21_next[7]) );
  XOR2X1 U779 ( .A(sa11_sr[6]), .B(sa21_sr[6]), .Y(n258) );
  XOR2X1 U781 ( .A(n258), .B(n257), .Y(sa11_next[7]) );
  XOR2X1 U717 ( .A(sa21_sr[7]), .B(sa31_sr[6]), .Y(n303) );
  XOR2X1 U719 ( .A(n303), .B(n302), .Y(sa31_next[7]) );
  XOR2X1 U680 ( .A(w2[31]), .B(sa12_sr[7]), .Y(n329) );
  XOR2X1 U682 ( .A(n329), .B(n328), .Y(sa02_next[7]) );
  XOR2X1 U639 ( .A(sa12_sr[6]), .B(sa22_sr[6]), .Y(n348) );
  XOR2X1 U641 ( .A(n348), .B(n347), .Y(sa12_next[7]) );
  XOR2X1 U604 ( .A(w2[15]), .B(sa32_sr[7]), .Y(n374) );
  XOR2X1 U606 ( .A(n374), .B(n373), .Y(sa22_next[7]) );
  XOR2X1 U960 ( .A(w0[31]), .B(sa10_sr[7]), .Y(n149) );
  XOR2X1 U962 ( .A(n149), .B(n148), .Y(sa00_next[7]) );
  XOR2X1 U919 ( .A(sa10_sr[6]), .B(sa20_sr[6]), .Y(n168) );
  XOR2X1 U921 ( .A(n168), .B(n167), .Y(sa10_next[7]) );
  XOR2X1 U857 ( .A(sa20_sr[7]), .B(sa30_sr[6]), .Y(n213) );
  XOR2X1 U859 ( .A(n213), .B(n212), .Y(sa30_next[7]) );
  XOR2X1 U577 ( .A(sa22_sr[7]), .B(sa32_sr[6]), .Y(n393) );
  XOR2X1 U579 ( .A(n393), .B(n392), .Y(sa32_next[7]) );
  XOR2X1 U762 ( .A(n273), .B(n272), .Y(n270) );
  XOR2X1 U763 ( .A(n271), .B(n270), .Y(sa11_next[3]) );
  XOR2X1 U704 ( .A(n543), .B(n538), .Y(n312) );
  XOR2X1 U706 ( .A(n312), .B(n311), .Y(sa31_next[4]) );
  XOR2X1 U766 ( .A(n526), .B(n529), .Y(n267) );
  XOR2X1 U768 ( .A(n267), .B(n266), .Y(sa11_next[4]) );
  XOR2X1 U798 ( .A(n535), .B(n540), .Y(n248) );
  XOR2X1 U800 ( .A(n248), .B(n247), .Y(sa01_next[3]) );
  XOR2X1 U732 ( .A(n531), .B(n294), .Y(n292) );
  XOR2X1 U733 ( .A(n293), .B(n292), .Y(sa21_next[3]) );
  XOR2X1 U658 ( .A(n553), .B(n558), .Y(n338) );
  XOR2X1 U660 ( .A(n338), .B(n337), .Y(sa02_next[3]) );
  XOR2X1 U592 ( .A(n549), .B(n384), .Y(n382) );
  XOR2X1 U593 ( .A(n383), .B(n382), .Y(sa22_next[3]) );
  XOR2X1 U622 ( .A(n363), .B(n362), .Y(n360) );
  XOR2X1 U623 ( .A(n361), .B(n360), .Y(sa12_next[3]) );
  XOR2X1 U564 ( .A(n561), .B(n556), .Y(n402) );
  XOR2X1 U566 ( .A(n402), .B(n401), .Y(sa32_next[4]) );
  XOR2X1 U626 ( .A(n544), .B(n547), .Y(n357) );
  XOR2X1 U628 ( .A(n357), .B(n356), .Y(sa12_next[4]) );
  XOR2X1 U938 ( .A(n517), .B(n522), .Y(n158) );
  XOR2X1 U940 ( .A(n158), .B(n157), .Y(sa00_next[3]) );
  XOR2X1 U902 ( .A(n183), .B(n182), .Y(n180) );
  XOR2X1 U903 ( .A(n181), .B(n180), .Y(sa10_next[3]) );
  XOR2X1 U906 ( .A(n508), .B(n511), .Y(n177) );
  XOR2X1 U908 ( .A(n177), .B(n176), .Y(sa10_next[4]) );
  XOR2X1 U844 ( .A(n525), .B(n520), .Y(n222) );
  XOR2X1 U846 ( .A(n222), .B(n221), .Y(sa30_next[4]) );
  XOR2X1 U872 ( .A(n513), .B(n204), .Y(n202) );
  XOR2X1 U873 ( .A(n203), .B(n202), .Y(sa20_next[3]) );
  XOR2X1 U752 ( .A(n526), .B(n532), .Y(n278) );
  XOR2X1 U754 ( .A(n278), .B(n277), .Y(sa11_next[1]) );
  XOR2X1 U788 ( .A(n532), .B(n254), .Y(n252) );
  XOR2X1 U789 ( .A(n253), .B(n252), .Y(sa01_next[1]) );
  XOR2X1 U724 ( .A(n534), .B(n541), .Y(n298) );
  XOR2X1 U726 ( .A(n298), .B(n297), .Y(sa21_next[1]) );
  XOR2X1 U648 ( .A(n550), .B(n344), .Y(n342) );
  XOR2X1 U649 ( .A(n343), .B(n342), .Y(sa02_next[1]) );
  XOR2X1 U584 ( .A(n552), .B(n559), .Y(n388) );
  XOR2X1 U586 ( .A(n388), .B(n387), .Y(sa22_next[1]) );
  XOR2X1 U612 ( .A(n544), .B(n550), .Y(n368) );
  XOR2X1 U614 ( .A(n368), .B(n367), .Y(sa12_next[1]) );
  XOR2X1 U928 ( .A(n514), .B(n164), .Y(n162) );
  XOR2X1 U929 ( .A(n163), .B(n162), .Y(sa00_next[1]) );
  XOR2X1 U892 ( .A(n508), .B(n514), .Y(n188) );
  XOR2X1 U894 ( .A(n188), .B(n187), .Y(sa10_next[1]) );
  XOR2X1 U864 ( .A(n516), .B(n523), .Y(n208) );
  XOR2X1 U866 ( .A(n208), .B(n207), .Y(sa20_next[1]) );
  XOR2X1 U815 ( .A(w1[30]), .B(sa11_sr[6]), .Y(n241) );
  XOR2X1 U817 ( .A(n241), .B(n240), .Y(sa01_next[6]) );
  XOR2X1 U741 ( .A(w1[14]), .B(sa31_sr[6]), .Y(n286) );
  XOR2X1 U743 ( .A(n286), .B(n285), .Y(sa21_next[6]) );
  XOR2X1 U713 ( .A(sa21_sr[6]), .B(sa31_sr[5]), .Y(n306) );
  XOR2X1 U715 ( .A(n306), .B(n305), .Y(sa31_next[6]) );
  XOR2X1 U675 ( .A(w2[30]), .B(sa12_sr[6]), .Y(n331) );
  XOR2X1 U677 ( .A(n331), .B(n330), .Y(sa02_next[6]) );
  XOR2X1 U601 ( .A(w2[14]), .B(sa32_sr[6]), .Y(n376) );
  XOR2X1 U603 ( .A(n376), .B(n375), .Y(sa22_next[6]) );
  XOR2X1 U573 ( .A(sa22_sr[6]), .B(sa32_sr[5]), .Y(n396) );
  XOR2X1 U575 ( .A(n396), .B(n395), .Y(sa32_next[6]) );
  XOR2X1 U881 ( .A(w0[14]), .B(sa30_sr[6]), .Y(n196) );
  XOR2X1 U883 ( .A(n196), .B(n195), .Y(sa20_next[6]) );
  XOR2X1 U955 ( .A(w0[30]), .B(sa10_sr[6]), .Y(n151) );
  XOR2X1 U957 ( .A(n151), .B(n150), .Y(sa00_next[6]) );
  XOR2X1 U853 ( .A(sa20_sr[6]), .B(sa30_sr[5]), .Y(n216) );
  XOR2X1 U855 ( .A(n216), .B(n215), .Y(sa30_next[6]) );
  XOR2X1 U523 ( .A(w3[28]), .B(sa13_sr[4]), .Y(n426) );
  XOR2X1 U703 ( .A(sa21_sr[4]), .B(sa31_sr[3]), .Y(n313) );
  XOR2X1 U702 ( .A(w1[4]), .B(sa01_sr[3]), .Y(n314) );
  XOR2X1 U705 ( .A(n314), .B(n313), .Y(n311) );
  XOR2X1 U423 ( .A(sa23_sr[4]), .B(sa33_sr[3]), .Y(n493) );
  XOR2X1 U422 ( .A(w3[4]), .B(sa03_sr[3]), .Y(n494) );
  XOR2X1 U425 ( .A(n494), .B(n493), .Y(n491) );
  XOR2X1 U563 ( .A(sa22_sr[4]), .B(sa32_sr[3]), .Y(n403) );
  XOR2X1 U562 ( .A(w2[4]), .B(sa02_sr[3]), .Y(n404) );
  XOR2X1 U565 ( .A(n404), .B(n403), .Y(n401) );
  XOR2X1 U843 ( .A(sa20_sr[4]), .B(sa30_sr[3]), .Y(n223) );
  XOR2X1 U842 ( .A(w0[4]), .B(sa00_sr[3]), .Y(n224) );
  XOR2X1 U845 ( .A(n224), .B(n223), .Y(n221) );
  XOR2X1 U450 ( .A(w3[11]), .B(sa33_sr[3]), .Y(n474) );
  DFFHQX1 done_reg ( .D(N21), .CK(clk), .Q(done) );
  DFFHQX1 \text_out_reg[127]  ( .D(N376), .CK(clk), .Q(text_out[127]) );
  DFFHQX1 \text_out_reg[126]  ( .D(N377), .CK(clk), .Q(text_out[126]) );
  DFFHQX1 \text_out_reg[125]  ( .D(N378), .CK(clk), .Q(text_out[125]) );
  DFFHQX1 \text_out_reg[124]  ( .D(N379), .CK(clk), .Q(text_out[124]) );
  DFFHQX1 \text_out_reg[123]  ( .D(N380), .CK(clk), .Q(text_out[123]) );
  DFFHQX1 \text_out_reg[122]  ( .D(N381), .CK(clk), .Q(text_out[122]) );
  DFFHQX1 \text_out_reg[121]  ( .D(N382), .CK(clk), .Q(text_out[121]) );
  DFFHQX1 \text_out_reg[120]  ( .D(N383), .CK(clk), .Q(text_out[120]) );
  DFFHQX1 \text_out_reg[95]  ( .D(N384), .CK(clk), .Q(text_out[95]) );
  DFFHQX1 \text_out_reg[94]  ( .D(N385), .CK(clk), .Q(text_out[94]) );
  DFFHQX1 \text_out_reg[93]  ( .D(N386), .CK(clk), .Q(text_out[93]) );
  DFFHQX1 \text_out_reg[92]  ( .D(N387), .CK(clk), .Q(text_out[92]) );
  DFFHQX1 \text_out_reg[91]  ( .D(N388), .CK(clk), .Q(text_out[91]) );
  DFFHQX1 \text_out_reg[90]  ( .D(N389), .CK(clk), .Q(text_out[90]) );
  DFFHQX1 \text_out_reg[89]  ( .D(N390), .CK(clk), .Q(text_out[89]) );
  DFFHQX1 \text_out_reg[88]  ( .D(N391), .CK(clk), .Q(text_out[88]) );
  DFFHQX1 \text_out_reg[63]  ( .D(N392), .CK(clk), .Q(text_out[63]) );
  DFFHQX1 \text_out_reg[62]  ( .D(N393), .CK(clk), .Q(text_out[62]) );
  DFFHQX1 \text_out_reg[61]  ( .D(N394), .CK(clk), .Q(text_out[61]) );
  DFFHQX1 \text_out_reg[60]  ( .D(N395), .CK(clk), .Q(text_out[60]) );
  DFFHQX1 \text_out_reg[59]  ( .D(N396), .CK(clk), .Q(text_out[59]) );
  DFFHQX1 \text_out_reg[58]  ( .D(N397), .CK(clk), .Q(text_out[58]) );
  DFFHQX1 \text_out_reg[57]  ( .D(N398), .CK(clk), .Q(text_out[57]) );
  DFFHQX1 \text_out_reg[56]  ( .D(N399), .CK(clk), .Q(text_out[56]) );
  DFFHQX1 \text_out_reg[31]  ( .D(N400), .CK(clk), .Q(text_out[31]) );
  DFFHQX1 \text_out_reg[30]  ( .D(N401), .CK(clk), .Q(text_out[30]) );
  DFFHQX1 \text_out_reg[29]  ( .D(N402), .CK(clk), .Q(text_out[29]) );
  DFFHQX1 \text_out_reg[28]  ( .D(N403), .CK(clk), .Q(text_out[28]) );
  DFFHQX1 \text_out_reg[27]  ( .D(N404), .CK(clk), .Q(text_out[27]) );
  DFFHQX1 \text_out_reg[26]  ( .D(N405), .CK(clk), .Q(text_out[26]) );
  DFFHQX1 \text_out_reg[25]  ( .D(N406), .CK(clk), .Q(text_out[25]) );
  DFFHQX1 \text_out_reg[24]  ( .D(N407), .CK(clk), .Q(text_out[24]) );
  DFFHQX1 \text_out_reg[119]  ( .D(N408), .CK(clk), .Q(text_out[119]) );
  DFFHQX1 \text_out_reg[118]  ( .D(N409), .CK(clk), .Q(text_out[118]) );
  DFFHQX1 \text_out_reg[117]  ( .D(N410), .CK(clk), .Q(text_out[117]) );
  DFFHQX1 \text_out_reg[116]  ( .D(N411), .CK(clk), .Q(text_out[116]) );
  DFFHQX1 \text_out_reg[115]  ( .D(N412), .CK(clk), .Q(text_out[115]) );
  DFFHQX1 \text_out_reg[114]  ( .D(N413), .CK(clk), .Q(text_out[114]) );
  DFFHQX1 \text_out_reg[113]  ( .D(N414), .CK(clk), .Q(text_out[113]) );
  DFFHQX1 \text_out_reg[112]  ( .D(N415), .CK(clk), .Q(text_out[112]) );
  DFFHQX1 \text_out_reg[87]  ( .D(N416), .CK(clk), .Q(text_out[87]) );
  DFFHQX1 \text_out_reg[86]  ( .D(N417), .CK(clk), .Q(text_out[86]) );
  DFFHQX1 \text_out_reg[85]  ( .D(N418), .CK(clk), .Q(text_out[85]) );
  DFFHQX1 \text_out_reg[84]  ( .D(N419), .CK(clk), .Q(text_out[84]) );
  DFFHQX1 \text_out_reg[83]  ( .D(N420), .CK(clk), .Q(text_out[83]) );
  DFFHQX1 \text_out_reg[82]  ( .D(N421), .CK(clk), .Q(text_out[82]) );
  DFFHQX1 \text_out_reg[81]  ( .D(N422), .CK(clk), .Q(text_out[81]) );
  DFFHQX1 \text_out_reg[80]  ( .D(N423), .CK(clk), .Q(text_out[80]) );
  DFFHQX1 \text_out_reg[55]  ( .D(N424), .CK(clk), .Q(text_out[55]) );
  DFFHQX1 \text_out_reg[54]  ( .D(N425), .CK(clk), .Q(text_out[54]) );
  DFFHQX1 \text_out_reg[53]  ( .D(N426), .CK(clk), .Q(text_out[53]) );
  DFFHQX1 \text_out_reg[52]  ( .D(N427), .CK(clk), .Q(text_out[52]) );
  DFFHQX1 \text_out_reg[51]  ( .D(N428), .CK(clk), .Q(text_out[51]) );
  DFFHQX1 \text_out_reg[50]  ( .D(N429), .CK(clk), .Q(text_out[50]) );
  DFFHQX1 \text_out_reg[49]  ( .D(N430), .CK(clk), .Q(text_out[49]) );
  DFFHQX1 \text_out_reg[48]  ( .D(N431), .CK(clk), .Q(text_out[48]) );
  DFFHQX1 \text_out_reg[23]  ( .D(N432), .CK(clk), .Q(text_out[23]) );
  DFFHQX1 \text_out_reg[22]  ( .D(N433), .CK(clk), .Q(text_out[22]) );
  DFFHQX1 \text_out_reg[21]  ( .D(N434), .CK(clk), .Q(text_out[21]) );
  DFFHQX1 \text_out_reg[20]  ( .D(N435), .CK(clk), .Q(text_out[20]) );
  DFFHQX1 \text_out_reg[19]  ( .D(N436), .CK(clk), .Q(text_out[19]) );
  DFFHQX1 \text_out_reg[18]  ( .D(N437), .CK(clk), .Q(text_out[18]) );
  DFFHQX1 \text_out_reg[17]  ( .D(N438), .CK(clk), .Q(text_out[17]) );
  DFFHQX1 \text_out_reg[16]  ( .D(N439), .CK(clk), .Q(text_out[16]) );
  DFFHQX1 \text_out_reg[111]  ( .D(N440), .CK(clk), .Q(text_out[111]) );
  DFFHQX1 \text_out_reg[110]  ( .D(N441), .CK(clk), .Q(text_out[110]) );
  DFFHQX1 \text_out_reg[109]  ( .D(N442), .CK(clk), .Q(text_out[109]) );
  DFFHQX1 \text_out_reg[108]  ( .D(N443), .CK(clk), .Q(text_out[108]) );
  DFFHQX1 \text_out_reg[107]  ( .D(N444), .CK(clk), .Q(text_out[107]) );
  DFFHQX1 \text_out_reg[106]  ( .D(N445), .CK(clk), .Q(text_out[106]) );
  DFFHQX1 \text_out_reg[105]  ( .D(N446), .CK(clk), .Q(text_out[105]) );
  DFFHQX1 \text_out_reg[104]  ( .D(N447), .CK(clk), .Q(text_out[104]) );
  DFFHQX1 \text_out_reg[79]  ( .D(N448), .CK(clk), .Q(text_out[79]) );
  DFFHQX1 \text_out_reg[78]  ( .D(N449), .CK(clk), .Q(text_out[78]) );
  DFFHQX1 \text_out_reg[77]  ( .D(N450), .CK(clk), .Q(text_out[77]) );
  DFFHQX1 \text_out_reg[76]  ( .D(N451), .CK(clk), .Q(text_out[76]) );
  DFFHQX1 \text_out_reg[75]  ( .D(N452), .CK(clk), .Q(text_out[75]) );
  DFFHQX1 \text_out_reg[74]  ( .D(N453), .CK(clk), .Q(text_out[74]) );
  DFFHQX1 \text_out_reg[73]  ( .D(N454), .CK(clk), .Q(text_out[73]) );
  DFFHQX1 \text_out_reg[72]  ( .D(N455), .CK(clk), .Q(text_out[72]) );
  DFFHQX1 \text_out_reg[47]  ( .D(N456), .CK(clk), .Q(text_out[47]) );
  DFFHQX1 \text_out_reg[46]  ( .D(N457), .CK(clk), .Q(text_out[46]) );
  DFFHQX1 \text_out_reg[45]  ( .D(N458), .CK(clk), .Q(text_out[45]) );
  DFFHQX1 \text_out_reg[44]  ( .D(N459), .CK(clk), .Q(text_out[44]) );
  DFFHQX1 \text_out_reg[43]  ( .D(N460), .CK(clk), .Q(text_out[43]) );
  DFFHQX1 \text_out_reg[42]  ( .D(N461), .CK(clk), .Q(text_out[42]) );
  DFFHQX1 \text_out_reg[41]  ( .D(N462), .CK(clk), .Q(text_out[41]) );
  DFFHQX1 \text_out_reg[40]  ( .D(N463), .CK(clk), .Q(text_out[40]) );
  DFFHQX1 \text_out_reg[15]  ( .D(N464), .CK(clk), .Q(text_out[15]) );
  DFFHQX1 \text_out_reg[14]  ( .D(N465), .CK(clk), .Q(text_out[14]) );
  DFFHQX1 \text_out_reg[13]  ( .D(N466), .CK(clk), .Q(text_out[13]) );
  DFFHQX1 \text_out_reg[12]  ( .D(N467), .CK(clk), .Q(text_out[12]) );
  DFFHQX1 \text_out_reg[11]  ( .D(N468), .CK(clk), .Q(text_out[11]) );
  DFFHQX1 \text_out_reg[10]  ( .D(N469), .CK(clk), .Q(text_out[10]) );
  DFFHQX1 \text_out_reg[9]  ( .D(N470), .CK(clk), .Q(text_out[9]) );
  DFFHQX1 \text_out_reg[8]  ( .D(N471), .CK(clk), .Q(text_out[8]) );
  DFFHQX1 \text_out_reg[103]  ( .D(N472), .CK(clk), .Q(text_out[103]) );
  DFFHQX1 \text_out_reg[102]  ( .D(N473), .CK(clk), .Q(text_out[102]) );
  DFFHQX1 \text_out_reg[101]  ( .D(N474), .CK(clk), .Q(text_out[101]) );
  DFFHQX1 \text_out_reg[100]  ( .D(N475), .CK(clk), .Q(text_out[100]) );
  DFFHQX1 \text_out_reg[99]  ( .D(N476), .CK(clk), .Q(text_out[99]) );
  DFFHQX1 \text_out_reg[98]  ( .D(N477), .CK(clk), .Q(text_out[98]) );
  DFFHQX1 \text_out_reg[97]  ( .D(N478), .CK(clk), .Q(text_out[97]) );
  DFFHQX1 \text_out_reg[96]  ( .D(N479), .CK(clk), .Q(text_out[96]) );
  DFFHQX1 \text_out_reg[71]  ( .D(N480), .CK(clk), .Q(text_out[71]) );
  DFFHQX1 \text_out_reg[70]  ( .D(N481), .CK(clk), .Q(text_out[70]) );
  DFFHQX1 \text_out_reg[69]  ( .D(N482), .CK(clk), .Q(text_out[69]) );
  DFFHQX1 \text_out_reg[68]  ( .D(N483), .CK(clk), .Q(text_out[68]) );
  DFFHQX1 \text_out_reg[67]  ( .D(N484), .CK(clk), .Q(text_out[67]) );
  DFFHQX1 \text_out_reg[66]  ( .D(N485), .CK(clk), .Q(text_out[66]) );
  DFFHQX1 \text_out_reg[65]  ( .D(N486), .CK(clk), .Q(text_out[65]) );
  DFFHQX1 \text_out_reg[64]  ( .D(N487), .CK(clk), .Q(text_out[64]) );
  DFFHQX1 \text_out_reg[39]  ( .D(N488), .CK(clk), .Q(text_out[39]) );
  DFFHQX1 \text_out_reg[38]  ( .D(N489), .CK(clk), .Q(text_out[38]) );
  DFFHQX1 \text_out_reg[37]  ( .D(N490), .CK(clk), .Q(text_out[37]) );
  DFFHQX1 \text_out_reg[36]  ( .D(N491), .CK(clk), .Q(text_out[36]) );
  DFFHQX1 \text_out_reg[35]  ( .D(N492), .CK(clk), .Q(text_out[35]) );
  DFFHQX1 \text_out_reg[34]  ( .D(N493), .CK(clk), .Q(text_out[34]) );
  DFFHQX1 \text_out_reg[33]  ( .D(N494), .CK(clk), .Q(text_out[33]) );
  DFFHQX1 \text_out_reg[32]  ( .D(N495), .CK(clk), .Q(text_out[32]) );
  DFFHQX1 \text_out_reg[7]  ( .D(N496), .CK(clk), .Q(text_out[7]) );
  DFFHQX1 \text_out_reg[6]  ( .D(N497), .CK(clk), .Q(text_out[6]) );
  DFFHQX1 \text_out_reg[5]  ( .D(N498), .CK(clk), .Q(text_out[5]) );
  DFFHQX1 \text_out_reg[4]  ( .D(N499), .CK(clk), .Q(text_out[4]) );
  DFFHQX1 \text_out_reg[3]  ( .D(N500), .CK(clk), .Q(text_out[3]) );
  DFFHQX1 \text_out_reg[2]  ( .D(N501), .CK(clk), .Q(text_out[2]) );
  DFFHQX1 \text_out_reg[1]  ( .D(N502), .CK(clk), .Q(text_out[1]) );
  DFFHQX1 \text_out_reg[0]  ( .D(N503), .CK(clk), .Q(text_out[0]) );
  DFFHQX1 \sa00_reg[0]  ( .D(N272), .CK(clk), .Q(sa00[0]) );
  DFFHQX1 \sa30_reg[0]  ( .D(N224), .CK(clk), .Q(sa30[0]) );
  DFFHQX1 \sa31_reg[0]  ( .D(N160), .CK(clk), .Q(sa31[0]) );
  DFFHQX1 \sa32_reg[0]  ( .D(N96), .CK(clk), .Q(sa32[0]) );
  DFFHQX1 \sa33_reg[0]  ( .D(N32), .CK(clk), .Q(sa33[0]) );
  DFFHQX1 \sa12_reg[0]  ( .D(N128), .CK(clk), .Q(sa12[0]) );
  DFFHQX1 \sa11_reg[0]  ( .D(N192), .CK(clk), .Q(sa11[0]) );
  DFFHQX1 \sa10_reg[0]  ( .D(N256), .CK(clk), .Q(sa10[0]) );
  DFFHQX1 \sa01_reg[0]  ( .D(N208), .CK(clk), .Q(sa01[0]) );
  DFFHQX1 \sa21_reg[0]  ( .D(N176), .CK(clk), .Q(sa21[0]) );
  DFFHQX1 \sa03_reg[0]  ( .D(N80), .CK(clk), .Q(sa03[0]) );
  DFFHQX1 \sa23_reg[0]  ( .D(N48), .CK(clk), .Q(sa23[0]) );
  DFFHQX1 \sa13_reg[0]  ( .D(N64), .CK(clk), .Q(sa13[0]) );
  DFFHQX1 \sa02_reg[0]  ( .D(N144), .CK(clk), .Q(sa02[0]) );
  DFFHQX1 \sa22_reg[0]  ( .D(N112), .CK(clk), .Q(sa22[0]) );
  DFFHQX1 \sa20_reg[0]  ( .D(N240), .CK(clk), .Q(sa20[0]) );
  XOR2X1 U698 ( .A(sa21_sr[3]), .B(sa31_sr[2]), .Y(n317) );
  XOR2X1 U418 ( .A(sa23_sr[3]), .B(sa33_sr[2]), .Y(n497) );
  XOR2X1 U558 ( .A(sa22_sr[3]), .B(sa32_sr[2]), .Y(n407) );
  XOR2X1 U838 ( .A(sa20_sr[3]), .B(sa30_sr[2]), .Y(n227) );
  XOR2X1 U801 ( .A(sa21_sr[3]), .B(sa31_sr[3]), .Y(n530) );
  XOR2X1 U521 ( .A(sa23_sr[3]), .B(sa33_sr[3]), .Y(n566) );
  XOR2X1 U661 ( .A(sa22_sr[3]), .B(sa32_sr[3]), .Y(n548) );
  XOR2X1 U941 ( .A(sa20_sr[3]), .B(sa30_sr[3]), .Y(n512) );
  XOR2X1 U925 ( .A(sa20_sr[0]), .B(sa30_sr[0]), .Y(n515) );
  XOR2X1 U645 ( .A(sa22_sr[0]), .B(sa32_sr[0]), .Y(n551) );
  XOR2X1 U785 ( .A(sa21_sr[0]), .B(sa31_sr[0]), .Y(n533) );
  XOR2X1 U505 ( .A(sa23_sr[0]), .B(sa33_sr[0]), .Y(n569) );
  DFFHQX1 \sa01_reg[2]  ( .D(N210), .CK(clk), .Q(sa01[2]) );
  DFFHQX1 \sa21_reg[2]  ( .D(N178), .CK(clk), .Q(sa21[2]) );
  DFFHQX1 \sa31_reg[2]  ( .D(N162), .CK(clk), .Q(sa31[2]) );
  DFFHQX1 \sa11_reg[2]  ( .D(N194), .CK(clk), .Q(sa11[2]) );
  DFFHQX1 \sa03_reg[2]  ( .D(N82), .CK(clk), .Q(sa03[2]) );
  DFFHQX1 \sa23_reg[2]  ( .D(N50), .CK(clk), .Q(sa23[2]) );
  DFFHQX1 \sa33_reg[2]  ( .D(N34), .CK(clk), .Q(sa33[2]) );
  DFFHQX1 \sa13_reg[2]  ( .D(N66), .CK(clk), .Q(sa13[2]) );
  DFFHQX1 \sa02_reg[2]  ( .D(N146), .CK(clk), .Q(sa02[2]) );
  DFFHQX1 \sa22_reg[2]  ( .D(N114), .CK(clk), .Q(sa22[2]) );
  DFFHQX1 \sa32_reg[2]  ( .D(N98), .CK(clk), .Q(sa32[2]) );
  DFFHQX1 \sa12_reg[2]  ( .D(N130), .CK(clk), .Q(sa12[2]) );
  DFFHQX1 \sa20_reg[2]  ( .D(N242), .CK(clk), .Q(sa20[2]) );
  DFFHQX1 \sa00_reg[2]  ( .D(N274), .CK(clk), .Q(sa00[2]) );
  DFFHQX1 \sa10_reg[2]  ( .D(N258), .CK(clk), .Q(sa10[2]) );
  DFFHQX1 \sa30_reg[2]  ( .D(N226), .CK(clk), .Q(sa30[2]) );
  XOR2X1 U699 ( .A(n543), .B(n539), .Y(n316) );
  XOR2X1 U419 ( .A(n579), .B(n575), .Y(n496) );
  XOR2X1 U559 ( .A(n561), .B(n557), .Y(n406) );
  XOR2X1 U839 ( .A(n525), .B(n521), .Y(n226) );
  XOR2X1 U761 ( .A(n526), .B(n530), .Y(n271) );
  XOR2X1 U481 ( .A(n562), .B(n566), .Y(n451) );
  XOR2X1 U621 ( .A(n544), .B(n548), .Y(n361) );
  XOR2X1 U901 ( .A(n508), .B(n512), .Y(n181) );
  XOR2X1 U804 ( .A(n535), .B(n539), .Y(n245) );
  XOR2X1 U731 ( .A(n534), .B(n539), .Y(n293) );
  XOR2X1 U524 ( .A(n571), .B(n575), .Y(n425) );
  XOR2X1 U451 ( .A(n570), .B(n575), .Y(n473) );
  XOR2X1 U664 ( .A(n553), .B(n557), .Y(n335) );
  XOR2X1 U591 ( .A(n552), .B(n557), .Y(n383) );
  XOR2X1 U944 ( .A(n517), .B(n521), .Y(n155) );
  XOR2X1 U871 ( .A(n516), .B(n521), .Y(n203) );
  XOR2X1 U787 ( .A(n535), .B(n542), .Y(n253) );
  XOR2X1 U507 ( .A(n571), .B(n578), .Y(n433) );
  XOR2X1 U647 ( .A(n553), .B(n560), .Y(n343) );
  XOR2X1 U927 ( .A(n517), .B(n524), .Y(n163) );
  XOR2X1 U923 ( .A(n517), .B(n515), .Y(n165) );
  XOR2X1 U608 ( .A(n544), .B(n551), .Y(n371) );
  XOR2X1 U748 ( .A(n526), .B(n533), .Y(n281) );
  XOR2X1 U888 ( .A(n508), .B(n515), .Y(n191) );
  XOR2X1 U783 ( .A(n535), .B(n533), .Y(n255) );
  XOR2X1 U503 ( .A(n571), .B(n569), .Y(n435) );
  XOR2X1 U468 ( .A(n562), .B(n569), .Y(n461) );
  XOR2X1 U643 ( .A(n553), .B(n551), .Y(n345) );
  XOR2X1 U826 ( .A(n525), .B(n524), .Y(n236) );
  XOR2X1 U686 ( .A(n543), .B(n542), .Y(n326) );
  XOR2X1 U546 ( .A(n561), .B(n560), .Y(n416) );
  XOR2X1 U406 ( .A(n579), .B(n578), .Y(n506) );
  XOR2X1 U721 ( .A(n534), .B(n542), .Y(n300) );
  XOR2X1 U441 ( .A(n570), .B(n578), .Y(n480) );
  XOR2X1 U581 ( .A(n552), .B(n560), .Y(n390) );
  XOR2X1 U861 ( .A(n516), .B(n524), .Y(n210) );
  XOR2X1 U760 ( .A(sa11_sr[2]), .B(sa21_sr[2]), .Y(n272) );
  XOR2X1 U480 ( .A(sa13_sr[2]), .B(sa23_sr[2]), .Y(n452) );
  XOR2X1 U620 ( .A(sa12_sr[2]), .B(sa22_sr[2]), .Y(n362) );
  XOR2X1 U900 ( .A(sa10_sr[2]), .B(sa20_sr[2]), .Y(n182) );
  XOR2X1 U819 ( .A(sa01_sr[5]), .B(sa11_sr[5]), .Y(n537) );
  XOR2X1 U539 ( .A(sa03_sr[5]), .B(sa13_sr[5]), .Y(n573) );
  XOR2X1 U679 ( .A(sa02_sr[5]), .B(sa12_sr[5]), .Y(n555) );
  XOR2X1 U959 ( .A(sa00_sr[5]), .B(sa10_sr[5]), .Y(n519) );
  XOR2X1 U847 ( .A(sa00_sr[7]), .B(sa30_sr[7]), .Y(n525) );
  XOR2X1 U707 ( .A(sa01_sr[7]), .B(sa31_sr[7]), .Y(n543) );
  XOR2X1 U567 ( .A(sa02_sr[7]), .B(sa32_sr[7]), .Y(n561) );
  XOR2X1 U427 ( .A(sa03_sr[7]), .B(sa33_sr[7]), .Y(n579) );
  XOR2X1 U629 ( .A(sa12_sr[7]), .B(sa22_sr[7]), .Y(n544) );
  XOR2X1 U769 ( .A(sa11_sr[7]), .B(sa21_sr[7]), .Y(n526) );
  XOR2X1 U909 ( .A(sa10_sr[7]), .B(sa20_sr[7]), .Y(n508) );
  XOR2X1 U489 ( .A(sa13_sr[7]), .B(sa23_sr[7]), .Y(n562) );
  XOR2X1 U823 ( .A(sa01_sr[6]), .B(sa11_sr[6]), .Y(n536) );
  XOR2X1 U543 ( .A(sa03_sr[6]), .B(sa13_sr[6]), .Y(n572) );
  XOR2X1 U683 ( .A(sa02_sr[6]), .B(sa12_sr[6]), .Y(n554) );
  XOR2X1 U963 ( .A(sa00_sr[6]), .B(sa10_sr[6]), .Y(n518) );
  XOR2X1 U795 ( .A(sa21_sr[2]), .B(sa31_sr[2]), .Y(n531) );
  XOR2X1 U515 ( .A(sa23_sr[2]), .B(sa33_sr[2]), .Y(n567) );
  XOR2X1 U655 ( .A(sa22_sr[2]), .B(sa32_sr[2]), .Y(n549) );
  XOR2X1 U935 ( .A(sa20_sr[2]), .B(sa30_sr[2]), .Y(n513) );
  XOR2X1 U802 ( .A(sa01_sr[2]), .B(sa11_sr[2]), .Y(n540) );
  XOR2X1 U522 ( .A(sa03_sr[2]), .B(sa13_sr[2]), .Y(n576) );
  XOR2X1 U662 ( .A(sa02_sr[2]), .B(sa12_sr[2]), .Y(n558) );
  XOR2X1 U942 ( .A(sa00_sr[2]), .B(sa10_sr[2]), .Y(n522) );
  XOR2X1 U796 ( .A(sa01_sr[1]), .B(sa11_sr[1]), .Y(n541) );
  XOR2X1 U516 ( .A(sa03_sr[1]), .B(sa13_sr[1]), .Y(n577) );
  XOR2X1 U656 ( .A(sa02_sr[1]), .B(sa12_sr[1]), .Y(n559) );
  XOR2X1 U936 ( .A(sa00_sr[1]), .B(sa10_sr[1]), .Y(n523) );
  XOR2X1 U813 ( .A(sa21_sr[5]), .B(sa31_sr[5]), .Y(n528) );
  XOR2X1 U533 ( .A(sa23_sr[5]), .B(sa33_sr[5]), .Y(n564) );
  XOR2X1 U673 ( .A(sa22_sr[5]), .B(sa32_sr[5]), .Y(n546) );
  XOR2X1 U953 ( .A(sa20_sr[5]), .B(sa30_sr[5]), .Y(n510) );
  XOR2X1 U790 ( .A(sa21_sr[1]), .B(sa31_sr[1]), .Y(n532) );
  XOR2X1 U510 ( .A(sa23_sr[1]), .B(sa33_sr[1]), .Y(n568) );
  XOR2X1 U650 ( .A(sa22_sr[1]), .B(sa32_sr[1]), .Y(n550) );
  XOR2X1 U930 ( .A(sa20_sr[1]), .B(sa30_sr[1]), .Y(n514) );
  XOR2X1 U958 ( .A(sa20_sr[6]), .B(sa30_sr[6]), .Y(n509) );
  XOR2X1 U538 ( .A(sa23_sr[6]), .B(sa33_sr[6]), .Y(n563) );
  XOR2X1 U818 ( .A(sa21_sr[6]), .B(sa31_sr[6]), .Y(n527) );
  XOR2X1 U678 ( .A(sa22_sr[6]), .B(sa32_sr[6]), .Y(n545) );
  XOR2X1 U807 ( .A(sa21_sr[4]), .B(sa31_sr[4]), .Y(n529) );
  XOR2X1 U527 ( .A(sa23_sr[4]), .B(sa33_sr[4]), .Y(n565) );
  XOR2X1 U667 ( .A(sa22_sr[4]), .B(sa32_sr[4]), .Y(n547) );
  XOR2X1 U947 ( .A(sa20_sr[4]), .B(sa30_sr[4]), .Y(n511) );
  XOR2X1 U814 ( .A(sa01_sr[4]), .B(sa11_sr[4]), .Y(n538) );
  XOR2X1 U534 ( .A(sa03_sr[4]), .B(sa13_sr[4]), .Y(n574) );
  XOR2X1 U674 ( .A(sa02_sr[4]), .B(sa12_sr[4]), .Y(n556) );
  XOR2X1 U954 ( .A(sa00_sr[4]), .B(sa10_sr[4]), .Y(n520) );
  XOR2X1 U949 ( .A(sa00_sr[7]), .B(sa10_sr[7]), .Y(n517) );
  XOR2X1 U809 ( .A(sa01_sr[7]), .B(sa11_sr[7]), .Y(n535) );
  XOR2X1 U824 ( .A(sa21_sr[7]), .B(sa31_sr[7]), .Y(n534) );
  XOR2X1 U529 ( .A(sa03_sr[7]), .B(sa13_sr[7]), .Y(n571) );
  XOR2X1 U544 ( .A(sa23_sr[7]), .B(sa33_sr[7]), .Y(n570) );
  XOR2X1 U669 ( .A(sa02_sr[7]), .B(sa12_sr[7]), .Y(n553) );
  XOR2X1 U684 ( .A(sa22_sr[7]), .B(sa32_sr[7]), .Y(n552) );
  XOR2X1 U964 ( .A(sa20_sr[7]), .B(sa30_sr[7]), .Y(n516) );
  XOR2X1 U793 ( .A(n541), .B(n531), .Y(n250) );
  XOR2X1 U513 ( .A(n577), .B(n567), .Y(n430) );
  XOR2X1 U653 ( .A(n559), .B(n549), .Y(n340) );
  XOR2X1 U933 ( .A(n523), .B(n513), .Y(n160) );
  XOR2X1 U821 ( .A(n534), .B(n536), .Y(n238) );
  XOR2X1 U541 ( .A(n570), .B(n572), .Y(n418) );
  XOR2X1 U681 ( .A(n552), .B(n554), .Y(n328) );
  XOR2X1 U961 ( .A(n516), .B(n518), .Y(n148) );
  XOR2X1 U885 ( .A(n517), .B(n509), .Y(n193) );
  XOR2X1 U465 ( .A(n571), .B(n563), .Y(n463) );
  XOR2X1 U745 ( .A(n535), .B(n527), .Y(n283) );
  XOR2X1 U605 ( .A(n553), .B(n545), .Y(n373) );
  XOR2X1 U816 ( .A(n537), .B(n527), .Y(n240) );
  XOR2X1 U536 ( .A(n573), .B(n563), .Y(n420) );
  XOR2X1 U676 ( .A(n555), .B(n545), .Y(n330) );
  XOR2X1 U956 ( .A(n519), .B(n509), .Y(n150) );
  XOR2X1 U739 ( .A(n537), .B(n529), .Y(n287) );
  XOR2X1 U459 ( .A(n573), .B(n565), .Y(n467) );
  XOR2X1 U599 ( .A(n555), .B(n547), .Y(n377) );
  XOR2X1 U879 ( .A(n519), .B(n511), .Y(n197) );
  XOR2X1 U811 ( .A(n538), .B(n528), .Y(n242) );
  XOR2X1 U531 ( .A(n574), .B(n564), .Y(n422) );
  XOR2X1 U671 ( .A(n556), .B(n546), .Y(n332) );
  XOR2X1 U951 ( .A(n520), .B(n510), .Y(n152) );
  XOR2X1 U728 ( .A(n540), .B(n532), .Y(n295) );
  XOR2X1 U448 ( .A(n576), .B(n568), .Y(n475) );
  XOR2X1 U588 ( .A(n558), .B(n550), .Y(n385) );
  XOR2X1 U868 ( .A(n522), .B(n514), .Y(n205) );
  XOR2X1 U742 ( .A(n536), .B(n528), .Y(n285) );
  XOR2X1 U462 ( .A(n572), .B(n564), .Y(n465) );
  XOR2X1 U602 ( .A(n554), .B(n546), .Y(n375) );
  XOR2X1 U882 ( .A(n518), .B(n510), .Y(n195) );
  XOR2X1 U808 ( .A(sa01_sr[3]), .B(sa11_sr[3]), .Y(n539) );
  XOR2X1 U528 ( .A(sa03_sr[3]), .B(sa13_sr[3]), .Y(n575) );
  XOR2X1 U668 ( .A(sa02_sr[3]), .B(sa12_sr[3]), .Y(n557) );
  XOR2X1 U948 ( .A(sa00_sr[3]), .B(sa10_sr[3]), .Y(n521) );
  XOR2X1 U931 ( .A(sa00_sr[0]), .B(sa10_sr[0]), .Y(n524) );
  XOR2X1 U791 ( .A(sa01_sr[0]), .B(sa11_sr[0]), .Y(n542) );
  XOR2X1 U651 ( .A(sa02_sr[0]), .B(sa12_sr[0]), .Y(n560) );
  XOR2X1 U511 ( .A(sa03_sr[0]), .B(sa13_sr[0]), .Y(n578) );
  DFFHQXL \dcnt_reg[2]  ( .D(n145), .CK(clk), .Q(n866) );
  DFFHQX1 \sa32_reg[4]  ( .D(N100), .CK(clk), .Q(sa32[4]) );
  DFFHQX1 \sa31_reg[4]  ( .D(N164), .CK(clk), .Q(sa31[4]) );
  DFFHQX1 \sa30_reg[4]  ( .D(N228), .CK(clk), .Q(sa30[4]) );
  DFFHQX1 \sa33_reg[4]  ( .D(N36), .CK(clk), .Q(sa33[4]) );
  DFFHQX1 \sa12_reg[4]  ( .D(N132), .CK(clk), .Q(sa12[4]) );
  DFFHQX1 \sa11_reg[4]  ( .D(N196), .CK(clk), .Q(sa11[4]) );
  DFFHQX1 \sa10_reg[4]  ( .D(N260), .CK(clk), .Q(sa10[4]) );
  DFFHQX1 \sa13_reg[4]  ( .D(N68), .CK(clk), .Q(sa13[4]) );
  DFFHQX1 \sa22_reg[4]  ( .D(N116), .CK(clk), .Q(sa22[4]) );
  DFFHQX1 \sa21_reg[4]  ( .D(N180), .CK(clk), .Q(sa21[4]) );
  DFFHQX1 \sa20_reg[4]  ( .D(N244), .CK(clk), .Q(sa20[4]) );
  DFFHQX1 \sa23_reg[4]  ( .D(N52), .CK(clk), .Q(sa23[4]) );
  DFFHQX1 \sa02_reg[4]  ( .D(N148), .CK(clk), .Q(sa02[4]) );
  DFFHQX1 \sa01_reg[4]  ( .D(N212), .CK(clk), .Q(sa01[4]) );
  DFFHQX1 \sa00_reg[4]  ( .D(N276), .CK(clk), .Q(sa00[4]) );
  DFFHQX1 \sa03_reg[4]  ( .D(N84), .CK(clk), .Q(sa03[4]) );
  XOR2X1 U454 ( .A(w3[12]), .B(sa33_sr[4]), .Y(n471) );
  XOR2X1 U1365 ( .A(w3[18]), .B(sa13_sr[2]), .Y(N437) );
  XOR2XL U1366 ( .A(n955), .B(w3[18]), .Y(n754) );
  XOR2X1 U1367 ( .A(w3[28]), .B(sa03_sr[4]), .Y(N403) );
  XOR2XL U1368 ( .A(n921), .B(w3[28]), .Y(n744) );
  XOR2X1 U1369 ( .A(w3[20]), .B(sa13_sr[4]), .Y(N435) );
  XOR2XL U1370 ( .A(n916), .B(w3[20]), .Y(n752) );
  XOR2X1 U1371 ( .A(w3[4]), .B(sa33_sr[4]), .Y(N499) );
  XOR2XL U1372 ( .A(n919), .B(w3[4]), .Y(n768) );
  XOR2XL U1373 ( .A(n918), .B(w3[12]), .Y(n760) );
  XOR2XL U1374 ( .A(n915), .B(w3[19]), .Y(n753) );
  XOR2XL U1375 ( .A(n922), .B(w3[27]), .Y(n745) );
  XOR2XL U1376 ( .A(n917), .B(w3[11]), .Y(n761) );
  XOR2XL U1377 ( .A(n920), .B(w3[3]), .Y(n769) );
  NOR2X1 U1378 ( .A(dcnt[1]), .B(dcnt[0]), .Y(n735) );
  NOR2X1 U1379 ( .A(n729), .B(n866), .Y(n731) );
  NAND2X1 U1380 ( .A(n1009), .B(rst), .Y(n733) );
  INVX1 U1381 ( .A(n735), .Y(n729) );
  CLKINVX3 U1382 ( .A(n996), .Y(n1004) );
  CLKINVX3 U1383 ( .A(n996), .Y(n1001) );
  CLKINVX3 U1384 ( .A(n996), .Y(n997) );
  CLKINVX3 U1385 ( .A(n996), .Y(n1002) );
  CLKINVX3 U1386 ( .A(n1008), .Y(n1000) );
  CLKINVX3 U1387 ( .A(n996), .Y(n998) );
  CLKINVX3 U1388 ( .A(n996), .Y(n1003) );
  CLKINVX3 U1389 ( .A(n1008), .Y(n999) );
  CLKINVX3 U1390 ( .A(n996), .Y(n1005) );
  CLKINVX3 U1391 ( .A(n996), .Y(n1007) );
  CLKINVX3 U1392 ( .A(n996), .Y(n1006) );
  INVX1 U1393 ( .A(n731), .Y(n728) );
  INVX12 U1394 ( .A(n1012), .Y(n1010) );
  INVX12 U1395 ( .A(n1012), .Y(n1011) );
  OAI2BB2X1 U1396 ( .B0(n6), .B1(n798), .A0N(sa30_next[6]), .A1N(n1007), .Y(
        N230) );
  XOR2X1 U1397 ( .A(n867), .B(w0[6]), .Y(n798) );
  OAI2BB2X1 U1398 ( .B0(n999), .B1(n774), .A0N(sa00_next[6]), .A1N(n1006), .Y(
        N278) );
  XOR2X1 U1399 ( .A(n869), .B(w0[30]), .Y(n774) );
  OAI2BB2X1 U1400 ( .B0(n1000), .B1(n790), .A0N(sa20_next[6]), .A1N(n1007), 
        .Y(N246) );
  XOR2X1 U1401 ( .A(n870), .B(w0[14]), .Y(n790) );
  OAI2BB2X1 U1402 ( .B0(n1001), .B1(n863), .A0N(sa32_next[6]), .A1N(n1004), 
        .Y(N102) );
  XOR2X1 U1403 ( .A(n872), .B(w2[6]), .Y(n863) );
  OAI2BB2X1 U1404 ( .B0(n1001), .B1(n855), .A0N(sa22_next[6]), .A1N(n1005), 
        .Y(N118) );
  XOR2X1 U1405 ( .A(n873), .B(w2[14]), .Y(n855) );
  OAI2BB2X1 U1406 ( .B0(n1003), .B1(n839), .A0N(sa02_next[6]), .A1N(n1007), 
        .Y(N150) );
  XOR2X1 U1407 ( .A(n874), .B(w2[30]), .Y(n839) );
  OAI2BB2X1 U1408 ( .B0(n1002), .B1(n831), .A0N(sa31_next[6]), .A1N(n1007), 
        .Y(N166) );
  XOR2X1 U1409 ( .A(n880), .B(w1[6]), .Y(n831) );
  OAI2BB2X1 U1410 ( .B0(n1001), .B1(n823), .A0N(sa21_next[6]), .A1N(n1002), 
        .Y(N182) );
  XOR2X1 U1411 ( .A(n881), .B(w1[14]), .Y(n823) );
  OAI2BB2X1 U1412 ( .B0(n6), .B1(n806), .A0N(sa01_next[6]), .A1N(n1002), .Y(
        N214) );
  XOR2X1 U1413 ( .A(n882), .B(w1[30]), .Y(n806) );
  OAI2BB2X1 U1414 ( .B0(n1000), .B1(n795), .A0N(sa20_next[1]), .A1N(n1007), 
        .Y(N241) );
  XOR2X1 U1415 ( .A(n883), .B(w0[9]), .Y(n795) );
  OAI2BB2X1 U1416 ( .B0(n1000), .B1(n787), .A0N(sa10_next[1]), .A1N(n1007), 
        .Y(N257) );
  XOR2X1 U1417 ( .A(n885), .B(w0[17]), .Y(n787) );
  OAI2BB2X1 U1418 ( .B0(n999), .B1(n779), .A0N(sa00_next[1]), .A1N(n1006), .Y(
        N273) );
  XOR2X1 U1419 ( .A(n886), .B(w0[25]), .Y(n779) );
  OAI2BB2X1 U1420 ( .B0(n1002), .B1(n852), .A0N(sa12_next[1]), .A1N(n1006), 
        .Y(N129) );
  XOR2X1 U1421 ( .A(n887), .B(w2[17]), .Y(n852) );
  OAI2BB2X1 U1422 ( .B0(n1002), .B1(n860), .A0N(sa22_next[1]), .A1N(n1004), 
        .Y(N113) );
  XOR2X1 U1423 ( .A(n889), .B(w2[9]), .Y(n860) );
  OAI2BB2X1 U1424 ( .B0(n1004), .B1(n844), .A0N(sa02_next[1]), .A1N(n1006), 
        .Y(N145) );
  XOR2X1 U1425 ( .A(n890), .B(w2[25]), .Y(n844) );
  OAI2BB2X1 U1426 ( .B0(n1002), .B1(n828), .A0N(sa21_next[1]), .A1N(n1002), 
        .Y(N177) );
  XOR2X1 U1427 ( .A(n895), .B(w1[9]), .Y(n828) );
  OAI2BB2X1 U1428 ( .B0(n997), .B1(n812), .A0N(sa01_next[1]), .A1N(n1001), .Y(
        N209) );
  XOR2X1 U1429 ( .A(n896), .B(w1[25]), .Y(n812) );
  OAI2BB2X1 U1430 ( .B0(n998), .B1(n820), .A0N(sa11_next[1]), .A1N(n1002), .Y(
        N193) );
  XOR2X1 U1431 ( .A(n897), .B(w1[17]), .Y(n820) );
  OAI2BB2X1 U1432 ( .B0(n1000), .B1(n793), .A0N(sa20_next[3]), .A1N(n1007), 
        .Y(N243) );
  XOR2X1 U1433 ( .A(n899), .B(w0[11]), .Y(n793) );
  OAI2BB2X1 U1434 ( .B0(n6), .B1(n800), .A0N(sa30_next[4]), .A1N(n1007), .Y(
        N228) );
  XOR2X1 U1435 ( .A(n901), .B(w0[4]), .Y(n800) );
  OAI2BB2X1 U1436 ( .B0(n999), .B1(n784), .A0N(sa10_next[4]), .A1N(n1006), .Y(
        N260) );
  XOR2X1 U1437 ( .A(n902), .B(w0[20]), .Y(n784) );
  OAI2BB2X1 U1438 ( .B0(n999), .B1(n785), .A0N(sa10_next[3]), .A1N(n1007), .Y(
        N259) );
  XOR2X1 U1439 ( .A(n905), .B(w0[19]), .Y(n785) );
  OAI2BB2X1 U1440 ( .B0(n999), .B1(n777), .A0N(sa00_next[3]), .A1N(n1006), .Y(
        N275) );
  XOR2X1 U1441 ( .A(n906), .B(w0[27]), .Y(n777) );
  OAI2BB2X1 U1442 ( .B0(n1002), .B1(n849), .A0N(sa12_next[4]), .A1N(n1006), 
        .Y(N132) );
  XOR2X1 U1443 ( .A(n907), .B(w2[20]), .Y(n849) );
  OAI2BB2X1 U1444 ( .B0(n1001), .B1(n865), .A0N(sa32_next[4]), .A1N(n1006), 
        .Y(N100) );
  XOR2X1 U1445 ( .A(n908), .B(w2[4]), .Y(n865) );
  OAI2BB2X1 U1446 ( .B0(n1004), .B1(n850), .A0N(sa12_next[3]), .A1N(n1006), 
        .Y(N131) );
  XOR2X1 U1447 ( .A(n910), .B(w2[19]), .Y(n850) );
  OAI2BB2X1 U1448 ( .B0(n1001), .B1(n858), .A0N(sa22_next[3]), .A1N(n1005), 
        .Y(N115) );
  XOR2X1 U1449 ( .A(n912), .B(w2[11]), .Y(n858) );
  OAI2BB2X1 U1450 ( .B0(n1004), .B1(n842), .A0N(sa02_next[3]), .A1N(n1006), 
        .Y(N147) );
  XOR2X1 U1451 ( .A(n914), .B(w2[27]), .Y(n842) );
  OAI2BB2X1 U1452 ( .B0(n1001), .B1(n826), .A0N(sa21_next[3]), .A1N(n1001), 
        .Y(N179) );
  XOR2X1 U1453 ( .A(n923), .B(w1[11]), .Y(n826) );
  OAI2BB2X1 U1454 ( .B0(n6), .B1(n809), .A0N(sa01_next[3]), .A1N(n1001), .Y(
        N211) );
  XOR2X1 U1455 ( .A(n925), .B(w1[27]), .Y(n809) );
  OAI2BB2X1 U1456 ( .B0(n997), .B1(n817), .A0N(sa11_next[4]), .A1N(n1002), .Y(
        N196) );
  XOR2X1 U1457 ( .A(n927), .B(w1[20]), .Y(n817) );
  OAI2BB2X1 U1458 ( .B0(n1003), .B1(n833), .A0N(sa31_next[4]), .A1N(n1007), 
        .Y(N164) );
  XOR2X1 U1459 ( .A(n928), .B(w1[4]), .Y(n833) );
  OAI2BB2X1 U1460 ( .B0(n998), .B1(n818), .A0N(sa11_next[3]), .A1N(n1001), .Y(
        N195) );
  XOR2X1 U1461 ( .A(n929), .B(w1[19]), .Y(n818) );
  OAI2BB2X1 U1462 ( .B0(n1002), .B1(n862), .A0N(sa32_next[7]), .A1N(n1005), 
        .Y(N103) );
  XOR2X1 U1463 ( .A(n931), .B(w2[7]), .Y(n862) );
  OAI2BB2X1 U1464 ( .B0(n1000), .B1(n797), .A0N(sa30_next[7]), .A1N(n1007), 
        .Y(N231) );
  XOR2X1 U1465 ( .A(n932), .B(w0[7]), .Y(n797) );
  OAI2BB2X1 U1466 ( .B0(n999), .B1(n781), .A0N(sa10_next[7]), .A1N(n1006), .Y(
        N263) );
  XOR2X1 U1467 ( .A(n933), .B(w0[23]), .Y(n781) );
  OAI2BB2X1 U1468 ( .B0(n998), .B1(n773), .A0N(sa00_next[7]), .A1N(n1006), .Y(
        N279) );
  XOR2X1 U1469 ( .A(n934), .B(w0[31]), .Y(n773) );
  OAI2BB2X1 U1470 ( .B0(n1003), .B1(n854), .A0N(sa22_next[7]), .A1N(n1005), 
        .Y(N119) );
  XOR2X1 U1471 ( .A(n935), .B(w2[15]), .Y(n854) );
  OAI2BB2X1 U1472 ( .B0(n1004), .B1(n846), .A0N(sa12_next[7]), .A1N(n1006), 
        .Y(N135) );
  XOR2X1 U1473 ( .A(n936), .B(w2[23]), .Y(n846) );
  OAI2BB2X1 U1474 ( .B0(n1003), .B1(n838), .A0N(sa02_next[7]), .A1N(n1007), 
        .Y(N151) );
  XOR2X1 U1475 ( .A(n937), .B(w2[31]), .Y(n838) );
  OAI2BB2X1 U1476 ( .B0(n1002), .B1(n830), .A0N(sa31_next[7]), .A1N(n1001), 
        .Y(N167) );
  XOR2X1 U1477 ( .A(n939), .B(w1[7]), .Y(n830) );
  OAI2BB2X1 U1478 ( .B0(n997), .B1(n814), .A0N(sa11_next[7]), .A1N(n1007), .Y(
        N199) );
  XOR2X1 U1479 ( .A(n942), .B(w1[23]), .Y(n814) );
  OAI2BB2X1 U1480 ( .B0(n999), .B1(n822), .A0N(sa21_next[7]), .A1N(n1004), .Y(
        N183) );
  XOR2X1 U1481 ( .A(n943), .B(w1[15]), .Y(n822) );
  OAI2BB2X1 U1482 ( .B0(n6), .B1(n805), .A0N(sa01_next[7]), .A1N(n1007), .Y(
        N215) );
  XOR2X1 U1483 ( .A(n944), .B(w1[31]), .Y(n805) );
  OAI2BB2X1 U1484 ( .B0(n1000), .B1(n789), .A0N(sa20_next[7]), .A1N(n1007), 
        .Y(N247) );
  XOR2X1 U1485 ( .A(n946), .B(w0[15]), .Y(n789) );
  OAI2BB2X1 U1486 ( .B0(n6), .B1(n802), .A0N(sa30_next[2]), .A1N(n1007), .Y(
        N226) );
  XOR2X1 U1487 ( .A(n947), .B(w0[2]), .Y(n802) );
  OAI2BB2X1 U1488 ( .B0(n999), .B1(n778), .A0N(sa00_next[2]), .A1N(n1006), .Y(
        N274) );
  XOR2X1 U1489 ( .A(n949), .B(w0[26]), .Y(n778) );
  OAI2BB2X1 U1490 ( .B0(n1000), .B1(n794), .A0N(sa20_next[2]), .A1N(n1007), 
        .Y(N242) );
  XOR2X1 U1491 ( .A(n950), .B(w0[10]), .Y(n794) );
  OAI2BB2X1 U1492 ( .B0(n1002), .B1(n738), .A0N(sa32_next[2]), .A1N(n1005), 
        .Y(N98) );
  XOR2X1 U1493 ( .A(n952), .B(w2[2]), .Y(n738) );
  OAI2BB2X1 U1494 ( .B0(n1002), .B1(n859), .A0N(sa22_next[2]), .A1N(n1005), 
        .Y(N114) );
  XOR2X1 U1495 ( .A(n953), .B(w2[10]), .Y(n859) );
  OAI2BB2X1 U1496 ( .B0(n1004), .B1(n843), .A0N(sa02_next[2]), .A1N(n1006), 
        .Y(N146) );
  XOR2X1 U1497 ( .A(n954), .B(w2[26]), .Y(n843) );
  OAI2BB2X1 U1498 ( .B0(n1003), .B1(n835), .A0N(sa31_next[2]), .A1N(n1007), 
        .Y(N162) );
  XOR2X1 U1499 ( .A(n960), .B(w1[2]), .Y(n835) );
  OAI2BB2X1 U1500 ( .B0(n1001), .B1(n827), .A0N(sa21_next[2]), .A1N(n1007), 
        .Y(N178) );
  XOR2X1 U1501 ( .A(n961), .B(w1[10]), .Y(n827) );
  OAI2BB2X1 U1502 ( .B0(n999), .B1(n810), .A0N(sa01_next[2]), .A1N(n1007), .Y(
        N210) );
  XOR2X1 U1503 ( .A(n962), .B(w1[26]), .Y(n810) );
  OAI2BB2X1 U1504 ( .B0(n999), .B1(n783), .A0N(sa10_next[5]), .A1N(n1006), .Y(
        N261) );
  XOR2X1 U1505 ( .A(n964), .B(w0[21]), .Y(n783) );
  OAI2BB2X1 U1506 ( .B0(n999), .B1(n775), .A0N(sa00_next[5]), .A1N(n1006), .Y(
        N277) );
  XOR2X1 U1507 ( .A(n965), .B(w0[29]), .Y(n775) );
  OAI2BB2X1 U1508 ( .B0(n1000), .B1(n791), .A0N(sa20_next[5]), .A1N(n1007), 
        .Y(N245) );
  XOR2X1 U1509 ( .A(n966), .B(w0[13]), .Y(n791) );
  OAI2BB2X1 U1510 ( .B0(n1004), .B1(n848), .A0N(sa12_next[5]), .A1N(n1006), 
        .Y(N133) );
  XOR2X1 U1511 ( .A(n967), .B(w2[21]), .Y(n848) );
  OAI2BB2X1 U1512 ( .B0(n1003), .B1(n856), .A0N(sa22_next[5]), .A1N(n1005), 
        .Y(N117) );
  XOR2X1 U1513 ( .A(n969), .B(w2[13]), .Y(n856) );
  OAI2BB2X1 U1514 ( .B0(n1003), .B1(n840), .A0N(sa02_next[5]), .A1N(n1007), 
        .Y(N149) );
  XOR2X1 U1515 ( .A(n970), .B(w2[29]), .Y(n840) );
  OAI2BB2X1 U1516 ( .B0(n6), .B1(n816), .A0N(sa11_next[5]), .A1N(n1001), .Y(
        N197) );
  XOR2X1 U1517 ( .A(n975), .B(w1[21]), .Y(n816) );
  OAI2BB2X1 U1518 ( .B0(n1001), .B1(n824), .A0N(sa21_next[5]), .A1N(n1002), 
        .Y(N181) );
  XOR2X1 U1519 ( .A(n977), .B(w1[13]), .Y(n824) );
  OAI2BB2X1 U1520 ( .B0(n6), .B1(n807), .A0N(sa01_next[5]), .A1N(n997), .Y(
        N213) );
  XOR2X1 U1521 ( .A(n978), .B(w1[29]), .Y(n807) );
  OAI2BB2X1 U1522 ( .B0(n1000), .B1(n796), .A0N(sa20_next[0]), .A1N(n1007), 
        .Y(N240) );
  XOR2X1 U1523 ( .A(n979), .B(w0[8]), .Y(n796) );
  OAI2BB2X1 U1524 ( .B0(n1002), .B1(n861), .A0N(sa22_next[0]), .A1N(n1004), 
        .Y(N112) );
  XOR2X1 U1525 ( .A(n980), .B(w2[8]), .Y(n861) );
  OAI2BB2X1 U1526 ( .B0(n1002), .B1(n845), .A0N(sa02_next[0]), .A1N(n1006), 
        .Y(N144) );
  XOR2X1 U1527 ( .A(n981), .B(w2[24]), .Y(n845) );
  OAI2BB2X1 U1528 ( .B0(n1002), .B1(n829), .A0N(sa21_next[0]), .A1N(n1000), 
        .Y(N176) );
  XOR2X1 U1529 ( .A(n985), .B(w1[8]), .Y(n829) );
  OAI2BB2X1 U1530 ( .B0(n1000), .B1(n813), .A0N(sa01_next[0]), .A1N(n997), .Y(
        N208) );
  XOR2X1 U1531 ( .A(n986), .B(w1[24]), .Y(n813) );
  OAI2BB2X1 U1532 ( .B0(n1000), .B1(n788), .A0N(sa10_next[0]), .A1N(n1007), 
        .Y(N256) );
  XOR2X1 U1533 ( .A(n987), .B(w0[16]), .Y(n788) );
  OAI2BB2X1 U1534 ( .B0(n999), .B1(n821), .A0N(sa11_next[0]), .A1N(n998), .Y(
        N192) );
  XOR2X1 U1535 ( .A(n988), .B(w1[16]), .Y(n821) );
  OAI2BB2X1 U1536 ( .B0(n1003), .B1(n853), .A0N(sa12_next[0]), .A1N(n1005), 
        .Y(N128) );
  XOR2X1 U1537 ( .A(n989), .B(w2[16]), .Y(n853) );
  OAI2BB2X1 U1538 ( .B0(n1001), .B1(n740), .A0N(sa32_next[0]), .A1N(n1004), 
        .Y(N96) );
  XOR2X1 U1539 ( .A(n991), .B(w2[0]), .Y(n740) );
  OAI2BB2X1 U1540 ( .B0(n1003), .B1(n837), .A0N(sa31_next[0]), .A1N(n1007), 
        .Y(N160) );
  XOR2X1 U1541 ( .A(n992), .B(w1[0]), .Y(n837) );
  OAI2BB2X1 U1542 ( .B0(n6), .B1(n804), .A0N(sa30_next[0]), .A1N(n1007), .Y(
        N224) );
  XOR2X1 U1543 ( .A(n993), .B(w0[0]), .Y(n804) );
  OAI2BB2X1 U1544 ( .B0(n999), .B1(n780), .A0N(sa00_next[0]), .A1N(n1006), .Y(
        N272) );
  XOR2X1 U1545 ( .A(n994), .B(w0[24]), .Y(n780) );
  OAI2BB2X1 U1546 ( .B0(n997), .B1(n750), .A0N(sa13_next[6]), .A1N(n1005), .Y(
        N70) );
  XOR2X1 U1547 ( .A(n875), .B(w3[22]), .Y(n750) );
  OAI2BB2X1 U1548 ( .B0(n998), .B1(n766), .A0N(sa33_next[6]), .A1N(n1006), .Y(
        N38) );
  XOR2X1 U1549 ( .A(n876), .B(w3[6]), .Y(n766) );
  OAI2BB2X1 U1550 ( .B0(n997), .B1(n758), .A0N(sa23_next[6]), .A1N(n1005), .Y(
        N54) );
  XOR2X1 U1551 ( .A(n877), .B(w3[14]), .Y(n758) );
  OAI2BB2X1 U1552 ( .B0(n1002), .B1(n742), .A0N(sa03_next[6]), .A1N(n1004), 
        .Y(N86) );
  XOR2X1 U1553 ( .A(n878), .B(w3[30]), .Y(n742) );
  OAI2BB2X1 U1554 ( .B0(n997), .B1(n755), .A0N(sa13_next[1]), .A1N(n1005), .Y(
        N65) );
  XOR2X1 U1555 ( .A(n891), .B(w3[17]), .Y(n755) );
  OAI2BB2X1 U1556 ( .B0(n998), .B1(n763), .A0N(sa23_next[1]), .A1N(n1005), .Y(
        N49) );
  XOR2X1 U1557 ( .A(n892), .B(w3[9]), .Y(n763) );
  OAI2BB2X1 U1558 ( .B0(n1000), .B1(n747), .A0N(sa03_next[1]), .A1N(n1005), 
        .Y(N81) );
  XOR2X1 U1559 ( .A(n894), .B(w3[25]), .Y(n747) );
  OAI2BB2X1 U1560 ( .B0(n997), .B1(n751), .A0N(sa13_next[5]), .A1N(n1005), .Y(
        N69) );
  XOR2X1 U1561 ( .A(n971), .B(w3[21]), .Y(n751) );
  OAI2BB2X1 U1562 ( .B0(n998), .B1(n767), .A0N(sa33_next[5]), .A1N(n1006), .Y(
        N37) );
  XOR2X1 U1563 ( .A(n972), .B(w3[5]), .Y(n767) );
  OAI2BB2X1 U1564 ( .B0(n997), .B1(n759), .A0N(sa23_next[5]), .A1N(n1005), .Y(
        N53) );
  XOR2X1 U1565 ( .A(n973), .B(w3[13]), .Y(n759) );
  OAI2BB2X1 U1566 ( .B0(n6), .B1(n743), .A0N(sa03_next[5]), .A1N(n1004), .Y(
        N85) );
  XOR2X1 U1567 ( .A(n974), .B(w3[29]), .Y(n743) );
  OAI2BB2X1 U1568 ( .B0(n998), .B1(n765), .A0N(sa33_next[7]), .A1N(n1006), .Y(
        N39) );
  XOR2X1 U1569 ( .A(n938), .B(w3[7]), .Y(n765) );
  OAI2BB2X1 U1570 ( .B0(n997), .B1(n749), .A0N(sa13_next[7]), .A1N(n1005), .Y(
        N71) );
  XOR2X1 U1571 ( .A(n940), .B(w3[23]), .Y(n749) );
  OAI2BB2X1 U1572 ( .B0(n998), .B1(n741), .A0N(sa03_next[7]), .A1N(n1005), .Y(
        N87) );
  XOR2X1 U1573 ( .A(n941), .B(w3[31]), .Y(n741) );
  OAI2BB2X1 U1574 ( .B0(n997), .B1(n757), .A0N(sa23_next[7]), .A1N(n1005), .Y(
        N55) );
  XOR2X1 U1575 ( .A(n945), .B(w3[15]), .Y(n757) );
  OAI2BB2X1 U1576 ( .B0(n997), .B1(n753), .A0N(sa13_next[3]), .A1N(n1005), .Y(
        N67) );
  OAI2BB2X1 U1577 ( .B0(n997), .B1(n752), .A0N(sa13_next[4]), .A1N(n1005), .Y(
        N68) );
  OAI2BB2X1 U1578 ( .B0(n997), .B1(n761), .A0N(sa23_next[3]), .A1N(n1005), .Y(
        N51) );
  OAI2BB2X1 U1579 ( .B0(n998), .B1(n768), .A0N(sa33_next[4]), .A1N(n1006), .Y(
        N36) );
  OAI2BB2X1 U1580 ( .B0(n1003), .B1(n745), .A0N(sa03_next[3]), .A1N(n1004), 
        .Y(N83) );
  OAI2BB2X1 U1581 ( .B0(n998), .B1(n770), .A0N(sa33_next[2]), .A1N(n1006), .Y(
        N34) );
  XOR2X1 U1582 ( .A(n956), .B(w3[2]), .Y(n770) );
  OAI2BB2X1 U1583 ( .B0(n998), .B1(n762), .A0N(sa23_next[2]), .A1N(n1005), .Y(
        N50) );
  XOR2X1 U1584 ( .A(n957), .B(w3[10]), .Y(n762) );
  OAI2BB2X1 U1585 ( .B0(n998), .B1(n746), .A0N(sa03_next[2]), .A1N(n1004), .Y(
        N82) );
  XOR2X1 U1586 ( .A(n958), .B(w3[26]), .Y(n746) );
  OAI2BB2X1 U1587 ( .B0(n997), .B1(n756), .A0N(sa13_next[0]), .A1N(n1005), .Y(
        N64) );
  XOR2X1 U1588 ( .A(n982), .B(w3[16]), .Y(n756) );
  OAI2BB2X1 U1589 ( .B0(n998), .B1(n764), .A0N(sa23_next[0]), .A1N(n1005), .Y(
        N48) );
  XOR2X1 U1590 ( .A(n983), .B(w3[8]), .Y(n764) );
  OAI2BB2X1 U1591 ( .B0(n999), .B1(n748), .A0N(sa03_next[0]), .A1N(n1005), .Y(
        N80) );
  XOR2X1 U1592 ( .A(n984), .B(w3[24]), .Y(n748) );
  OAI2BB2X1 U1593 ( .B0(n998), .B1(n772), .A0N(sa33_next[0]), .A1N(n1006), .Y(
        N32) );
  XOR2X1 U1594 ( .A(n990), .B(w3[0]), .Y(n772) );
  OAI2BB2X1 U1595 ( .B0(n999), .B1(n782), .A0N(sa10_next[6]), .A1N(n1006), .Y(
        N262) );
  XOR2X1 U1596 ( .A(n868), .B(w0[22]), .Y(n782) );
  OAI2BB2X1 U1597 ( .B0(n1004), .B1(n847), .A0N(sa12_next[6]), .A1N(n1006), 
        .Y(N134) );
  XOR2X1 U1598 ( .A(n871), .B(w2[22]), .Y(n847) );
  OAI2BB2X1 U1599 ( .B0(n6), .B1(n815), .A0N(sa11_next[6]), .A1N(n1003), .Y(
        N198) );
  XOR2X1 U1600 ( .A(n879), .B(w1[22]), .Y(n815) );
  OAI2BB2X1 U1601 ( .B0(n6), .B1(n803), .A0N(sa30_next[1]), .A1N(n1007), .Y(
        N225) );
  XOR2X1 U1602 ( .A(n884), .B(w0[1]), .Y(n803) );
  OAI2BB2X1 U1603 ( .B0(n1000), .B1(n739), .A0N(sa32_next[1]), .A1N(n1005), 
        .Y(N97) );
  XOR2X1 U1604 ( .A(n888), .B(w2[1]), .Y(n739) );
  OAI2BB2X1 U1605 ( .B0(n998), .B1(n771), .A0N(sa33_next[1]), .A1N(n1006), .Y(
        N33) );
  XOR2X1 U1606 ( .A(n893), .B(w3[1]), .Y(n771) );
  OAI2BB2X1 U1607 ( .B0(n1001), .B1(n836), .A0N(sa31_next[1]), .A1N(n1007), 
        .Y(N161) );
  XOR2X1 U1608 ( .A(n898), .B(w1[1]), .Y(n836) );
  OAI2BB2X1 U1609 ( .B0(n1000), .B1(n792), .A0N(sa20_next[4]), .A1N(n1007), 
        .Y(N244) );
  XOR2X1 U1610 ( .A(n900), .B(w0[12]), .Y(n792) );
  OAI2BB2X1 U1611 ( .B0(n999), .B1(n776), .A0N(sa00_next[4]), .A1N(n1006), .Y(
        N276) );
  XOR2X1 U1612 ( .A(n903), .B(w0[28]), .Y(n776) );
  OAI2BB2X1 U1613 ( .B0(n1001), .B1(n801), .A0N(sa30_next[3]), .A1N(n1007), 
        .Y(N227) );
  XOR2X1 U1614 ( .A(n904), .B(w0[3]), .Y(n801) );
  OAI2BB2X1 U1615 ( .B0(n1003), .B1(n857), .A0N(sa22_next[4]), .A1N(n1005), 
        .Y(N116) );
  XOR2X1 U1616 ( .A(n909), .B(w2[12]), .Y(n857) );
  OAI2BB2X1 U1617 ( .B0(n6), .B1(n737), .A0N(sa32_next[3]), .A1N(n1004), .Y(
        N99) );
  XOR2X1 U1618 ( .A(n911), .B(w2[3]), .Y(n737) );
  OAI2BB2X1 U1619 ( .B0(n1003), .B1(n841), .A0N(sa02_next[4]), .A1N(n1007), 
        .Y(N148) );
  XOR2X1 U1620 ( .A(n913), .B(w2[28]), .Y(n841) );
  OAI2BB2X1 U1621 ( .B0(n997), .B1(n760), .A0N(sa23_next[4]), .A1N(n1005), .Y(
        N52) );
  OAI2BB2X1 U1622 ( .B0(n998), .B1(n769), .A0N(sa33_next[3]), .A1N(n1006), .Y(
        N35) );
  OAI2BB2X1 U1623 ( .B0(n6), .B1(n744), .A0N(sa03_next[4]), .A1N(n1005), .Y(
        N84) );
  OAI2BB2X1 U1624 ( .B0(n1001), .B1(n825), .A0N(sa21_next[4]), .A1N(n1000), 
        .Y(N180) );
  XOR2X1 U1625 ( .A(n924), .B(w1[12]), .Y(n825) );
  OAI2BB2X1 U1626 ( .B0(n6), .B1(n808), .A0N(sa01_next[4]), .A1N(n999), .Y(
        N212) );
  XOR2X1 U1627 ( .A(n926), .B(w1[28]), .Y(n808) );
  OAI2BB2X1 U1628 ( .B0(n1003), .B1(n834), .A0N(sa31_next[3]), .A1N(n1007), 
        .Y(N163) );
  XOR2X1 U1629 ( .A(n930), .B(w1[3]), .Y(n834) );
  OAI2BB2X1 U1630 ( .B0(n1000), .B1(n786), .A0N(sa10_next[2]), .A1N(n1007), 
        .Y(N258) );
  XOR2X1 U1631 ( .A(n948), .B(w0[18]), .Y(n786) );
  OAI2BB2X1 U1632 ( .B0(n1004), .B1(n851), .A0N(sa12_next[2]), .A1N(n1005), 
        .Y(N130) );
  XOR2X1 U1633 ( .A(n951), .B(w2[18]), .Y(n851) );
  OAI2BB2X1 U1634 ( .B0(n997), .B1(n754), .A0N(sa13_next[2]), .A1N(n1005), .Y(
        N66) );
  OAI2BB2X1 U1635 ( .B0(n1000), .B1(n819), .A0N(sa11_next[2]), .A1N(n1001), 
        .Y(N194) );
  XOR2X1 U1636 ( .A(n959), .B(w1[18]), .Y(n819) );
  OAI2BB2X1 U1637 ( .B0(n6), .B1(n799), .A0N(sa30_next[5]), .A1N(n1007), .Y(
        N229) );
  XOR2X1 U1638 ( .A(n963), .B(w0[5]), .Y(n799) );
  OAI2BB2X1 U1639 ( .B0(n1001), .B1(n864), .A0N(sa32_next[5]), .A1N(n1004), 
        .Y(N101) );
  XOR2X1 U1640 ( .A(n968), .B(w2[5]), .Y(n864) );
  OAI2BB2X1 U1641 ( .B0(n1002), .B1(n832), .A0N(sa31_next[5]), .A1N(n1007), 
        .Y(N165) );
  XOR2X1 U1642 ( .A(n976), .B(w1[5]), .Y(n832) );
  XOR2X1 U1643 ( .A(w3[3]), .B(sa33_sr[3]), .Y(N500) );
  XOR2X1 U1644 ( .A(w3[11]), .B(sa23_sr[3]), .Y(N468) );
  XOR2X1 U1645 ( .A(w3[19]), .B(sa13_sr[3]), .Y(N436) );
  XOR2X1 U1646 ( .A(w3[27]), .B(sa03_sr[3]), .Y(N404) );
  XOR2XL U1647 ( .A(w3[0]), .B(sa33_sr[0]), .Y(N503) );
  XOR2XL U1648 ( .A(w3[8]), .B(sa23_sr[0]), .Y(N471) );
  XOR2XL U1649 ( .A(w3[16]), .B(sa13_sr[0]), .Y(N439) );
  XOR2XL U1650 ( .A(w3[24]), .B(sa03_sr[0]), .Y(N407) );
  XOR2X1 U1651 ( .A(w3[12]), .B(sa23_sr[4]), .Y(N467) );
  XOR2XL U1652 ( .A(w3[2]), .B(sa33_sr[2]), .Y(N501) );
  XOR2X1 U1653 ( .A(w3[10]), .B(sa23_sr[2]), .Y(N469) );
  XOR2XL U1654 ( .A(w3[26]), .B(sa03_sr[2]), .Y(N405) );
  XOR2XL U1655 ( .A(w2[0]), .B(sa32_sr[0]), .Y(N495) );
  XOR2XL U1656 ( .A(w1[0]), .B(sa31_sr[0]), .Y(N487) );
  XOR2XL U1657 ( .A(w0[0]), .B(sa30_sr[0]), .Y(N479) );
  XOR2XL U1658 ( .A(w2[2]), .B(sa32_sr[2]), .Y(N493) );
  XOR2XL U1659 ( .A(w2[4]), .B(sa32_sr[4]), .Y(N491) );
  XOR2XL U1660 ( .A(w1[2]), .B(sa31_sr[2]), .Y(N485) );
  XOR2XL U1661 ( .A(w1[4]), .B(sa31_sr[4]), .Y(N483) );
  XOR2XL U1662 ( .A(w0[2]), .B(sa30_sr[2]), .Y(N477) );
  XOR2XL U1663 ( .A(w0[4]), .B(sa30_sr[4]), .Y(N475) );
  XOR2XL U1664 ( .A(w2[8]), .B(sa22_sr[0]), .Y(N463) );
  XOR2XL U1665 ( .A(w1[8]), .B(sa21_sr[0]), .Y(N455) );
  XOR2XL U1666 ( .A(w0[8]), .B(sa20_sr[0]), .Y(N447) );
  XOR2XL U1667 ( .A(w2[16]), .B(sa12_sr[0]), .Y(N431) );
  XOR2XL U1668 ( .A(w1[16]), .B(sa11_sr[0]), .Y(N423) );
  XOR2XL U1669 ( .A(w0[16]), .B(sa10_sr[0]), .Y(N415) );
  XOR2XL U1670 ( .A(w2[24]), .B(sa02_sr[0]), .Y(N399) );
  XOR2XL U1671 ( .A(w1[24]), .B(sa01_sr[0]), .Y(N391) );
  XOR2XL U1672 ( .A(w0[24]), .B(sa00_sr[0]), .Y(N383) );
  XOR2XL U1673 ( .A(w2[18]), .B(sa12_sr[2]), .Y(N429) );
  XOR2XL U1674 ( .A(w2[20]), .B(sa12_sr[4]), .Y(N427) );
  XOR2XL U1675 ( .A(w1[18]), .B(sa11_sr[2]), .Y(N421) );
  XOR2XL U1676 ( .A(w1[20]), .B(sa11_sr[4]), .Y(N419) );
  XOR2XL U1677 ( .A(w0[18]), .B(sa10_sr[2]), .Y(N413) );
  XOR2XL U1678 ( .A(w0[20]), .B(sa10_sr[4]), .Y(N411) );
  XOR2XL U1679 ( .A(w2[26]), .B(sa02_sr[2]), .Y(N397) );
  XOR2XL U1680 ( .A(w2[28]), .B(sa02_sr[4]), .Y(N395) );
  XOR2XL U1681 ( .A(w1[26]), .B(sa01_sr[2]), .Y(N389) );
  XOR2XL U1682 ( .A(w1[28]), .B(sa01_sr[4]), .Y(N387) );
  XOR2XL U1683 ( .A(w0[26]), .B(sa00_sr[2]), .Y(N381) );
  XOR2XL U1684 ( .A(w0[28]), .B(sa00_sr[4]), .Y(N379) );
  XOR2XL U1685 ( .A(w3[6]), .B(sa33_sr[6]), .Y(N497) );
  XOR2XL U1686 ( .A(w2[6]), .B(sa32_sr[6]), .Y(N489) );
  XOR2XL U1687 ( .A(w1[6]), .B(sa31_sr[6]), .Y(N481) );
  XOR2XL U1688 ( .A(w0[6]), .B(sa30_sr[6]), .Y(N473) );
  XOR2XL U1689 ( .A(w3[7]), .B(sa33_sr[7]), .Y(N496) );
  XOR2XL U1690 ( .A(w2[7]), .B(sa32_sr[7]), .Y(N488) );
  XOR2XL U1691 ( .A(w1[7]), .B(sa31_sr[7]), .Y(N480) );
  XOR2XL U1692 ( .A(w0[7]), .B(sa30_sr[7]), .Y(N472) );
  XOR2X1 U1693 ( .A(w3[15]), .B(sa23_sr[7]), .Y(N464) );
  XOR2X1 U1694 ( .A(w3[23]), .B(sa13_sr[7]), .Y(N432) );
  XOR2X1 U1695 ( .A(w3[31]), .B(sa03_sr[7]), .Y(N400) );
  XOR2X1 U1696 ( .A(w2[10]), .B(sa22_sr[2]), .Y(N461) );
  XOR2X1 U1697 ( .A(w2[12]), .B(sa22_sr[4]), .Y(N459) );
  XOR2X1 U1698 ( .A(w1[10]), .B(sa21_sr[2]), .Y(N453) );
  XOR2X1 U1699 ( .A(w1[12]), .B(sa21_sr[4]), .Y(N451) );
  XOR2X1 U1700 ( .A(w0[10]), .B(sa20_sr[2]), .Y(N445) );
  XOR2X1 U1701 ( .A(w0[12]), .B(sa20_sr[4]), .Y(N443) );
  XOR2X1 U1702 ( .A(w3[22]), .B(sa13_sr[6]), .Y(N433) );
  XOR2X1 U1703 ( .A(w2[22]), .B(sa12_sr[6]), .Y(N425) );
  XOR2X1 U1704 ( .A(w1[22]), .B(sa11_sr[6]), .Y(N417) );
  XOR2X1 U1705 ( .A(w0[22]), .B(sa10_sr[6]), .Y(N409) );
  XOR2X1 U1706 ( .A(w3[30]), .B(sa03_sr[6]), .Y(N401) );
  XOR2X1 U1707 ( .A(w2[30]), .B(sa02_sr[6]), .Y(N393) );
  XOR2X1 U1708 ( .A(w1[30]), .B(sa01_sr[6]), .Y(N385) );
  XOR2X1 U1709 ( .A(w0[30]), .B(sa00_sr[6]), .Y(N377) );
  XOR2X1 U1710 ( .A(w2[23]), .B(sa12_sr[7]), .Y(N424) );
  XOR2X1 U1711 ( .A(w1[23]), .B(sa11_sr[7]), .Y(N416) );
  XOR2X1 U1712 ( .A(w0[23]), .B(sa10_sr[7]), .Y(N408) );
  XOR2X1 U1713 ( .A(w3[14]), .B(sa23_sr[6]), .Y(N465) );
  XOR2X1 U1714 ( .A(w2[14]), .B(sa22_sr[6]), .Y(N457) );
  XOR2X1 U1715 ( .A(w1[14]), .B(sa21_sr[6]), .Y(N449) );
  XOR2X1 U1716 ( .A(w0[14]), .B(sa20_sr[6]), .Y(N441) );
  XOR2X1 U1717 ( .A(w2[15]), .B(sa22_sr[7]), .Y(N456) );
  XOR2X1 U1718 ( .A(w1[15]), .B(sa21_sr[7]), .Y(N448) );
  XOR2X1 U1719 ( .A(w0[15]), .B(sa20_sr[7]), .Y(N440) );
  XOR2X1 U1720 ( .A(w2[31]), .B(sa02_sr[7]), .Y(N392) );
  XOR2X1 U1721 ( .A(w1[31]), .B(sa01_sr[7]), .Y(N384) );
  XOR2X1 U1722 ( .A(w0[31]), .B(sa00_sr[7]), .Y(N376) );
  XOR2X1 U1723 ( .A(w3[1]), .B(sa33_sr[1]), .Y(N502) );
  XOR2X1 U1724 ( .A(w3[5]), .B(sa33_sr[5]), .Y(N498) );
  XOR2X1 U1725 ( .A(w3[9]), .B(sa23_sr[1]), .Y(N470) );
  XOR2X1 U1726 ( .A(w3[13]), .B(sa23_sr[5]), .Y(N466) );
  XOR2X1 U1727 ( .A(w3[17]), .B(sa13_sr[1]), .Y(N438) );
  XOR2X1 U1728 ( .A(w3[21]), .B(sa13_sr[5]), .Y(N434) );
  XOR2X1 U1729 ( .A(w3[25]), .B(sa03_sr[1]), .Y(N406) );
  XOR2X1 U1730 ( .A(w3[29]), .B(sa03_sr[5]), .Y(N402) );
  XOR2X1 U1731 ( .A(w2[3]), .B(sa32_sr[3]), .Y(N492) );
  XOR2X1 U1732 ( .A(w1[3]), .B(sa31_sr[3]), .Y(N484) );
  XOR2X1 U1733 ( .A(w0[3]), .B(sa30_sr[3]), .Y(N476) );
  XOR2X1 U1734 ( .A(w2[1]), .B(sa32_sr[1]), .Y(N494) );
  XOR2X1 U1735 ( .A(w1[1]), .B(sa31_sr[1]), .Y(N486) );
  XOR2X1 U1736 ( .A(w0[1]), .B(sa30_sr[1]), .Y(N478) );
  XOR2X1 U1737 ( .A(w2[5]), .B(sa32_sr[5]), .Y(N490) );
  XOR2X1 U1738 ( .A(w1[5]), .B(sa31_sr[5]), .Y(N482) );
  XOR2X1 U1739 ( .A(w0[5]), .B(sa30_sr[5]), .Y(N474) );
  XOR2X1 U1740 ( .A(w2[9]), .B(sa22_sr[1]), .Y(N462) );
  XOR2X1 U1741 ( .A(w2[11]), .B(sa22_sr[3]), .Y(N460) );
  XOR2X1 U1742 ( .A(w2[13]), .B(sa22_sr[5]), .Y(N458) );
  XOR2X1 U1743 ( .A(w1[9]), .B(sa21_sr[1]), .Y(N454) );
  XOR2X1 U1744 ( .A(w1[11]), .B(sa21_sr[3]), .Y(N452) );
  XOR2X1 U1745 ( .A(w1[13]), .B(sa21_sr[5]), .Y(N450) );
  XOR2X1 U1746 ( .A(w0[9]), .B(sa20_sr[1]), .Y(N446) );
  XOR2X1 U1747 ( .A(w0[11]), .B(sa20_sr[3]), .Y(N444) );
  XOR2X1 U1748 ( .A(w0[13]), .B(sa20_sr[5]), .Y(N442) );
  XOR2X1 U1749 ( .A(w2[17]), .B(sa12_sr[1]), .Y(N430) );
  XOR2X1 U1750 ( .A(w2[19]), .B(sa12_sr[3]), .Y(N428) );
  XOR2X1 U1751 ( .A(w2[21]), .B(sa12_sr[5]), .Y(N426) );
  XOR2X1 U1752 ( .A(w1[17]), .B(sa11_sr[1]), .Y(N422) );
  XOR2X1 U1753 ( .A(w1[19]), .B(sa11_sr[3]), .Y(N420) );
  XOR2X1 U1754 ( .A(w1[21]), .B(sa11_sr[5]), .Y(N418) );
  XOR2X1 U1755 ( .A(w0[17]), .B(sa10_sr[1]), .Y(N414) );
  XOR2X1 U1756 ( .A(w0[19]), .B(sa10_sr[3]), .Y(N412) );
  XOR2X1 U1757 ( .A(w0[21]), .B(sa10_sr[5]), .Y(N410) );
  XOR2X1 U1758 ( .A(w2[25]), .B(sa02_sr[1]), .Y(N398) );
  XOR2X1 U1759 ( .A(w2[27]), .B(sa02_sr[3]), .Y(N396) );
  XOR2X1 U1760 ( .A(w2[29]), .B(sa02_sr[5]), .Y(N394) );
  XOR2X1 U1761 ( .A(w1[25]), .B(sa01_sr[1]), .Y(N390) );
  XOR2X1 U1762 ( .A(w1[27]), .B(sa01_sr[3]), .Y(N388) );
  XOR2X1 U1763 ( .A(w1[29]), .B(sa01_sr[5]), .Y(N386) );
  XOR2X1 U1764 ( .A(w0[25]), .B(sa00_sr[1]), .Y(N382) );
  XOR2X1 U1765 ( .A(w0[27]), .B(sa00_sr[3]), .Y(N380) );
  XOR2X1 U1766 ( .A(w0[29]), .B(sa00_sr[5]), .Y(N378) );
  OAI211X1 U1767 ( .A0(dcnt[3]), .A1(n728), .B0(n1012), .C0(rst), .Y(n732) );
  OAI21XL U1768 ( .A0(n734), .A1(n732), .B0(n733), .Y(n146) );
  AOI21X1 U1769 ( .A0(dcnt[1]), .A1(dcnt[0]), .B0(n735), .Y(n734) );
  OAI21XL U1770 ( .A0(dcnt[0]), .A1(n732), .B0(n733), .Y(n147) );
  AOI21X1 U1771 ( .A0(n728), .A1(n736), .B0(n732), .Y(n145) );
  NAND2X1 U1772 ( .A(n866), .B(n729), .Y(n736) );
  OAI31X1 U1773 ( .A0(n727), .A1(n731), .A2(n732), .B0(n733), .Y(n995) );
  INVX1 U1774 ( .A(dcnt[3]), .Y(n727) );
  INVX1 U1775 ( .A(n6), .Y(n1008) );
  NOR3BX1 U1776 ( .AN(dcnt[0]), .B(n811), .C(dcnt[1]), .Y(N21) );
  OR3XL U1777 ( .A(n866), .B(n1009), .C(dcnt[3]), .Y(n811) );
  INVX8 U1778 ( .A(n1013), .Y(n1009) );
  INVX1 U1779 ( .A(ld), .Y(n1013) );
  INVX1 U1780 ( .A(ld), .Y(n1012) );
endmodule

