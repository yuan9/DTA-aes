module aes_rcon ( clk, kld, out );
  output [31:0] out;
  input clk, kld;
  wire   N45, N46, N47, N48, N49, N51, N52, n1, n2, n5, n6, n3, n4, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22;
  wire   [3:0] rcnt;

  DFFX1 \rcnt_reg[0]  ( .D(N52), .CK(clk), .Q(rcnt[0]), .QN(n3) );
  DFFTRX1 \rcnt_reg[2]  ( .D(n4), .RN(n5), .CK(clk), .Q(rcnt[2]) );
  DFFTRX1 \rcnt_reg[3]  ( .D(n4), .RN(n1), .CK(clk), .Q(rcnt[3]) );
  DFFTRX1 \out_reg[30]  ( .D(n6), .RN(n2), .CK(clk), .Q(out[30]) );
  DFFHQX1 \out_reg[31]  ( .D(N51), .CK(clk), .Q(out[31]) );
  DFFHQX1 \out_reg[25]  ( .D(N45), .CK(clk), .Q(out[25]) );
  DFFHQX1 \out_reg[28]  ( .D(N48), .CK(clk), .Q(out[28]) );
  DFFHQX1 \out_reg[29]  ( .D(N49), .CK(clk), .Q(out[29]) );
  DFFHQX1 \out_reg[26]  ( .D(N46), .CK(clk), .Q(out[26]) );
  DFFHQX1 \out_reg[27]  ( .D(N47), .CK(clk), .Q(out[27]) );
  DFFTRX1 \rcnt_reg[1]  ( .D(n4), .RN(n6), .CK(clk), .Q(rcnt[1]) );
  DFFTRXL \out_reg[24]  ( .D(n22), .RN(n4), .CK(clk), .QN(out[24]) );
  INVX1 U3 ( .A(kld), .Y(n4) );
  NOR2XL U4 ( .A(n1), .B(n5), .Y(n18) );
  INVX1 U5 ( .A(n21), .Y(n5) );
  INVX1 U6 ( .A(n10), .Y(n7) );
  NAND4XL U7 ( .A(rcnt[0]), .B(n18), .C(n4), .D(n10), .Y(n11) );
  NAND3XL U8 ( .A(rcnt[1]), .B(n18), .C(N52), .Y(n12) );
  OAI2BB1XL U9 ( .A0N(n2), .A1N(n15), .B0(n14), .Y(N48) );
  AOI211XL U10 ( .A0(n5), .A1(n19), .B0(n18), .C0(n17), .Y(N49) );
  NOR3XL U11 ( .A(n1), .B(n21), .C(n20), .Y(N51) );
  NOR3XL U12 ( .A(n1), .B(n21), .C(n13), .Y(n2) );
  INVXL U13 ( .A(n16), .Y(n19) );
  INVXL U14 ( .A(n6), .Y(n15) );
  NAND2XL U15 ( .A(rcnt[1]), .B(N52), .Y(n20) );
  NAND2XL U16 ( .A(n8), .B(N52), .Y(n17) );
  NAND2XL U17 ( .A(rcnt[0]), .B(n4), .Y(n13) );
  NOR2XL U18 ( .A(rcnt[0]), .B(rcnt[1]), .Y(n8) );
  NAND2X1 U19 ( .A(rcnt[0]), .B(rcnt[1]), .Y(n10) );
  OAI21X1 U20 ( .A0(n7), .A1(rcnt[2]), .B0(n22), .Y(n21) );
  NAND2X1 U21 ( .A(rcnt[2]), .B(n7), .Y(n22) );
  NOR2X1 U22 ( .A(n7), .B(n8), .Y(n6) );
  NOR2X1 U23 ( .A(rcnt[0]), .B(kld), .Y(N52) );
  INVX1 U24 ( .A(n22), .Y(n9) );
  NOR2X1 U25 ( .A(n9), .B(rcnt[3]), .Y(n16) );
  AOI21X1 U26 ( .A0(rcnt[3]), .A1(n9), .B0(n16), .Y(n1) );
  NAND4X1 U27 ( .A(n1), .B(n4), .C(n21), .D(n15), .Y(n14) );
  OAI21XL U28 ( .A0(n5), .A1(n17), .B0(n14), .Y(N45) );
  OAI21XL U29 ( .A0(rcnt[0]), .A1(n14), .B0(n11), .Y(N46) );
  OAI21XL U30 ( .A0(n14), .A1(n3), .B0(n12), .Y(N47) );
endmodule


module aes_sbox_0 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368;

  INVX1 U1 ( .A(n93), .Y(n341) );
  NOR2BX1 U2 ( .AN(n349), .B(n311), .Y(n250) );
  AOI211XL U3 ( .A0(n287), .A1(n286), .B0(n285), .C0(n284), .Y(n288) );
  AOI31XL U4 ( .A0(n263), .A1(n262), .A2(n261), .B0(n341), .Y(n285) );
  AOI211X1 U5 ( .A0(n287), .A1(n222), .B0(n221), .C0(n220), .Y(n223) );
  NAND2XL U6 ( .A(n239), .B(n268), .Y(n339) );
  NOR2XL U7 ( .A(n328), .B(n146), .Y(n358) );
  NOR2X1 U8 ( .A(n199), .B(n273), .Y(n165) );
  INVX1 U9 ( .A(n325), .Y(n268) );
  NOR2X1 U10 ( .A(a[2]), .B(n278), .Y(n70) );
  AOI31XL U11 ( .A0(n29), .A1(n28), .A2(n27), .B0(n341), .Y(n30) );
  AOI31XL U12 ( .A0(n125), .A1(n124), .A2(n123), .B0(n341), .Y(n126) );
  AOI211X1 U13 ( .A0(n1), .A1(n308), .B0(n183), .C0(n182), .Y(n224) );
  AOI211XL U14 ( .A0(n189), .A1(n188), .B0(n187), .C0(n186), .Y(n195) );
  AOI21XL U15 ( .A0(n340), .A1(n339), .B0(n338), .Y(n342) );
  AOI2BB2XL U16 ( .B0(n360), .B1(n291), .A0N(n350), .A1N(n290), .Y(n302) );
  INVXL U17 ( .A(n260), .Y(n291) );
  NOR2XL U18 ( .A(n228), .B(n327), .Y(n260) );
  AOI32XL U19 ( .A0(n113), .A1(a[7]), .A2(n269), .B0(n163), .B1(n267), .Y(n197) );
  NAND2XL U20 ( .A(n113), .B(n82), .Y(n162) );
  INVXL U21 ( .A(n154), .Y(n312) );
  NAND2XL U22 ( .A(n144), .B(n24), .Y(n155) );
  NAND2XL U23 ( .A(a[1]), .B(n295), .Y(n86) );
  NOR2X1 U24 ( .A(a[1]), .B(n295), .Y(n320) );
  NOR2XL U25 ( .A(n325), .B(n135), .Y(n265) );
  NAND2XL U26 ( .A(n198), .B(n277), .Y(n345) );
  NOR2X1 U27 ( .A(n295), .B(n5), .Y(n154) );
  NAND2XL U28 ( .A(n313), .B(n240), .Y(n347) );
  AOI2BB2XL U29 ( .B0(n360), .B1(n164), .A0N(n303), .A1N(n163), .Y(n169) );
  NAND2XL U30 ( .A(n330), .B(n5), .Y(n249) );
  CLKINVX3 U31 ( .A(n328), .Y(n2) );
  INVX1 U32 ( .A(n298), .Y(n355) );
  INVXL U33 ( .A(n270), .Y(n334) );
  CLKINVX3 U34 ( .A(n269), .Y(n330) );
  NOR2XL U35 ( .A(n5), .B(n269), .Y(n191) );
  NOR2X1 U36 ( .A(a[1]), .B(n107), .Y(n332) );
  NOR2XL U37 ( .A(a[1]), .B(n246), .Y(n190) );
  NAND2X1 U38 ( .A(a[1]), .B(n35), .Y(n353) );
  NAND2X1 U39 ( .A(a[6]), .B(a[0]), .Y(n361) );
  INVX1 U40 ( .A(a[3]), .Y(n35) );
  AOI211XL U41 ( .A0(n129), .A1(n128), .B0(n127), .C0(n126), .Y(n130) );
  AOI211XL U42 ( .A0(n129), .A1(n32), .B0(n31), .C0(n30), .Y(n33) );
  AOI211XL U43 ( .A0(n329), .A1(n260), .B0(n259), .C0(n258), .Y(n261) );
  AOI211XL U44 ( .A0(n129), .A1(n62), .B0(n61), .C0(n60), .Y(n63) );
  OAI211XL U45 ( .A0(n249), .A1(n355), .B0(n248), .C0(n247), .Y(n286) );
  AOI211XL U46 ( .A0(n93), .A1(n92), .B0(n91), .C0(n90), .Y(n94) );
  OR4X2 U47 ( .A(n368), .B(n367), .C(n366), .D(n365), .Y(d[0]) );
  AOI31XL U48 ( .A0(n23), .A1(n22), .A2(n21), .B0(n299), .Y(n31) );
  AOI31XL U49 ( .A0(n59), .A1(n58), .A2(n57), .B0(n341), .Y(n60) );
  AOI31XL U50 ( .A0(n246), .A1(n256), .A2(n245), .B0(n244), .Y(n248) );
  OAI22XL U51 ( .A0(n257), .A1(n350), .B0(n256), .B1(n255), .Y(n258) );
  AOI31XL U52 ( .A0(n89), .A1(n88), .A2(n87), .B0(n299), .Y(n90) );
  OAI211XL U53 ( .A0(n74), .A1(n121), .B0(n73), .C0(n72), .Y(n92) );
  AOI31XL U54 ( .A0(n302), .A1(n301), .A2(n300), .B0(n299), .Y(n368) );
  AOI31XL U55 ( .A0(n344), .A1(n343), .A2(n342), .B0(n341), .Y(n366) );
  AOI211XL U56 ( .A0(n260), .A1(n360), .B0(n19), .C0(n18), .Y(n21) );
  AOI31XL U57 ( .A0(n170), .A1(n169), .A2(n168), .B0(n341), .Y(n171) );
  AOI211XL U58 ( .A0(n192), .A1(n4), .B0(n143), .C0(n142), .Y(n175) );
  OAI211XL U59 ( .A0(n197), .A1(n196), .B0(n195), .C0(n194), .Y(n222) );
  AOI22XL U60 ( .A0(n257), .A1(n298), .B0(n268), .B1(n106), .Y(n109) );
  AOI31XL U61 ( .A0(n212), .A1(n211), .A2(n210), .B0(n361), .Y(n221) );
  AOI31XL U62 ( .A0(n161), .A1(n160), .A2(n159), .B0(n321), .Y(n172) );
  AOI211XL U63 ( .A0(n4), .A1(n339), .B0(n358), .C0(n148), .Y(n151) );
  AOI31XL U64 ( .A0(n219), .A1(n218), .A2(n217), .B0(n321), .Y(n220) );
  OAI211XL U65 ( .A0(n350), .A1(n268), .B0(n141), .C0(n140), .Y(n142) );
  AOI211XL U66 ( .A0(n1), .A1(n207), .B0(n206), .C0(n205), .Y(n211) );
  AOI211XL U67 ( .A0(n250), .A1(n240), .B0(n178), .C0(n56), .Y(n57) );
  NAND2XL U68 ( .A(n298), .B(n105), .Y(n98) );
  INVXL U69 ( .A(n105), .Y(n257) );
  AOI211XL U70 ( .A0(n326), .A1(n188), .B0(n52), .C0(n167), .Y(n53) );
  AOI211XL U71 ( .A0(n3), .A1(n86), .B0(n51), .C0(n50), .Y(n54) );
  OAI211XL U72 ( .A0(n337), .A1(n237), .B0(n181), .C0(n180), .Y(n182) );
  AOI31XL U73 ( .A0(n118), .A1(n117), .A2(n247), .B0(n361), .Y(n127) );
  AOI211XL U74 ( .A0(n298), .A1(n105), .B0(n40), .C0(n39), .Y(n64) );
  AOI211XL U75 ( .A0(n329), .A1(n162), .B0(n85), .C0(n84), .Y(n88) );
  AOI31XL U76 ( .A0(n283), .A1(n282), .A2(n281), .B0(n361), .Y(n284) );
  AOI211XL U77 ( .A0(n346), .A1(n268), .B0(n143), .C0(n119), .Y(n125) );
  AOI31XL U78 ( .A0(n81), .A1(n80), .A2(n97), .B0(n321), .Y(n91) );
  AOI211XL U79 ( .A0(n329), .A1(n198), .B0(n71), .C0(n143), .Y(n72) );
  AOI21X1 U80 ( .A0(n360), .A1(n227), .B0(n69), .Y(n95) );
  AOI22XL U81 ( .A0(n2), .A1(n207), .B0(n192), .B1(n122), .Y(n123) );
  AOI31XL U82 ( .A0(n324), .A1(n323), .A2(n322), .B0(n321), .Y(n367) );
  AOI211XL U83 ( .A0(n2), .A1(n291), .B0(n167), .C0(n166), .Y(n168) );
  AOI31XL U84 ( .A0(n364), .A1(n363), .A2(n362), .B0(n361), .Y(n365) );
  AOI211XL U85 ( .A0(a[7]), .A1(n339), .B0(n96), .C0(n115), .Y(n19) );
  AOI211XL U86 ( .A0(n350), .A1(n303), .B0(n185), .C0(n264), .Y(n186) );
  AOI211XL U87 ( .A0(n329), .A1(n266), .B0(n216), .C0(n215), .Y(n218) );
  AOI211XL U88 ( .A0(n298), .A1(n179), .B0(n178), .C0(n177), .Y(n181) );
  AOI211XL U89 ( .A0(n320), .A1(n1), .B0(n319), .C0(n318), .Y(n322) );
  AOI211XL U90 ( .A0(n360), .A1(n359), .B0(n358), .C0(n357), .Y(n362) );
  AOI22XL U91 ( .A0(n2), .A1(n227), .B0(n3), .B1(n226), .Y(n234) );
  AOI211XL U92 ( .A0(n4), .A1(n251), .B0(n250), .C0(n314), .Y(n263) );
  AOI2BB2XL U93 ( .B0(n264), .B1(n360), .A0N(n350), .A1N(n265), .Y(n283) );
  OAI211XL U94 ( .A0(n252), .A1(n336), .B0(n68), .C0(n67), .Y(n69) );
  AOI221XL U95 ( .A0(n346), .A1(n330), .B0(n3), .B1(n269), .C0(n116), .Y(n117)
         );
  NAND2XL U96 ( .A(n239), .B(n277), .Y(n188) );
  AOI2BB2XL U97 ( .B0(n4), .B1(n337), .A0N(n350), .A1N(n179), .Y(n48) );
  AOI211XL U98 ( .A0(n298), .A1(n290), .B0(n79), .C0(n78), .Y(n80) );
  AOI211XL U99 ( .A0(n2), .A1(n139), .B0(n138), .C0(n137), .Y(n140) );
  AOI211XL U100 ( .A0(a[2]), .A1(n134), .B0(n317), .C0(n133), .Y(n138) );
  AOI22XL U101 ( .A0(n1), .A1(n24), .B0(n346), .B1(n320), .Y(n9) );
  AOI2BB2XL U102 ( .B0(n4), .B1(n86), .A0N(n237), .A1N(n104), .Y(n55) );
  NOR2XL U103 ( .A(n228), .B(n154), .Y(n120) );
  NOR2XL U104 ( .A(n185), .B(n99), .Y(n178) );
  AOI22XL U105 ( .A0(n4), .A1(n162), .B0(n329), .B1(n179), .Y(n170) );
  AOI22XL U106 ( .A0(n1), .A1(n214), .B0(n329), .B1(n268), .Y(n58) );
  AOI22XL U107 ( .A0(n1), .A1(n290), .B0(n346), .B1(n269), .Y(n157) );
  AOI22XL U108 ( .A0(n3), .A1(n134), .B0(n360), .B1(n266), .Y(n13) );
  AOI22XL U109 ( .A0(n3), .A1(n192), .B0(n360), .B1(n154), .Y(n161) );
  NAND2XL U110 ( .A(n268), .B(n349), .Y(n251) );
  INVXL U111 ( .A(n156), .Y(n226) );
  AOI22XL U112 ( .A0(n1), .A1(n104), .B0(n326), .B1(n176), .Y(n38) );
  OAI22XL U113 ( .A0(n35), .A1(n328), .B0(n201), .B1(n155), .Y(n40) );
  AOI22XL U114 ( .A0(n330), .A1(n3), .B0(n298), .B1(n139), .Y(n68) );
  AOI22XL U115 ( .A0(n1), .A1(n307), .B0(n4), .B1(n42), .Y(n29) );
  AOI22XL U116 ( .A0(n1), .A1(n293), .B0(n259), .B1(n268), .Y(n83) );
  AOI22XL U117 ( .A0(n96), .A1(n1), .B0(n4), .B1(n305), .Y(n81) );
  AOI22XL U118 ( .A0(n165), .A1(n2), .B0(n17), .B1(n268), .Y(n22) );
  AOI2BB2XL U119 ( .B0(n4), .B1(n104), .A0N(n196), .A1N(n103), .Y(n110) );
  AOI22XL U120 ( .A0(n3), .A1(n44), .B0(n346), .B1(n290), .Y(n45) );
  AOI22XL U121 ( .A0(n228), .A1(n329), .B0(n298), .B1(n103), .Y(n47) );
  AOI22XL U122 ( .A0(n1), .A1(n295), .B0(n298), .B1(n327), .Y(n15) );
  AOI211XL U123 ( .A0(n298), .A1(n352), .B0(n297), .C0(n296), .Y(n300) );
  AOI2BB2XL U124 ( .B0(n2), .B1(n293), .A0N(n316), .A1N(n292), .Y(n301) );
  OAI22XL U125 ( .A0(n356), .A1(n354), .B0(n176), .B1(n184), .Y(n177) );
  AOI31XL U126 ( .A0(n2), .A1(n353), .A2(n352), .B0(n310), .Y(n323) );
  AOI22XL U127 ( .A0(n192), .A1(n276), .B0(n237), .B1(n316), .Y(n193) );
  AOI22XL U128 ( .A0(a[3]), .A1(n4), .B0(n1), .B1(n349), .Y(n363) );
  NOR3XL U129 ( .A(n325), .B(n252), .C(n328), .Y(n253) );
  AOI22XL U130 ( .A0(n1), .A1(n230), .B0(n252), .B1(n329), .Y(n233) );
  AOI22XL U131 ( .A0(a[1]), .A1(n4), .B0(n1), .B1(n334), .Y(n219) );
  AOI22XL U132 ( .A0(n2), .A1(n96), .B0(n346), .B1(n5), .Y(n49) );
  NOR2XL U133 ( .A(n295), .B(n294), .Y(n296) );
  INVXL U134 ( .A(n314), .Y(n315) );
  AOI22XL U135 ( .A0(n298), .A1(n154), .B0(n4), .B1(n265), .Y(n8) );
  AOI22XL U136 ( .A0(n2), .A1(n43), .B0(n360), .B1(n42), .Y(n46) );
  AOI22XL U137 ( .A0(n3), .A1(n43), .B0(n346), .B1(n65), .Y(n23) );
  NOR2XL U138 ( .A(n165), .B(n311), .Y(n166) );
  NAND2XL U139 ( .A(n2), .B(n269), .Y(n99) );
  OAI22XL U140 ( .A0(n165), .A1(n303), .B0(n96), .B1(n237), .Y(n102) );
  NOR2XL U141 ( .A(n154), .B(n332), .Y(n134) );
  AOI22XL U142 ( .A0(n271), .A1(n4), .B0(n2), .B1(n155), .Y(n160) );
  AOI22XL U143 ( .A0(n298), .A1(n146), .B0(n4), .B1(n163), .Y(n89) );
  OAI211XL U144 ( .A0(n277), .A1(n276), .B0(n275), .C0(n274), .Y(n279) );
  OAI2BB1XL U145 ( .A0N(n214), .A1N(n326), .B0(n247), .Y(n215) );
  AOI22XL U146 ( .A0(n70), .A1(n154), .B0(n4), .B1(n266), .Y(n73) );
  AOI22XL U147 ( .A0(n2), .A1(n121), .B0(n329), .B1(n155), .Y(n28) );
  INVXL U148 ( .A(n184), .Y(n187) );
  AOI211XL U149 ( .A0(n2), .A1(n271), .B0(n66), .C0(n297), .Y(n67) );
  AOI22XL U150 ( .A0(n3), .A1(n230), .B0(n4), .B1(n225), .Y(n203) );
  NAND2XL U151 ( .A(n113), .B(n246), .Y(n139) );
  AOI22XL U152 ( .A0(n199), .A1(n333), .B0(n329), .B1(n345), .Y(n212) );
  INVXL U153 ( .A(n86), .Y(n176) );
  AOI22XL U154 ( .A0(n330), .A1(n329), .B0(n2), .B1(n327), .Y(n343) );
  AOI22XL U155 ( .A0(n3), .A1(n347), .B0(n346), .B1(n345), .Y(n364) );
  NAND2XL U156 ( .A(n353), .B(n352), .Y(n359) );
  NAND3XL U157 ( .A(n3), .B(n144), .C(n86), .Y(n87) );
  NOR2XL U158 ( .A(n213), .B(n237), .Y(n259) );
  AOI22XL U159 ( .A0(n2), .A1(n292), .B0(n334), .B1(n4), .Y(n241) );
  AOI22XL U160 ( .A0(n189), .A1(n320), .B0(n2), .B1(n265), .Y(n114) );
  NAND2XL U161 ( .A(n107), .B(n256), .Y(n307) );
  AOI22XL U162 ( .A0(n3), .A1(n266), .B0(n329), .B1(n265), .Y(n282) );
  AOI22XL U163 ( .A0(a[3]), .A1(n346), .B0(n2), .B1(n202), .Y(n204) );
  AOI22XL U164 ( .A0(n185), .A1(n4), .B0(n329), .B1(n272), .Y(n100) );
  AOI22XL U165 ( .A0(n271), .A1(n360), .B0(n340), .B1(n332), .Y(n147) );
  AOI22XL U166 ( .A0(a[1]), .A1(n298), .B0(n3), .B1(n144), .Y(n153) );
  INVXL U167 ( .A(n135), .Y(n352) );
  NOR2XL U168 ( .A(n185), .B(n272), .Y(n317) );
  AOI22XL U169 ( .A0(n298), .A1(n132), .B0(n360), .B1(n308), .Y(n141) );
  OAI22XL U170 ( .A0(n327), .A1(n237), .B0(n201), .B1(n200), .Y(n206) );
  NAND2XL U171 ( .A(n4), .B(n249), .Y(n184) );
  NAND2XL U172 ( .A(n313), .B(n200), .Y(n44) );
  NOR2XL U173 ( .A(n41), .B(n149), .Y(n103) );
  AOI22XL U174 ( .A0(n190), .A1(n360), .B0(n329), .B1(n107), .Y(n37) );
  AOI22XL U175 ( .A0(n230), .A1(n209), .B0(n360), .B1(n313), .Y(n10) );
  AND2X2 U176 ( .A(n305), .B(n82), .Y(n225) );
  NOR2XL U177 ( .A(n295), .B(n230), .Y(n43) );
  AOI31XL U178 ( .A0(n355), .A1(n237), .A2(n180), .B0(n330), .Y(n71) );
  NOR2XL U179 ( .A(n271), .B(n355), .Y(n17) );
  NOR3XL U180 ( .A(n185), .B(n264), .C(n311), .Y(n297) );
  AOI211XL U181 ( .A0(a[7]), .A1(n65), .B0(n191), .C0(n115), .Y(n66) );
  AOI22XL U182 ( .A0(n230), .A1(n4), .B0(n340), .B1(n356), .Y(n124) );
  OAI22XL U183 ( .A0(n355), .A1(n198), .B0(n308), .B1(n316), .Y(n119) );
  AOI22XL U184 ( .A0(n4), .A1(n353), .B0(n112), .B1(n111), .Y(n118) );
  AOI22XL U185 ( .A0(a[4]), .A1(n298), .B0(n346), .B1(n308), .Y(n25) );
  AOI22XL U186 ( .A0(n271), .A1(n326), .B0(n331), .B1(n270), .Y(n275) );
  NOR2XL U187 ( .A(n191), .B(n190), .Y(n292) );
  NAND2XL U188 ( .A(n111), .B(n349), .Y(n179) );
  AOI22XL U189 ( .A0(n334), .A1(n333), .B0(n332), .B1(n331), .Y(n335) );
  AOI22XL U190 ( .A0(n326), .A1(n325), .B0(n3), .B1(n5), .Y(n344) );
  NAND3XL U191 ( .A(n3), .B(a[3]), .C(n208), .Y(n77) );
  OR2X2 U192 ( .A(a[7]), .B(n115), .Y(n350) );
  NAND2XL U193 ( .A(n313), .B(n305), .Y(n42) );
  AOI22XL U194 ( .A0(n145), .A1(n333), .B0(n254), .B1(n331), .Y(n152) );
  NOR2XL U195 ( .A(n237), .B(n332), .Y(n112) );
  NOR2XL U196 ( .A(a[1]), .B(n330), .Y(n272) );
  NOR2XL U197 ( .A(a[1]), .B(n252), .Y(n135) );
  AOI22XL U198 ( .A0(n191), .A1(n209), .B0(n329), .B1(n309), .Y(n16) );
  NAND2XL U199 ( .A(n308), .B(n270), .Y(n65) );
  NOR2XL U200 ( .A(n41), .B(a[1]), .Y(n199) );
  NAND3XL U201 ( .A(n209), .B(n246), .C(n208), .Y(n210) );
  INVXL U202 ( .A(n299), .Y(n287) );
  INVXL U203 ( .A(n333), .Y(n238) );
  INVXL U204 ( .A(n201), .Y(n189) );
  NAND2XL U205 ( .A(n329), .B(n313), .Y(n354) );
  NAND3XL U206 ( .A(n333), .B(n76), .C(n246), .Y(n75) );
  NAND2XL U207 ( .A(a[1]), .B(n264), .Y(n305) );
  INVXL U208 ( .A(n196), .Y(n209) );
  OR2X2 U209 ( .A(n267), .B(n196), .Y(n328) );
  NAND2XL U210 ( .A(a[2]), .B(n278), .Y(n196) );
  NOR2XL U211 ( .A(a[1]), .B(n202), .Y(n164) );
  NAND2XL U212 ( .A(n267), .B(n278), .Y(n255) );
  NOR2XL U213 ( .A(n267), .B(n276), .Y(n331) );
  INVXL U214 ( .A(n277), .Y(n254) );
  AOI22XL U215 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n276), .Y(n136) );
  AOI22XL U216 ( .A0(a[1]), .A1(a[7]), .B0(n267), .B1(n5), .Y(n76) );
  INVX2 U217 ( .A(a[4]), .Y(n202) );
  INVX2 U218 ( .A(a[5]), .Y(n278) );
  INVX2 U219 ( .A(a[2]), .Y(n276) );
  NAND2XL U220 ( .A(a[3]), .B(a[1]), .Y(n24) );
  NOR2XL U221 ( .A(a[3]), .B(a[1]), .Y(n229) );
  NAND2XL U222 ( .A(a[4]), .B(a[1]), .Y(n277) );
  NAND2X2 U223 ( .A(n278), .B(n276), .Y(n201) );
  NOR2X2 U224 ( .A(n35), .B(n202), .Y(n264) );
  NOR2X2 U225 ( .A(n41), .B(n5), .Y(n185) );
  NAND2X2 U226 ( .A(a[1]), .B(n246), .Y(n308) );
  NAND2X2 U227 ( .A(a[3]), .B(n202), .Y(n246) );
  NOR2X2 U228 ( .A(n276), .B(a[7]), .Y(n326) );
  NOR2X2 U229 ( .A(n252), .B(n330), .Y(n295) );
  NOR2X2 U230 ( .A(n330), .B(n5), .Y(n230) );
  NAND2X2 U231 ( .A(n202), .B(n5), .Y(n313) );
  CLKINVX3 U232 ( .A(n237), .Y(n360) );
  NAND2X2 U233 ( .A(a[5]), .B(n326), .Y(n237) );
  CLKINVX3 U234 ( .A(n350), .Y(n1) );
  NOR2X4 U235 ( .A(a[2]), .B(n133), .Y(n329) );
  BUFX3 U236 ( .A(n348), .Y(n3) );
  NOR2X4 U237 ( .A(a[7]), .B(n201), .Y(n298) );
  CLKINVX3 U238 ( .A(a[1]), .Y(n5) );
  CLKINVX3 U239 ( .A(n311), .Y(n346) );
  NAND2X2 U240 ( .A(n278), .B(n326), .Y(n311) );
  BUFX3 U241 ( .A(n351), .Y(n4) );
  AOI21XL U242 ( .A0(n313), .A1(n312), .B0(n311), .Y(n319) );
  AOI21XL U243 ( .A0(n309), .A1(n308), .B0(n336), .Y(n310) );
  AOI21XL U244 ( .A0(n360), .A1(n307), .B0(n306), .Y(n324) );
  AOI21XL U245 ( .A0(n305), .A1(n304), .B0(n303), .Y(n306) );
  AOI21XL U246 ( .A0(n4), .A1(n308), .B0(n3), .Y(n294) );
  AOI21XL U247 ( .A0(n213), .A1(n308), .B0(n328), .Y(n216) );
  AOI21XL U248 ( .A0(n270), .A1(n353), .B0(n311), .Y(n183) );
  AOI21XL U249 ( .A0(n329), .A1(n226), .B0(n158), .Y(n159) );
  AOI21XL U250 ( .A0(n136), .A1(n352), .B0(n311), .Y(n137) );
  AOI21XL U251 ( .A0(n240), .A1(n249), .B0(n328), .Y(n85) );
  AOI21XL U252 ( .A0(n209), .A1(n320), .B0(n346), .Y(n74) );
  AOI21XL U253 ( .A0(n54), .A1(n53), .B0(n361), .Y(n61) );
  AOI21XL U254 ( .A0(n240), .A1(n82), .B0(n316), .Y(n51) );
  AOI21XL U255 ( .A0(n360), .A1(n290), .B0(n26), .Y(n27) );
  AOI21XL U256 ( .A0(n146), .A1(n353), .B0(n336), .Y(n18) );
  AOI21XL U257 ( .A0(n2), .A1(n251), .B0(n52), .Y(n14) );
  AOI21XL U258 ( .A0(n313), .A1(n200), .B0(n336), .Y(n52) );
  AOI21XL U259 ( .A0(n269), .A1(n268), .B0(n267), .Y(n280) );
  AOI21XL U260 ( .A0(n254), .A1(n3), .B0(n253), .Y(n262) );
  AOI21XL U261 ( .A0(n346), .A1(n347), .B0(n242), .Y(n243) );
  NOR2X1 U262 ( .A(n276), .B(n133), .Y(n348) );
  NOR2X1 U263 ( .A(n267), .B(n201), .Y(n351) );
  INVX1 U264 ( .A(a[7]), .Y(n267) );
  OAI21XL U265 ( .A0(n224), .A1(n341), .B0(n223), .Y(d[2]) );
  OAI21XL U266 ( .A0(n175), .A1(n361), .B0(n174), .Y(d[3]) );
  OAI21XL U267 ( .A0(n95), .A1(n361), .B0(n94), .Y(d[5]) );
  OAI21XL U268 ( .A0(n64), .A1(n299), .B0(n63), .Y(d[6]) );
  OAI21XL U269 ( .A0(n34), .A1(n361), .B0(n33), .Y(d[7]) );
  OAI21XL U270 ( .A0(n131), .A1(n299), .B0(n130), .Y(d[4]) );
  OAI21XL U271 ( .A0(n289), .A1(n321), .B0(n288), .Y(d[1]) );
  NAND2X1 U272 ( .A(a[7]), .B(a[5]), .Y(n133) );
  NOR2X1 U273 ( .A(n5), .B(n246), .Y(n214) );
  NAND2X1 U274 ( .A(a[4]), .B(n35), .Y(n269) );
  NOR2X1 U275 ( .A(a[4]), .B(n5), .Y(n273) );
  OAI21XL U276 ( .A0(n273), .A1(n229), .B0(n3), .Y(n7) );
  NOR2X1 U277 ( .A(a[7]), .B(a[2]), .Y(n340) );
  INVX1 U278 ( .A(n246), .Y(n252) );
  OAI21XL U279 ( .A0(n70), .A1(n340), .B0(n135), .Y(n6) );
  NAND3X1 U280 ( .A(n99), .B(n7), .C(n6), .Y(n12) );
  INVX1 U281 ( .A(n70), .Y(n115) );
  NOR2X1 U282 ( .A(n264), .B(n5), .Y(n325) );
  NAND3X1 U283 ( .A(n10), .B(n9), .C(n8), .Y(n11) );
  AOI211X1 U284 ( .A0(n329), .A1(n214), .B0(n12), .C0(n11), .Y(n34) );
  INVX1 U285 ( .A(a[6]), .Y(n20) );
  NOR2X1 U286 ( .A(a[0]), .B(n20), .Y(n129) );
  INVX1 U287 ( .A(n264), .Y(n309) );
  INVX1 U288 ( .A(n24), .Y(n327) );
  NAND2X1 U289 ( .A(n264), .B(n5), .Y(n349) );
  INVX1 U290 ( .A(n191), .Y(n200) );
  INVX1 U291 ( .A(n4), .Y(n336) );
  NAND2X1 U292 ( .A(n35), .B(n202), .Y(n107) );
  NAND2X1 U293 ( .A(n24), .B(n249), .Y(n266) );
  NAND4X1 U294 ( .A(n16), .B(n15), .C(n14), .D(n13), .Y(n32) );
  NAND2X1 U295 ( .A(a[3]), .B(n5), .Y(n270) );
  INVX1 U296 ( .A(n107), .Y(n41) );
  INVX1 U297 ( .A(n313), .Y(n271) );
  INVX1 U298 ( .A(n295), .Y(n213) );
  NOR2X1 U299 ( .A(a[1]), .B(n213), .Y(n228) );
  INVX1 U300 ( .A(n228), .Y(n239) );
  NAND2X1 U301 ( .A(n5), .B(n309), .Y(n144) );
  NOR2BX1 U302 ( .AN(n144), .B(n185), .Y(n96) );
  INVX1 U303 ( .A(n199), .Y(n146) );
  NAND2X1 U304 ( .A(a[0]), .B(n20), .Y(n299) );
  INVX1 U305 ( .A(n230), .Y(n256) );
  NAND2X1 U306 ( .A(n200), .B(n349), .Y(n121) );
  NAND2X1 U307 ( .A(n309), .B(n86), .Y(n290) );
  INVX1 U308 ( .A(n3), .Y(n303) );
  NAND2X1 U309 ( .A(n239), .B(n353), .Y(n105) );
  OAI21XL U310 ( .A0(n303), .A1(n105), .B0(n25), .Y(n26) );
  NOR2X1 U311 ( .A(a[6]), .B(a[0]), .Y(n93) );
  INVX1 U312 ( .A(n185), .Y(n113) );
  INVX1 U313 ( .A(n229), .Y(n304) );
  NAND2X1 U314 ( .A(n113), .B(n304), .Y(n104) );
  OAI21XL U315 ( .A0(n273), .A1(n164), .B0(n3), .Y(n36) );
  NAND4BXL U316 ( .AN(n250), .B(n38), .C(n37), .D(n36), .Y(n39) );
  INVX1 U317 ( .A(n353), .Y(n145) );
  NOR2X1 U318 ( .A(n145), .B(n332), .Y(n337) );
  INVX1 U319 ( .A(n273), .Y(n111) );
  INVX1 U320 ( .A(n308), .Y(n149) );
  NAND4X1 U321 ( .A(n48), .B(n47), .C(n46), .D(n45), .Y(n62) );
  INVX1 U322 ( .A(n214), .Y(n240) );
  INVX1 U323 ( .A(n332), .Y(n82) );
  INVX1 U324 ( .A(n329), .Y(n316) );
  OAI21XL U325 ( .A0(a[4]), .A1(n350), .B0(n49), .Y(n50) );
  NAND2X1 U326 ( .A(n313), .B(n256), .Y(n293) );
  NOR2X1 U327 ( .A(n355), .B(n293), .Y(n167) );
  OAI21XL U328 ( .A0(n325), .A1(n229), .B0(n298), .Y(n59) );
  OAI21XL U329 ( .A0(n120), .A1(n303), .B0(n55), .Y(n56) );
  NAND2X1 U330 ( .A(n270), .B(n312), .Y(n227) );
  INVX1 U331 ( .A(n190), .Y(n198) );
  NAND2X1 U332 ( .A(n3), .B(n313), .Y(n180) );
  NOR2X1 U333 ( .A(n350), .B(n313), .Y(n143) );
  NOR2X1 U334 ( .A(n278), .B(n276), .Y(n333) );
  OAI21XL U335 ( .A0(n353), .A1(n328), .B0(n75), .Y(n79) );
  INVX1 U336 ( .A(n76), .Y(n208) );
  OAI21XL U337 ( .A0(n225), .A1(n316), .B0(n77), .Y(n78) );
  NAND2X1 U338 ( .A(n346), .B(n213), .Y(n97) );
  INVX1 U339 ( .A(n129), .Y(n321) );
  NAND2X1 U340 ( .A(n111), .B(n270), .Y(n163) );
  OAI21XL U341 ( .A0(n120), .A1(n311), .B0(n83), .Y(n84) );
  NOR2X1 U342 ( .A(n149), .B(n320), .Y(n156) );
  NAND4X1 U343 ( .A(n100), .B(n99), .C(n98), .D(n97), .Y(n101) );
  AOI211X1 U344 ( .A0(n1), .A1(n156), .B0(n102), .C0(n101), .Y(n131) );
  OAI21XL U345 ( .A0(n252), .A1(n350), .B0(n180), .Y(n106) );
  NOR2X1 U346 ( .A(n107), .B(n5), .Y(n356) );
  OAI21XL U347 ( .A0(n190), .A1(n356), .B0(n329), .Y(n108) );
  NAND4BXL U348 ( .AN(n112), .B(n110), .C(n109), .D(n108), .Y(n128) );
  OAI21XL U349 ( .A0(n115), .A1(n197), .B0(n114), .Y(n116) );
  NAND2X1 U350 ( .A(n298), .B(n230), .Y(n247) );
  INVX1 U351 ( .A(n120), .Y(n207) );
  INVX1 U352 ( .A(n121), .Y(n192) );
  OAI21XL U353 ( .A0(n198), .A1(n238), .B0(n237), .Y(n122) );
  OAI21XL U354 ( .A0(a[1]), .A1(n136), .B0(n308), .Y(n132) );
  OAI21XL U355 ( .A0(n311), .A1(n304), .B0(n147), .Y(n148) );
  OAI21XL U356 ( .A0(n330), .A1(n149), .B0(n329), .Y(n150) );
  NAND4X1 U357 ( .A(n153), .B(n152), .C(n151), .D(n150), .Y(n173) );
  OAI21XL U358 ( .A0(n213), .A1(n255), .B0(n157), .Y(n158) );
  AOI211X1 U359 ( .A0(n287), .A1(n173), .B0(n172), .C0(n171), .Y(n174) );
  OAI21XL U360 ( .A0(n292), .A1(n276), .B0(n193), .Y(n194) );
  OAI21XL U361 ( .A0(n204), .A1(n208), .B0(n203), .Y(n205) );
  OAI21XL U362 ( .A0(n320), .A1(n356), .B0(n3), .Y(n217) );
  NOR2X1 U363 ( .A(n225), .B(n336), .Y(n236) );
  OAI21XL U364 ( .A0(n228), .A1(n273), .B0(n346), .Y(n232) );
  OAI21XL U365 ( .A0(n230), .A1(n229), .B0(n360), .Y(n231) );
  NAND4X1 U366 ( .A(n234), .B(n233), .C(n232), .D(n231), .Y(n235) );
  AOI211X1 U367 ( .A0(n337), .A1(n298), .B0(n236), .C0(n235), .Y(n289) );
  OAI21XL U368 ( .A0(n239), .A1(n238), .B0(n237), .Y(n245) );
  OAI21XL U369 ( .A0(n330), .A1(n316), .B0(n241), .Y(n242) );
  OAI21XL U370 ( .A0(n350), .A1(n347), .B0(n243), .Y(n244) );
  NOR2X1 U371 ( .A(n355), .B(n304), .Y(n314) );
  OAI21XL U372 ( .A0(n273), .A1(n272), .B0(n340), .Y(n274) );
  OAI21XL U373 ( .A0(n280), .A1(n279), .B0(n278), .Y(n281) );
  OAI21XL U374 ( .A0(n317), .A1(n316), .B0(n315), .Y(n318) );
  OAI21XL U375 ( .A0(n337), .A1(n336), .B0(n335), .Y(n338) );
  OAI21XL U376 ( .A0(n356), .A1(n355), .B0(n354), .Y(n357) );
endmodule


module aes_sbox_1 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368;

  INVX1 U1 ( .A(n93), .Y(n341) );
  NOR2BX1 U2 ( .AN(n349), .B(n311), .Y(n250) );
  AOI211XL U3 ( .A0(n287), .A1(n286), .B0(n285), .C0(n284), .Y(n288) );
  AOI31XL U4 ( .A0(n263), .A1(n262), .A2(n261), .B0(n341), .Y(n285) );
  AOI211X1 U5 ( .A0(n287), .A1(n222), .B0(n221), .C0(n220), .Y(n223) );
  NAND2XL U6 ( .A(n239), .B(n268), .Y(n339) );
  INVX1 U7 ( .A(n325), .Y(n268) );
  NOR2X1 U8 ( .A(a[2]), .B(n278), .Y(n70) );
  CLKINVX3 U9 ( .A(a[5]), .Y(n278) );
  AOI31XL U10 ( .A0(n29), .A1(n28), .A2(n27), .B0(n341), .Y(n30) );
  AOI211X1 U11 ( .A0(n1), .A1(n308), .B0(n183), .C0(n182), .Y(n224) );
  AOI31XL U12 ( .A0(n125), .A1(n124), .A2(n123), .B0(n341), .Y(n126) );
  AOI21XL U13 ( .A0(n340), .A1(n339), .B0(n338), .Y(n342) );
  AOI2BB2XL U14 ( .B0(n360), .B1(n291), .A0N(n350), .A1N(n290), .Y(n302) );
  AOI211XL U15 ( .A0(n189), .A1(n188), .B0(n187), .C0(n186), .Y(n195) );
  INVXL U16 ( .A(n260), .Y(n291) );
  NOR2XL U17 ( .A(n228), .B(n327), .Y(n260) );
  AOI32XL U18 ( .A0(n113), .A1(a[7]), .A2(n269), .B0(n163), .B1(n267), .Y(n197) );
  INVXL U19 ( .A(n154), .Y(n312) );
  NAND2XL U20 ( .A(n113), .B(n82), .Y(n162) );
  NAND2XL U21 ( .A(a[1]), .B(n295), .Y(n86) );
  NAND2XL U22 ( .A(n313), .B(n240), .Y(n347) );
  AOI2BB2XL U23 ( .B0(n360), .B1(n164), .A0N(n303), .A1N(n163), .Y(n169) );
  NOR2X1 U24 ( .A(n295), .B(n5), .Y(n154) );
  NAND2XL U25 ( .A(n144), .B(n24), .Y(n155) );
  NOR2X1 U26 ( .A(a[1]), .B(n295), .Y(n320) );
  NOR2XL U27 ( .A(n325), .B(n135), .Y(n265) );
  NAND2XL U28 ( .A(n198), .B(n277), .Y(n345) );
  INVX1 U29 ( .A(n298), .Y(n355) );
  NAND2XL U30 ( .A(n330), .B(n5), .Y(n249) );
  CLKINVX3 U31 ( .A(n328), .Y(n2) );
  NOR2X1 U32 ( .A(a[1]), .B(n107), .Y(n332) );
  NOR2XL U33 ( .A(n5), .B(n269), .Y(n191) );
  CLKINVX3 U34 ( .A(n269), .Y(n330) );
  NOR2XL U35 ( .A(a[1]), .B(n246), .Y(n190) );
  INVXL U36 ( .A(n270), .Y(n334) );
  NAND2X1 U37 ( .A(a[1]), .B(n35), .Y(n353) );
  NAND2X1 U38 ( .A(a[6]), .B(a[0]), .Y(n361) );
  INVX1 U39 ( .A(a[3]), .Y(n35) );
  AOI211XL U40 ( .A0(n129), .A1(n128), .B0(n127), .C0(n126), .Y(n130) );
  AOI211XL U41 ( .A0(n129), .A1(n32), .B0(n31), .C0(n30), .Y(n33) );
  AOI31XL U42 ( .A0(n23), .A1(n22), .A2(n21), .B0(n299), .Y(n31) );
  AOI211XL U43 ( .A0(n129), .A1(n62), .B0(n61), .C0(n60), .Y(n63) );
  OAI211XL U44 ( .A0(n249), .A1(n355), .B0(n248), .C0(n247), .Y(n286) );
  AOI211XL U45 ( .A0(n329), .A1(n260), .B0(n259), .C0(n258), .Y(n261) );
  AOI211XL U46 ( .A0(n93), .A1(n92), .B0(n91), .C0(n90), .Y(n94) );
  OR4X2 U47 ( .A(n368), .B(n367), .C(n366), .D(n365), .Y(d[0]) );
  AOI31XL U48 ( .A0(n161), .A1(n160), .A2(n159), .B0(n321), .Y(n172) );
  AOI211XL U49 ( .A0(n260), .A1(n360), .B0(n19), .C0(n18), .Y(n21) );
  AOI31XL U50 ( .A0(n170), .A1(n169), .A2(n168), .B0(n341), .Y(n171) );
  AOI22XL U51 ( .A0(n257), .A1(n298), .B0(n268), .B1(n106), .Y(n109) );
  AOI31XL U52 ( .A0(n302), .A1(n301), .A2(n300), .B0(n299), .Y(n368) );
  AOI31XL U53 ( .A0(n344), .A1(n343), .A2(n342), .B0(n341), .Y(n366) );
  AOI31XL U54 ( .A0(n246), .A1(n256), .A2(n245), .B0(n244), .Y(n248) );
  OAI22XL U55 ( .A0(n257), .A1(n350), .B0(n256), .B1(n255), .Y(n258) );
  OAI211XL U56 ( .A0(n197), .A1(n196), .B0(n195), .C0(n194), .Y(n222) );
  AOI31XL U57 ( .A0(n212), .A1(n211), .A2(n210), .B0(n361), .Y(n221) );
  AOI211XL U58 ( .A0(n192), .A1(n4), .B0(n143), .C0(n142), .Y(n175) );
  AOI31XL U59 ( .A0(n89), .A1(n88), .A2(n87), .B0(n299), .Y(n90) );
  OAI211XL U60 ( .A0(n74), .A1(n121), .B0(n73), .C0(n72), .Y(n92) );
  AOI31XL U61 ( .A0(n59), .A1(n58), .A2(n57), .B0(n341), .Y(n60) );
  AOI211XL U62 ( .A0(n298), .A1(n105), .B0(n40), .C0(n39), .Y(n64) );
  AOI31XL U63 ( .A0(n219), .A1(n218), .A2(n217), .B0(n321), .Y(n220) );
  AOI211XL U64 ( .A0(n1), .A1(n207), .B0(n206), .C0(n205), .Y(n211) );
  AOI211XL U65 ( .A0(n3), .A1(n86), .B0(n51), .C0(n50), .Y(n54) );
  AOI211XL U66 ( .A0(n326), .A1(n188), .B0(n52), .C0(n167), .Y(n53) );
  OAI211XL U67 ( .A0(n337), .A1(n237), .B0(n181), .C0(n180), .Y(n182) );
  AOI211XL U68 ( .A0(n250), .A1(n240), .B0(n178), .C0(n56), .Y(n57) );
  AOI31XL U69 ( .A0(n283), .A1(n282), .A2(n281), .B0(n361), .Y(n284) );
  AOI211XL U70 ( .A0(a[7]), .A1(n339), .B0(n96), .C0(n115), .Y(n19) );
  AOI211XL U71 ( .A0(n2), .A1(n291), .B0(n167), .C0(n166), .Y(n168) );
  NAND2XL U72 ( .A(n298), .B(n105), .Y(n98) );
  INVXL U73 ( .A(n105), .Y(n257) );
  AOI31XL U74 ( .A0(n118), .A1(n117), .A2(n247), .B0(n361), .Y(n127) );
  AOI211XL U75 ( .A0(n346), .A1(n268), .B0(n143), .C0(n119), .Y(n125) );
  AOI22XL U76 ( .A0(n2), .A1(n207), .B0(n192), .B1(n122), .Y(n123) );
  AOI211XL U77 ( .A0(n4), .A1(n339), .B0(n358), .C0(n148), .Y(n151) );
  AOI21X1 U78 ( .A0(n360), .A1(n227), .B0(n69), .Y(n95) );
  AOI211XL U79 ( .A0(n329), .A1(n198), .B0(n71), .C0(n143), .Y(n72) );
  AOI31XL U80 ( .A0(n81), .A1(n80), .A2(n97), .B0(n321), .Y(n91) );
  OAI211XL U81 ( .A0(n350), .A1(n268), .B0(n141), .C0(n140), .Y(n142) );
  AOI211XL U82 ( .A0(n329), .A1(n162), .B0(n85), .C0(n84), .Y(n88) );
  AOI31XL U83 ( .A0(n364), .A1(n363), .A2(n362), .B0(n361), .Y(n365) );
  AOI31XL U84 ( .A0(n324), .A1(n323), .A2(n322), .B0(n321), .Y(n367) );
  AOI211XL U85 ( .A0(n350), .A1(n303), .B0(n185), .C0(n264), .Y(n186) );
  AOI2BB2XL U86 ( .B0(n264), .B1(n360), .A0N(n350), .A1N(n265), .Y(n283) );
  AOI211XL U87 ( .A0(n298), .A1(n179), .B0(n178), .C0(n177), .Y(n181) );
  NAND2XL U88 ( .A(n239), .B(n277), .Y(n188) );
  AOI211XL U89 ( .A0(n320), .A1(n1), .B0(n319), .C0(n318), .Y(n322) );
  AOI211XL U90 ( .A0(n360), .A1(n359), .B0(n358), .C0(n357), .Y(n362) );
  AOI22XL U91 ( .A0(n2), .A1(n227), .B0(n3), .B1(n226), .Y(n234) );
  AOI211XL U92 ( .A0(n4), .A1(n251), .B0(n250), .C0(n314), .Y(n263) );
  AOI221XL U93 ( .A0(n346), .A1(n330), .B0(n3), .B1(n269), .C0(n116), .Y(n117)
         );
  AOI211XL U94 ( .A0(n298), .A1(n290), .B0(n79), .C0(n78), .Y(n80) );
  AOI211XL U95 ( .A0(n2), .A1(n139), .B0(n138), .C0(n137), .Y(n140) );
  OAI211XL U96 ( .A0(n252), .A1(n336), .B0(n68), .C0(n67), .Y(n69) );
  AOI2BB2XL U97 ( .B0(n4), .B1(n337), .A0N(n350), .A1N(n179), .Y(n48) );
  AOI211XL U98 ( .A0(n329), .A1(n266), .B0(n216), .C0(n215), .Y(n218) );
  AOI22XL U99 ( .A0(n165), .A1(n2), .B0(n17), .B1(n268), .Y(n22) );
  AOI2BB2XL U100 ( .B0(n4), .B1(n86), .A0N(n237), .A1N(n104), .Y(n55) );
  NOR2XL U101 ( .A(n228), .B(n154), .Y(n120) );
  AOI2BB2XL U102 ( .B0(n2), .B1(n293), .A0N(n316), .A1N(n292), .Y(n301) );
  AOI22XL U103 ( .A0(n3), .A1(n134), .B0(n360), .B1(n266), .Y(n13) );
  AOI211XL U104 ( .A0(n298), .A1(n352), .B0(n297), .C0(n296), .Y(n300) );
  NAND2XL U105 ( .A(n268), .B(n349), .Y(n251) );
  AOI22XL U106 ( .A0(n1), .A1(n295), .B0(n298), .B1(n327), .Y(n15) );
  AOI22XL U107 ( .A0(n1), .A1(n24), .B0(n346), .B1(n320), .Y(n9) );
  AOI31XL U108 ( .A0(n2), .A1(n353), .A2(n352), .B0(n310), .Y(n323) );
  AOI22XL U109 ( .A0(n1), .A1(n307), .B0(n4), .B1(n42), .Y(n29) );
  AOI2BB2XL U110 ( .B0(n4), .B1(n104), .A0N(n196), .A1N(n103), .Y(n110) );
  NOR3XL U111 ( .A(n325), .B(n252), .C(n328), .Y(n253) );
  AOI22XL U112 ( .A0(n1), .A1(n293), .B0(n259), .B1(n268), .Y(n83) );
  AOI22XL U113 ( .A0(a[1]), .A1(n4), .B0(n1), .B1(n334), .Y(n219) );
  OAI22XL U114 ( .A0(n35), .A1(n328), .B0(n201), .B1(n155), .Y(n40) );
  AOI22XL U115 ( .A0(n1), .A1(n104), .B0(n326), .B1(n176), .Y(n38) );
  OAI22XL U116 ( .A0(n356), .A1(n354), .B0(n176), .B1(n184), .Y(n177) );
  AOI22XL U117 ( .A0(n330), .A1(n3), .B0(n298), .B1(n139), .Y(n68) );
  AOI22XL U118 ( .A0(n192), .A1(n276), .B0(n237), .B1(n316), .Y(n193) );
  AOI22XL U119 ( .A0(n96), .A1(n1), .B0(n4), .B1(n305), .Y(n81) );
  AOI22XL U120 ( .A0(n228), .A1(n329), .B0(n298), .B1(n103), .Y(n47) );
  AOI22XL U121 ( .A0(n3), .A1(n192), .B0(n360), .B1(n154), .Y(n161) );
  AOI22XL U122 ( .A0(n3), .A1(n44), .B0(n346), .B1(n290), .Y(n45) );
  AOI22XL U123 ( .A0(a[3]), .A1(n4), .B0(n1), .B1(n349), .Y(n363) );
  AOI22XL U124 ( .A0(n1), .A1(n214), .B0(n329), .B1(n268), .Y(n58) );
  AOI22XL U125 ( .A0(n4), .A1(n162), .B0(n329), .B1(n179), .Y(n170) );
  AOI211XL U126 ( .A0(a[2]), .A1(n134), .B0(n317), .C0(n133), .Y(n138) );
  AOI22XL U127 ( .A0(n1), .A1(n290), .B0(n346), .B1(n269), .Y(n157) );
  NOR2XL U128 ( .A(n185), .B(n99), .Y(n178) );
  AOI22XL U129 ( .A0(n1), .A1(n230), .B0(n252), .B1(n329), .Y(n233) );
  INVXL U130 ( .A(n156), .Y(n226) );
  AOI22XL U131 ( .A0(n3), .A1(n230), .B0(n4), .B1(n225), .Y(n203) );
  AOI22XL U132 ( .A0(a[3]), .A1(n346), .B0(n2), .B1(n202), .Y(n204) );
  INVXL U133 ( .A(n314), .Y(n315) );
  OAI2BB1XL U134 ( .A0N(n214), .A1N(n326), .B0(n247), .Y(n215) );
  NOR2XL U135 ( .A(n295), .B(n294), .Y(n296) );
  NAND2XL U136 ( .A(n353), .B(n352), .Y(n359) );
  AOI22XL U137 ( .A0(n3), .A1(n266), .B0(n329), .B1(n265), .Y(n282) );
  AOI22XL U138 ( .A0(n2), .A1(n292), .B0(n334), .B1(n4), .Y(n241) );
  AOI22XL U139 ( .A0(n330), .A1(n329), .B0(n2), .B1(n327), .Y(n343) );
  AOI22XL U140 ( .A0(n199), .A1(n333), .B0(n329), .B1(n345), .Y(n212) );
  INVXL U141 ( .A(n184), .Y(n187) );
  AOI22XL U142 ( .A0(n3), .A1(n347), .B0(n346), .B1(n345), .Y(n364) );
  OAI211XL U143 ( .A0(n277), .A1(n276), .B0(n275), .C0(n274), .Y(n279) );
  NAND2XL U144 ( .A(n2), .B(n269), .Y(n99) );
  AOI22XL U145 ( .A0(n298), .A1(n154), .B0(n4), .B1(n265), .Y(n8) );
  NOR2XL U146 ( .A(n154), .B(n332), .Y(n134) );
  AOI22XL U147 ( .A0(n3), .A1(n43), .B0(n346), .B1(n65), .Y(n23) );
  NAND2XL U148 ( .A(n107), .B(n256), .Y(n307) );
  AOI22XL U149 ( .A0(n2), .A1(n121), .B0(n329), .B1(n155), .Y(n28) );
  NOR2XL U150 ( .A(n165), .B(n311), .Y(n166) );
  INVXL U151 ( .A(n86), .Y(n176) );
  NAND3XL U152 ( .A(n3), .B(n144), .C(n86), .Y(n87) );
  NOR2XL U153 ( .A(n213), .B(n237), .Y(n259) );
  OAI22XL U154 ( .A0(n165), .A1(n303), .B0(n96), .B1(n237), .Y(n102) );
  AOI22XL U155 ( .A0(n298), .A1(n146), .B0(n4), .B1(n163), .Y(n89) );
  AOI22XL U156 ( .A0(n70), .A1(n154), .B0(n4), .B1(n266), .Y(n73) );
  AOI22XL U157 ( .A0(n189), .A1(n320), .B0(n2), .B1(n265), .Y(n114) );
  AOI211XL U158 ( .A0(n2), .A1(n271), .B0(n66), .C0(n297), .Y(n67) );
  NAND2XL U159 ( .A(n113), .B(n246), .Y(n139) );
  AOI22XL U160 ( .A0(n2), .A1(n96), .B0(n346), .B1(n5), .Y(n49) );
  AOI22XL U161 ( .A0(n2), .A1(n43), .B0(n360), .B1(n42), .Y(n46) );
  AOI22XL U162 ( .A0(n271), .A1(n4), .B0(n2), .B1(n155), .Y(n160) );
  AOI22XL U163 ( .A0(a[4]), .A1(n298), .B0(n346), .B1(n308), .Y(n25) );
  NOR2XL U164 ( .A(n295), .B(n230), .Y(n43) );
  NOR2XL U165 ( .A(n271), .B(n355), .Y(n17) );
  NAND2XL U166 ( .A(n4), .B(n249), .Y(n184) );
  OAI22XL U167 ( .A0(n327), .A1(n237), .B0(n201), .B1(n200), .Y(n206) );
  AOI22XL U168 ( .A0(n298), .A1(n132), .B0(n360), .B1(n308), .Y(n141) );
  NOR2XL U169 ( .A(n185), .B(n272), .Y(n317) );
  INVXL U170 ( .A(n135), .Y(n352) );
  AOI22XL U171 ( .A0(a[1]), .A1(n298), .B0(n3), .B1(n144), .Y(n153) );
  AOI22XL U172 ( .A0(n271), .A1(n360), .B0(n340), .B1(n332), .Y(n147) );
  AOI211XL U173 ( .A0(a[7]), .A1(n65), .B0(n191), .C0(n115), .Y(n66) );
  AOI31XL U174 ( .A0(n355), .A1(n237), .A2(n180), .B0(n330), .Y(n71) );
  AND2X2 U175 ( .A(n305), .B(n82), .Y(n225) );
  AOI22XL U176 ( .A0(n190), .A1(n360), .B0(n329), .B1(n107), .Y(n37) );
  NOR2XL U177 ( .A(n41), .B(n149), .Y(n103) );
  NAND2XL U178 ( .A(n313), .B(n200), .Y(n44) );
  AOI22XL U179 ( .A0(n230), .A1(n209), .B0(n360), .B1(n313), .Y(n10) );
  NOR3XL U180 ( .A(n185), .B(n264), .C(n311), .Y(n297) );
  AOI22XL U181 ( .A0(n185), .A1(n4), .B0(n329), .B1(n272), .Y(n100) );
  AOI22XL U182 ( .A0(n4), .A1(n353), .B0(n112), .B1(n111), .Y(n118) );
  OAI22XL U183 ( .A0(n355), .A1(n198), .B0(n308), .B1(n316), .Y(n119) );
  AOI22XL U184 ( .A0(n230), .A1(n4), .B0(n340), .B1(n356), .Y(n124) );
  NAND2XL U185 ( .A(n111), .B(n349), .Y(n179) );
  AOI22XL U186 ( .A0(n271), .A1(n326), .B0(n331), .B1(n270), .Y(n275) );
  AOI22XL U187 ( .A0(n334), .A1(n333), .B0(n332), .B1(n331), .Y(n335) );
  NOR2XL U188 ( .A(a[1]), .B(n330), .Y(n272) );
  NOR2XL U189 ( .A(n191), .B(n190), .Y(n292) );
  AOI22XL U190 ( .A0(n145), .A1(n333), .B0(n254), .B1(n331), .Y(n152) );
  NAND3XL U191 ( .A(n209), .B(n246), .C(n208), .Y(n210) );
  NAND2XL U192 ( .A(n313), .B(n305), .Y(n42) );
  NAND2XL U193 ( .A(n308), .B(n270), .Y(n65) );
  OR2X2 U194 ( .A(a[7]), .B(n115), .Y(n350) );
  NOR2XL U195 ( .A(n41), .B(a[1]), .Y(n199) );
  AOI22XL U196 ( .A0(n326), .A1(n325), .B0(n3), .B1(n5), .Y(n344) );
  NAND3XL U197 ( .A(n3), .B(a[3]), .C(n208), .Y(n77) );
  NOR2XL U198 ( .A(n237), .B(n332), .Y(n112) );
  AOI22XL U199 ( .A0(n191), .A1(n209), .B0(n329), .B1(n309), .Y(n16) );
  NOR2XL U200 ( .A(a[1]), .B(n252), .Y(n135) );
  NAND2XL U201 ( .A(a[1]), .B(n264), .Y(n305) );
  OR2X2 U202 ( .A(n267), .B(n196), .Y(n328) );
  NAND2XL U203 ( .A(n329), .B(n313), .Y(n354) );
  INVXL U204 ( .A(n201), .Y(n189) );
  INVXL U205 ( .A(n333), .Y(n238) );
  INVXL U206 ( .A(n299), .Y(n287) );
  NAND3XL U207 ( .A(n333), .B(n76), .C(n246), .Y(n75) );
  INVXL U208 ( .A(n196), .Y(n209) );
  NOR2XL U209 ( .A(n267), .B(n276), .Y(n331) );
  INVXL U210 ( .A(n277), .Y(n254) );
  AOI22XL U211 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n276), .Y(n136) );
  NOR2XL U212 ( .A(a[1]), .B(n202), .Y(n164) );
  NAND2XL U213 ( .A(a[2]), .B(n278), .Y(n196) );
  NAND2XL U214 ( .A(n267), .B(n278), .Y(n255) );
  AOI22XL U215 ( .A0(a[1]), .A1(a[7]), .B0(n267), .B1(n5), .Y(n76) );
  NOR2XL U216 ( .A(a[3]), .B(a[1]), .Y(n229) );
  NAND2XL U217 ( .A(a[3]), .B(a[1]), .Y(n24) );
  INVX2 U218 ( .A(a[4]), .Y(n202) );
  INVX2 U219 ( .A(a[2]), .Y(n276) );
  NAND2XL U220 ( .A(a[4]), .B(a[1]), .Y(n277) );
  NAND2X2 U221 ( .A(n278), .B(n276), .Y(n201) );
  NOR2X2 U222 ( .A(n35), .B(n202), .Y(n264) );
  NOR2X2 U223 ( .A(n41), .B(n5), .Y(n185) );
  NAND2X2 U224 ( .A(a[1]), .B(n246), .Y(n308) );
  NAND2X2 U225 ( .A(a[3]), .B(n202), .Y(n246) );
  NOR2X2 U226 ( .A(n276), .B(a[7]), .Y(n326) );
  NOR2X2 U227 ( .A(n252), .B(n330), .Y(n295) );
  NOR2X2 U228 ( .A(n330), .B(n5), .Y(n230) );
  NAND2X2 U229 ( .A(n202), .B(n5), .Y(n313) );
  CLKINVX3 U230 ( .A(n237), .Y(n360) );
  NAND2X2 U231 ( .A(a[5]), .B(n326), .Y(n237) );
  CLKINVX3 U232 ( .A(n350), .Y(n1) );
  NOR2X4 U233 ( .A(a[2]), .B(n133), .Y(n329) );
  BUFX3 U234 ( .A(n348), .Y(n3) );
  NOR2X4 U235 ( .A(a[7]), .B(n201), .Y(n298) );
  CLKINVX3 U236 ( .A(a[1]), .Y(n5) );
  CLKINVX3 U237 ( .A(n311), .Y(n346) );
  NAND2X2 U238 ( .A(n278), .B(n326), .Y(n311) );
  BUFX3 U239 ( .A(n351), .Y(n4) );
  AOI21XL U240 ( .A0(n313), .A1(n312), .B0(n311), .Y(n319) );
  AOI21XL U241 ( .A0(n309), .A1(n308), .B0(n336), .Y(n310) );
  AOI21XL U242 ( .A0(n360), .A1(n307), .B0(n306), .Y(n324) );
  AOI21XL U243 ( .A0(n305), .A1(n304), .B0(n303), .Y(n306) );
  AOI21XL U244 ( .A0(n4), .A1(n308), .B0(n3), .Y(n294) );
  AOI21XL U245 ( .A0(n213), .A1(n308), .B0(n328), .Y(n216) );
  AOI21XL U246 ( .A0(n270), .A1(n353), .B0(n311), .Y(n183) );
  AOI21XL U247 ( .A0(n329), .A1(n226), .B0(n158), .Y(n159) );
  AOI21XL U248 ( .A0(n136), .A1(n352), .B0(n311), .Y(n137) );
  AOI21XL U249 ( .A0(n240), .A1(n249), .B0(n328), .Y(n85) );
  AOI21XL U250 ( .A0(n209), .A1(n320), .B0(n346), .Y(n74) );
  AOI21XL U251 ( .A0(n54), .A1(n53), .B0(n361), .Y(n61) );
  AOI21XL U252 ( .A0(n240), .A1(n82), .B0(n316), .Y(n51) );
  AOI21XL U253 ( .A0(n360), .A1(n290), .B0(n26), .Y(n27) );
  AOI21XL U254 ( .A0(n146), .A1(n353), .B0(n336), .Y(n18) );
  AOI21XL U255 ( .A0(n2), .A1(n251), .B0(n52), .Y(n14) );
  AOI21XL U256 ( .A0(n313), .A1(n200), .B0(n336), .Y(n52) );
  AOI21XL U257 ( .A0(n269), .A1(n268), .B0(n267), .Y(n280) );
  AOI21XL U258 ( .A0(n254), .A1(n3), .B0(n253), .Y(n262) );
  AOI21XL U259 ( .A0(n346), .A1(n347), .B0(n242), .Y(n243) );
  NOR2X1 U260 ( .A(n276), .B(n133), .Y(n348) );
  NOR2X1 U261 ( .A(n267), .B(n201), .Y(n351) );
  INVX1 U262 ( .A(a[7]), .Y(n267) );
  OAI21XL U263 ( .A0(n224), .A1(n341), .B0(n223), .Y(d[2]) );
  OAI21XL U264 ( .A0(n175), .A1(n361), .B0(n174), .Y(d[3]) );
  OAI21XL U265 ( .A0(n95), .A1(n361), .B0(n94), .Y(d[5]) );
  OAI21XL U266 ( .A0(n64), .A1(n299), .B0(n63), .Y(d[6]) );
  OAI21XL U267 ( .A0(n34), .A1(n361), .B0(n33), .Y(d[7]) );
  OAI21XL U268 ( .A0(n131), .A1(n299), .B0(n130), .Y(d[4]) );
  OAI21XL U269 ( .A0(n289), .A1(n321), .B0(n288), .Y(d[1]) );
  NAND2X1 U270 ( .A(a[7]), .B(a[5]), .Y(n133) );
  NOR2X1 U271 ( .A(n5), .B(n246), .Y(n214) );
  NAND2X1 U272 ( .A(a[4]), .B(n35), .Y(n269) );
  NOR2X1 U273 ( .A(a[4]), .B(n5), .Y(n273) );
  OAI21XL U274 ( .A0(n273), .A1(n229), .B0(n3), .Y(n7) );
  NOR2X1 U275 ( .A(a[7]), .B(a[2]), .Y(n340) );
  INVX1 U276 ( .A(n246), .Y(n252) );
  OAI21XL U277 ( .A0(n70), .A1(n340), .B0(n135), .Y(n6) );
  NAND3X1 U278 ( .A(n99), .B(n7), .C(n6), .Y(n12) );
  INVX1 U279 ( .A(n70), .Y(n115) );
  NOR2X1 U280 ( .A(n264), .B(n5), .Y(n325) );
  NAND3X1 U281 ( .A(n10), .B(n9), .C(n8), .Y(n11) );
  AOI211X1 U282 ( .A0(n329), .A1(n214), .B0(n12), .C0(n11), .Y(n34) );
  INVX1 U283 ( .A(a[6]), .Y(n20) );
  NOR2X1 U284 ( .A(a[0]), .B(n20), .Y(n129) );
  INVX1 U285 ( .A(n264), .Y(n309) );
  INVX1 U286 ( .A(n24), .Y(n327) );
  NAND2X1 U287 ( .A(n264), .B(n5), .Y(n349) );
  INVX1 U288 ( .A(n191), .Y(n200) );
  INVX1 U289 ( .A(n4), .Y(n336) );
  NAND2X1 U290 ( .A(n35), .B(n202), .Y(n107) );
  NAND2X1 U291 ( .A(n24), .B(n249), .Y(n266) );
  NAND4X1 U292 ( .A(n16), .B(n15), .C(n14), .D(n13), .Y(n32) );
  NAND2X1 U293 ( .A(a[3]), .B(n5), .Y(n270) );
  INVX1 U294 ( .A(n107), .Y(n41) );
  NOR2X1 U295 ( .A(n199), .B(n273), .Y(n165) );
  INVX1 U296 ( .A(n313), .Y(n271) );
  INVX1 U297 ( .A(n295), .Y(n213) );
  NOR2X1 U298 ( .A(a[1]), .B(n213), .Y(n228) );
  INVX1 U299 ( .A(n228), .Y(n239) );
  NAND2X1 U300 ( .A(n5), .B(n309), .Y(n144) );
  NOR2BX1 U301 ( .AN(n144), .B(n185), .Y(n96) );
  INVX1 U302 ( .A(n199), .Y(n146) );
  NAND2X1 U303 ( .A(a[0]), .B(n20), .Y(n299) );
  INVX1 U304 ( .A(n230), .Y(n256) );
  NAND2X1 U305 ( .A(n200), .B(n349), .Y(n121) );
  NAND2X1 U306 ( .A(n309), .B(n86), .Y(n290) );
  INVX1 U307 ( .A(n3), .Y(n303) );
  NAND2X1 U308 ( .A(n239), .B(n353), .Y(n105) );
  OAI21XL U309 ( .A0(n303), .A1(n105), .B0(n25), .Y(n26) );
  NOR2X1 U310 ( .A(a[6]), .B(a[0]), .Y(n93) );
  INVX1 U311 ( .A(n185), .Y(n113) );
  INVX1 U312 ( .A(n229), .Y(n304) );
  NAND2X1 U313 ( .A(n113), .B(n304), .Y(n104) );
  OAI21XL U314 ( .A0(n273), .A1(n164), .B0(n3), .Y(n36) );
  NAND4BXL U315 ( .AN(n250), .B(n38), .C(n37), .D(n36), .Y(n39) );
  INVX1 U316 ( .A(n353), .Y(n145) );
  NOR2X1 U317 ( .A(n145), .B(n332), .Y(n337) );
  INVX1 U318 ( .A(n273), .Y(n111) );
  INVX1 U319 ( .A(n308), .Y(n149) );
  NAND4X1 U320 ( .A(n48), .B(n47), .C(n46), .D(n45), .Y(n62) );
  INVX1 U321 ( .A(n214), .Y(n240) );
  INVX1 U322 ( .A(n332), .Y(n82) );
  INVX1 U323 ( .A(n329), .Y(n316) );
  OAI21XL U324 ( .A0(a[4]), .A1(n350), .B0(n49), .Y(n50) );
  NAND2X1 U325 ( .A(n313), .B(n256), .Y(n293) );
  NOR2X1 U326 ( .A(n355), .B(n293), .Y(n167) );
  OAI21XL U327 ( .A0(n325), .A1(n229), .B0(n298), .Y(n59) );
  OAI21XL U328 ( .A0(n120), .A1(n303), .B0(n55), .Y(n56) );
  NAND2X1 U329 ( .A(n270), .B(n312), .Y(n227) );
  INVX1 U330 ( .A(n190), .Y(n198) );
  NAND2X1 U331 ( .A(n3), .B(n313), .Y(n180) );
  NOR2X1 U332 ( .A(n350), .B(n313), .Y(n143) );
  NOR2X1 U333 ( .A(n278), .B(n276), .Y(n333) );
  OAI21XL U334 ( .A0(n353), .A1(n328), .B0(n75), .Y(n79) );
  INVX1 U335 ( .A(n76), .Y(n208) );
  OAI21XL U336 ( .A0(n225), .A1(n316), .B0(n77), .Y(n78) );
  NAND2X1 U337 ( .A(n346), .B(n213), .Y(n97) );
  INVX1 U338 ( .A(n129), .Y(n321) );
  NAND2X1 U339 ( .A(n111), .B(n270), .Y(n163) );
  OAI21XL U340 ( .A0(n120), .A1(n311), .B0(n83), .Y(n84) );
  NOR2X1 U341 ( .A(n149), .B(n320), .Y(n156) );
  NAND4X1 U342 ( .A(n100), .B(n99), .C(n98), .D(n97), .Y(n101) );
  AOI211X1 U343 ( .A0(n1), .A1(n156), .B0(n102), .C0(n101), .Y(n131) );
  OAI21XL U344 ( .A0(n252), .A1(n350), .B0(n180), .Y(n106) );
  NOR2X1 U345 ( .A(n107), .B(n5), .Y(n356) );
  OAI21XL U346 ( .A0(n190), .A1(n356), .B0(n329), .Y(n108) );
  NAND4BXL U347 ( .AN(n112), .B(n110), .C(n109), .D(n108), .Y(n128) );
  OAI21XL U348 ( .A0(n115), .A1(n197), .B0(n114), .Y(n116) );
  NAND2X1 U349 ( .A(n298), .B(n230), .Y(n247) );
  INVX1 U350 ( .A(n120), .Y(n207) );
  INVX1 U351 ( .A(n121), .Y(n192) );
  OAI21XL U352 ( .A0(n198), .A1(n238), .B0(n237), .Y(n122) );
  OAI21XL U353 ( .A0(a[1]), .A1(n136), .B0(n308), .Y(n132) );
  NOR2X1 U354 ( .A(n328), .B(n146), .Y(n358) );
  OAI21XL U355 ( .A0(n311), .A1(n304), .B0(n147), .Y(n148) );
  OAI21XL U356 ( .A0(n330), .A1(n149), .B0(n329), .Y(n150) );
  NAND4X1 U357 ( .A(n153), .B(n152), .C(n151), .D(n150), .Y(n173) );
  OAI21XL U358 ( .A0(n213), .A1(n255), .B0(n157), .Y(n158) );
  AOI211X1 U359 ( .A0(n287), .A1(n173), .B0(n172), .C0(n171), .Y(n174) );
  OAI21XL U360 ( .A0(n292), .A1(n276), .B0(n193), .Y(n194) );
  OAI21XL U361 ( .A0(n204), .A1(n208), .B0(n203), .Y(n205) );
  OAI21XL U362 ( .A0(n320), .A1(n356), .B0(n3), .Y(n217) );
  NOR2X1 U363 ( .A(n225), .B(n336), .Y(n236) );
  OAI21XL U364 ( .A0(n228), .A1(n273), .B0(n346), .Y(n232) );
  OAI21XL U365 ( .A0(n230), .A1(n229), .B0(n360), .Y(n231) );
  NAND4X1 U366 ( .A(n234), .B(n233), .C(n232), .D(n231), .Y(n235) );
  AOI211X1 U367 ( .A0(n337), .A1(n298), .B0(n236), .C0(n235), .Y(n289) );
  OAI21XL U368 ( .A0(n239), .A1(n238), .B0(n237), .Y(n245) );
  OAI21XL U369 ( .A0(n330), .A1(n316), .B0(n241), .Y(n242) );
  OAI21XL U370 ( .A0(n350), .A1(n347), .B0(n243), .Y(n244) );
  NOR2X1 U371 ( .A(n355), .B(n304), .Y(n314) );
  OAI21XL U372 ( .A0(n273), .A1(n272), .B0(n340), .Y(n274) );
  OAI21XL U373 ( .A0(n280), .A1(n279), .B0(n278), .Y(n281) );
  OAI21XL U374 ( .A0(n317), .A1(n316), .B0(n315), .Y(n318) );
  OAI21XL U375 ( .A0(n337), .A1(n336), .B0(n335), .Y(n338) );
  OAI21XL U376 ( .A0(n356), .A1(n355), .B0(n354), .Y(n357) );
endmodule


module aes_sbox_2 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368;

  INVX1 U1 ( .A(n93), .Y(n341) );
  NOR2BX1 U2 ( .AN(n349), .B(n311), .Y(n250) );
  AOI211XL U3 ( .A0(n287), .A1(n286), .B0(n285), .C0(n284), .Y(n288) );
  AOI31XL U4 ( .A0(n263), .A1(n262), .A2(n261), .B0(n341), .Y(n285) );
  AOI211X1 U5 ( .A0(n287), .A1(n222), .B0(n221), .C0(n220), .Y(n223) );
  NAND2XL U6 ( .A(n239), .B(n268), .Y(n339) );
  INVX1 U7 ( .A(n325), .Y(n268) );
  INVX1 U8 ( .A(n353), .Y(n145) );
  NOR2X1 U9 ( .A(a[2]), .B(n278), .Y(n70) );
  AOI31XL U10 ( .A0(n29), .A1(n28), .A2(n27), .B0(n341), .Y(n30) );
  AOI211X1 U11 ( .A0(n1), .A1(n308), .B0(n183), .C0(n182), .Y(n224) );
  AOI31XL U12 ( .A0(n125), .A1(n124), .A2(n123), .B0(n341), .Y(n126) );
  AOI2BB2XL U13 ( .B0(n360), .B1(n291), .A0N(n350), .A1N(n290), .Y(n302) );
  AOI21XL U14 ( .A0(n340), .A1(n339), .B0(n338), .Y(n342) );
  AOI211XL U15 ( .A0(n189), .A1(n188), .B0(n187), .C0(n186), .Y(n195) );
  INVXL U16 ( .A(n260), .Y(n291) );
  NOR2XL U17 ( .A(n228), .B(n327), .Y(n260) );
  INVXL U18 ( .A(n154), .Y(n312) );
  AOI32XL U19 ( .A0(n113), .A1(a[7]), .A2(n269), .B0(n163), .B1(n267), .Y(n197) );
  NAND2XL U20 ( .A(n113), .B(n82), .Y(n162) );
  NAND2XL U21 ( .A(a[1]), .B(n295), .Y(n86) );
  NAND2XL U22 ( .A(n144), .B(n24), .Y(n155) );
  AOI2BB2XL U23 ( .B0(n360), .B1(n164), .A0N(n303), .A1N(n163), .Y(n169) );
  NAND2XL U24 ( .A(n198), .B(n277), .Y(n345) );
  NOR2X1 U25 ( .A(a[1]), .B(n295), .Y(n320) );
  NAND2XL U26 ( .A(n313), .B(n240), .Y(n347) );
  NOR2XL U27 ( .A(n325), .B(n135), .Y(n265) );
  NOR2X1 U28 ( .A(n295), .B(n5), .Y(n154) );
  CLKINVX3 U29 ( .A(n328), .Y(n2) );
  INVX1 U30 ( .A(n298), .Y(n355) );
  NAND2XL U31 ( .A(n330), .B(n5), .Y(n249) );
  INVXL U32 ( .A(n270), .Y(n334) );
  NOR2XL U33 ( .A(n5), .B(n269), .Y(n191) );
  NOR2X1 U34 ( .A(a[1]), .B(n107), .Y(n332) );
  CLKINVX3 U35 ( .A(n269), .Y(n330) );
  NOR2XL U36 ( .A(a[1]), .B(n246), .Y(n190) );
  NAND2X1 U37 ( .A(a[1]), .B(n35), .Y(n353) );
  INVX1 U38 ( .A(a[3]), .Y(n35) );
  NAND2X1 U39 ( .A(a[6]), .B(a[0]), .Y(n361) );
  AOI211XL U40 ( .A0(n129), .A1(n128), .B0(n127), .C0(n126), .Y(n130) );
  AOI211XL U41 ( .A0(n129), .A1(n32), .B0(n31), .C0(n30), .Y(n33) );
  AOI31XL U42 ( .A0(n23), .A1(n22), .A2(n21), .B0(n299), .Y(n31) );
  AOI211XL U43 ( .A0(n93), .A1(n92), .B0(n91), .C0(n90), .Y(n94) );
  AOI211XL U44 ( .A0(n129), .A1(n62), .B0(n61), .C0(n60), .Y(n63) );
  OAI211XL U45 ( .A0(n249), .A1(n355), .B0(n248), .C0(n247), .Y(n286) );
  AOI211XL U46 ( .A0(n329), .A1(n260), .B0(n259), .C0(n258), .Y(n261) );
  OR4X2 U47 ( .A(n368), .B(n367), .C(n366), .D(n365), .Y(d[0]) );
  AOI31XL U48 ( .A0(n212), .A1(n211), .A2(n210), .B0(n361), .Y(n221) );
  AOI211XL U49 ( .A0(n260), .A1(n360), .B0(n19), .C0(n18), .Y(n21) );
  AOI211XL U50 ( .A0(n192), .A1(n4), .B0(n143), .C0(n142), .Y(n175) );
  AOI31XL U51 ( .A0(n344), .A1(n343), .A2(n342), .B0(n341), .Y(n366) );
  AOI31XL U52 ( .A0(n302), .A1(n301), .A2(n300), .B0(n299), .Y(n368) );
  AOI31XL U53 ( .A0(n246), .A1(n256), .A2(n245), .B0(n244), .Y(n248) );
  OAI22XL U54 ( .A0(n257), .A1(n350), .B0(n256), .B1(n255), .Y(n258) );
  OAI211XL U55 ( .A0(n197), .A1(n196), .B0(n195), .C0(n194), .Y(n222) );
  AOI31XL U56 ( .A0(n161), .A1(n160), .A2(n159), .B0(n321), .Y(n172) );
  AOI22XL U57 ( .A0(n257), .A1(n298), .B0(n268), .B1(n106), .Y(n109) );
  AOI31XL U58 ( .A0(n89), .A1(n88), .A2(n87), .B0(n299), .Y(n90) );
  AOI31XL U59 ( .A0(n170), .A1(n169), .A2(n168), .B0(n341), .Y(n171) );
  OAI211XL U60 ( .A0(n74), .A1(n121), .B0(n73), .C0(n72), .Y(n92) );
  AOI31XL U61 ( .A0(n59), .A1(n58), .A2(n57), .B0(n341), .Y(n60) );
  AOI31XL U62 ( .A0(n364), .A1(n363), .A2(n362), .B0(n361), .Y(n365) );
  AOI21X1 U63 ( .A0(n360), .A1(n227), .B0(n69), .Y(n95) );
  AOI22XL U64 ( .A0(n2), .A1(n207), .B0(n192), .B1(n122), .Y(n123) );
  AOI211XL U65 ( .A0(n346), .A1(n268), .B0(n143), .C0(n119), .Y(n125) );
  AOI31XL U66 ( .A0(n118), .A1(n117), .A2(n247), .B0(n361), .Y(n127) );
  INVXL U67 ( .A(n105), .Y(n257) );
  NAND2XL U68 ( .A(n298), .B(n105), .Y(n98) );
  AOI211XL U69 ( .A0(n2), .A1(n291), .B0(n167), .C0(n166), .Y(n168) );
  AOI211XL U70 ( .A0(n4), .A1(n339), .B0(n358), .C0(n148), .Y(n151) );
  OAI211XL U71 ( .A0(n350), .A1(n268), .B0(n141), .C0(n140), .Y(n142) );
  AOI31XL U72 ( .A0(n219), .A1(n218), .A2(n217), .B0(n321), .Y(n220) );
  AOI211XL U73 ( .A0(a[7]), .A1(n339), .B0(n96), .C0(n115), .Y(n19) );
  AOI211XL U74 ( .A0(n250), .A1(n240), .B0(n178), .C0(n56), .Y(n57) );
  AOI211XL U75 ( .A0(n326), .A1(n188), .B0(n52), .C0(n167), .Y(n53) );
  AOI211XL U76 ( .A0(n3), .A1(n86), .B0(n51), .C0(n50), .Y(n54) );
  AOI211XL U77 ( .A0(n298), .A1(n105), .B0(n40), .C0(n39), .Y(n64) );
  AOI211XL U78 ( .A0(n329), .A1(n162), .B0(n85), .C0(n84), .Y(n88) );
  AOI31XL U79 ( .A0(n81), .A1(n80), .A2(n97), .B0(n321), .Y(n91) );
  AOI211XL U80 ( .A0(n329), .A1(n198), .B0(n71), .C0(n143), .Y(n72) );
  OAI211XL U81 ( .A0(n337), .A1(n237), .B0(n181), .C0(n180), .Y(n182) );
  AOI31XL U82 ( .A0(n324), .A1(n323), .A2(n322), .B0(n321), .Y(n367) );
  AOI211XL U83 ( .A0(n1), .A1(n207), .B0(n206), .C0(n205), .Y(n211) );
  AOI31XL U84 ( .A0(n283), .A1(n282), .A2(n281), .B0(n361), .Y(n284) );
  AOI221XL U85 ( .A0(n346), .A1(n330), .B0(n3), .B1(n269), .C0(n116), .Y(n117)
         );
  AOI211XL U86 ( .A0(n360), .A1(n359), .B0(n358), .C0(n357), .Y(n362) );
  AOI211XL U87 ( .A0(n320), .A1(n1), .B0(n319), .C0(n318), .Y(n322) );
  AOI22XL U88 ( .A0(n2), .A1(n227), .B0(n3), .B1(n226), .Y(n234) );
  AOI211XL U89 ( .A0(n4), .A1(n251), .B0(n250), .C0(n314), .Y(n263) );
  AOI2BB2XL U90 ( .B0(n264), .B1(n360), .A0N(n350), .A1N(n265), .Y(n283) );
  AOI211XL U91 ( .A0(n298), .A1(n179), .B0(n178), .C0(n177), .Y(n181) );
  AOI211XL U92 ( .A0(n350), .A1(n303), .B0(n185), .C0(n264), .Y(n186) );
  AOI211XL U93 ( .A0(n329), .A1(n266), .B0(n216), .C0(n215), .Y(n218) );
  AOI211XL U94 ( .A0(n2), .A1(n139), .B0(n138), .C0(n137), .Y(n140) );
  AOI211XL U95 ( .A0(n298), .A1(n290), .B0(n79), .C0(n78), .Y(n80) );
  AOI2BB2XL U96 ( .B0(n4), .B1(n337), .A0N(n350), .A1N(n179), .Y(n48) );
  NAND2XL U97 ( .A(n239), .B(n277), .Y(n188) );
  OAI211XL U98 ( .A0(n252), .A1(n336), .B0(n68), .C0(n67), .Y(n69) );
  AOI22XL U99 ( .A0(n3), .A1(n192), .B0(n360), .B1(n154), .Y(n161) );
  AOI22XL U100 ( .A0(a[1]), .A1(n4), .B0(n1), .B1(n334), .Y(n219) );
  NOR2XL U101 ( .A(n185), .B(n99), .Y(n178) );
  INVXL U102 ( .A(n156), .Y(n226) );
  AOI2BB2XL U103 ( .B0(n4), .B1(n104), .A0N(n196), .A1N(n103), .Y(n110) );
  AOI211XL U104 ( .A0(a[2]), .A1(n134), .B0(n317), .C0(n133), .Y(n138) );
  AOI22XL U105 ( .A0(n1), .A1(n290), .B0(n346), .B1(n269), .Y(n157) );
  AOI22XL U106 ( .A0(n4), .A1(n162), .B0(n329), .B1(n179), .Y(n170) );
  AOI22XL U107 ( .A0(n1), .A1(n307), .B0(n4), .B1(n42), .Y(n29) );
  AOI22XL U108 ( .A0(n1), .A1(n293), .B0(n259), .B1(n268), .Y(n83) );
  AOI22XL U109 ( .A0(n165), .A1(n2), .B0(n17), .B1(n268), .Y(n22) );
  OAI22XL U110 ( .A0(n35), .A1(n328), .B0(n201), .B1(n155), .Y(n40) );
  AOI22XL U111 ( .A0(n3), .A1(n134), .B0(n360), .B1(n266), .Y(n13) );
  AOI22XL U112 ( .A0(n1), .A1(n104), .B0(n326), .B1(n176), .Y(n38) );
  NAND2XL U113 ( .A(n268), .B(n349), .Y(n251) );
  AOI22XL U114 ( .A0(n1), .A1(n295), .B0(n298), .B1(n327), .Y(n15) );
  AOI22XL U115 ( .A0(n1), .A1(n230), .B0(n252), .B1(n329), .Y(n233) );
  AOI22XL U116 ( .A0(n228), .A1(n329), .B0(n298), .B1(n103), .Y(n47) );
  AOI22XL U117 ( .A0(n1), .A1(n24), .B0(n346), .B1(n320), .Y(n9) );
  AOI22XL U118 ( .A0(n3), .A1(n44), .B0(n346), .B1(n290), .Y(n45) );
  AOI22XL U119 ( .A0(a[3]), .A1(n4), .B0(n1), .B1(n349), .Y(n363) );
  AOI2BB2XL U120 ( .B0(n2), .B1(n293), .A0N(n316), .A1N(n292), .Y(n301) );
  AOI211XL U121 ( .A0(n298), .A1(n352), .B0(n297), .C0(n296), .Y(n300) );
  AOI2BB2XL U122 ( .B0(n4), .B1(n86), .A0N(n237), .A1N(n104), .Y(n55) );
  AOI31XL U123 ( .A0(n2), .A1(n353), .A2(n352), .B0(n310), .Y(n323) );
  AOI22XL U124 ( .A0(n1), .A1(n214), .B0(n329), .B1(n268), .Y(n58) );
  NOR2XL U125 ( .A(n228), .B(n154), .Y(n120) );
  AOI22XL U126 ( .A0(n192), .A1(n276), .B0(n237), .B1(n316), .Y(n193) );
  AOI22XL U127 ( .A0(n330), .A1(n3), .B0(n298), .B1(n139), .Y(n68) );
  OAI22XL U128 ( .A0(n356), .A1(n354), .B0(n176), .B1(n184), .Y(n177) );
  AOI22XL U129 ( .A0(n96), .A1(n1), .B0(n4), .B1(n305), .Y(n81) );
  NOR3XL U130 ( .A(n325), .B(n252), .C(n328), .Y(n253) );
  NOR2XL U131 ( .A(n295), .B(n294), .Y(n296) );
  INVXL U132 ( .A(n314), .Y(n315) );
  AOI22XL U133 ( .A0(n330), .A1(n329), .B0(n2), .B1(n327), .Y(n343) );
  AOI22XL U134 ( .A0(n3), .A1(n347), .B0(n346), .B1(n345), .Y(n364) );
  NAND2XL U135 ( .A(n353), .B(n352), .Y(n359) );
  AOI22XL U136 ( .A0(n2), .A1(n292), .B0(n334), .B1(n4), .Y(n241) );
  AOI22XL U137 ( .A0(n3), .A1(n266), .B0(n329), .B1(n265), .Y(n282) );
  OAI211XL U138 ( .A0(n277), .A1(n276), .B0(n275), .C0(n274), .Y(n279) );
  INVXL U139 ( .A(n184), .Y(n187) );
  AOI22XL U140 ( .A0(n199), .A1(n333), .B0(n329), .B1(n345), .Y(n212) );
  AOI22XL U141 ( .A0(a[3]), .A1(n346), .B0(n2), .B1(n202), .Y(n204) );
  AOI22XL U142 ( .A0(n3), .A1(n230), .B0(n4), .B1(n225), .Y(n203) );
  OAI2BB1XL U143 ( .A0N(n214), .A1N(n326), .B0(n247), .Y(n215) );
  AOI22XL U144 ( .A0(n2), .A1(n96), .B0(n346), .B1(n5), .Y(n49) );
  NAND2XL U145 ( .A(n2), .B(n269), .Y(n99) );
  AOI22XL U146 ( .A0(n298), .A1(n154), .B0(n4), .B1(n265), .Y(n8) );
  NOR2XL U147 ( .A(n154), .B(n332), .Y(n134) );
  AOI22XL U148 ( .A0(n2), .A1(n43), .B0(n360), .B1(n42), .Y(n46) );
  AOI22XL U149 ( .A0(n3), .A1(n43), .B0(n346), .B1(n65), .Y(n23) );
  NAND2XL U150 ( .A(n107), .B(n256), .Y(n307) );
  AOI22XL U151 ( .A0(n2), .A1(n121), .B0(n329), .B1(n155), .Y(n28) );
  AOI22XL U152 ( .A0(n271), .A1(n4), .B0(n2), .B1(n155), .Y(n160) );
  NOR2XL U153 ( .A(n165), .B(n311), .Y(n166) );
  OAI22XL U154 ( .A0(n165), .A1(n303), .B0(n96), .B1(n237), .Y(n102) );
  AOI22XL U155 ( .A0(n189), .A1(n320), .B0(n2), .B1(n265), .Y(n114) );
  NAND2XL U156 ( .A(n113), .B(n246), .Y(n139) );
  AOI211XL U157 ( .A0(n2), .A1(n271), .B0(n66), .C0(n297), .Y(n67) );
  AOI22XL U158 ( .A0(n70), .A1(n154), .B0(n4), .B1(n266), .Y(n73) );
  AOI22XL U159 ( .A0(n298), .A1(n146), .B0(n4), .B1(n163), .Y(n89) );
  NOR2XL U160 ( .A(n213), .B(n237), .Y(n259) );
  NAND3XL U161 ( .A(n3), .B(n144), .C(n86), .Y(n87) );
  INVXL U162 ( .A(n86), .Y(n176) );
  AND2X2 U163 ( .A(n305), .B(n82), .Y(n225) );
  NOR3XL U164 ( .A(n185), .B(n264), .C(n311), .Y(n297) );
  AOI31XL U165 ( .A0(n355), .A1(n237), .A2(n180), .B0(n330), .Y(n71) );
  NOR2XL U166 ( .A(n41), .B(n149), .Y(n103) );
  AOI22XL U167 ( .A0(n190), .A1(n360), .B0(n329), .B1(n107), .Y(n37) );
  NAND2XL U168 ( .A(n313), .B(n200), .Y(n44) );
  OAI22XL U169 ( .A0(n327), .A1(n237), .B0(n201), .B1(n200), .Y(n206) );
  AOI22XL U170 ( .A0(n230), .A1(n209), .B0(n360), .B1(n313), .Y(n10) );
  AOI22XL U171 ( .A0(n185), .A1(n4), .B0(n329), .B1(n272), .Y(n100) );
  AOI22XL U172 ( .A0(n298), .A1(n132), .B0(n360), .B1(n308), .Y(n141) );
  NOR2XL U173 ( .A(n185), .B(n272), .Y(n317) );
  INVXL U174 ( .A(n135), .Y(n352) );
  AOI22XL U175 ( .A0(a[1]), .A1(n298), .B0(n3), .B1(n144), .Y(n153) );
  NOR2XL U176 ( .A(n271), .B(n355), .Y(n17) );
  AOI22XL U177 ( .A0(n271), .A1(n360), .B0(n340), .B1(n332), .Y(n147) );
  NOR2XL U178 ( .A(n295), .B(n230), .Y(n43) );
  AOI211XL U179 ( .A0(a[7]), .A1(n65), .B0(n191), .C0(n115), .Y(n66) );
  AOI22XL U180 ( .A0(a[4]), .A1(n298), .B0(n346), .B1(n308), .Y(n25) );
  AOI22XL U181 ( .A0(n230), .A1(n4), .B0(n340), .B1(n356), .Y(n124) );
  OAI22XL U182 ( .A0(n355), .A1(n198), .B0(n308), .B1(n316), .Y(n119) );
  AOI22XL U183 ( .A0(n4), .A1(n353), .B0(n112), .B1(n111), .Y(n118) );
  NAND2XL U184 ( .A(n4), .B(n249), .Y(n184) );
  NAND2XL U185 ( .A(n308), .B(n270), .Y(n65) );
  NOR2XL U186 ( .A(a[1]), .B(n252), .Y(n135) );
  AOI22XL U187 ( .A0(n191), .A1(n209), .B0(n329), .B1(n309), .Y(n16) );
  AOI22XL U188 ( .A0(n145), .A1(n333), .B0(n254), .B1(n331), .Y(n152) );
  OR2X2 U189 ( .A(a[7]), .B(n115), .Y(n350) );
  NAND3XL U190 ( .A(n209), .B(n246), .C(n208), .Y(n210) );
  NAND2XL U191 ( .A(n313), .B(n305), .Y(n42) );
  AOI22XL U192 ( .A0(n271), .A1(n326), .B0(n331), .B1(n270), .Y(n275) );
  NOR2XL U193 ( .A(n41), .B(a[1]), .Y(n199) );
  NOR2XL U194 ( .A(n191), .B(n190), .Y(n292) );
  NOR2XL U195 ( .A(a[1]), .B(n330), .Y(n272) );
  NOR2XL U196 ( .A(n237), .B(n332), .Y(n112) );
  NAND2XL U197 ( .A(n111), .B(n349), .Y(n179) );
  AOI22XL U198 ( .A0(n334), .A1(n333), .B0(n332), .B1(n331), .Y(n335) );
  NAND3XL U199 ( .A(n3), .B(a[3]), .C(n208), .Y(n77) );
  AOI22XL U200 ( .A0(n326), .A1(n325), .B0(n3), .B1(n5), .Y(n344) );
  NAND2XL U201 ( .A(n329), .B(n313), .Y(n354) );
  INVXL U202 ( .A(n201), .Y(n189) );
  INVXL U203 ( .A(n333), .Y(n238) );
  INVXL U204 ( .A(n299), .Y(n287) );
  NAND3XL U205 ( .A(n333), .B(n76), .C(n246), .Y(n75) );
  OR2X2 U206 ( .A(n267), .B(n196), .Y(n328) );
  NAND2XL U207 ( .A(a[1]), .B(n264), .Y(n305) );
  INVXL U208 ( .A(n196), .Y(n209) );
  NOR2XL U209 ( .A(n267), .B(n276), .Y(n331) );
  INVXL U210 ( .A(n277), .Y(n254) );
  AOI22XL U211 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n276), .Y(n136) );
  AOI22XL U212 ( .A0(a[1]), .A1(a[7]), .B0(n267), .B1(n5), .Y(n76) );
  NAND2XL U213 ( .A(a[2]), .B(n278), .Y(n196) );
  NOR2XL U214 ( .A(a[1]), .B(n202), .Y(n164) );
  NAND2XL U215 ( .A(n267), .B(n278), .Y(n255) );
  INVX2 U216 ( .A(a[4]), .Y(n202) );
  INVX2 U217 ( .A(a[2]), .Y(n276) );
  INVX2 U218 ( .A(a[5]), .Y(n278) );
  NAND2XL U219 ( .A(a[3]), .B(a[1]), .Y(n24) );
  NOR2XL U220 ( .A(a[3]), .B(a[1]), .Y(n229) );
  NAND2XL U221 ( .A(a[4]), .B(a[1]), .Y(n277) );
  NAND2X2 U222 ( .A(n278), .B(n276), .Y(n201) );
  NOR2X2 U223 ( .A(n35), .B(n202), .Y(n264) );
  NOR2X2 U224 ( .A(n41), .B(n5), .Y(n185) );
  NAND2X2 U225 ( .A(a[1]), .B(n246), .Y(n308) );
  NAND2X2 U226 ( .A(a[3]), .B(n202), .Y(n246) );
  NOR2X2 U227 ( .A(n276), .B(a[7]), .Y(n326) );
  NOR2X2 U228 ( .A(n252), .B(n330), .Y(n295) );
  NOR2X2 U229 ( .A(n330), .B(n5), .Y(n230) );
  NAND2X2 U230 ( .A(n202), .B(n5), .Y(n313) );
  CLKINVX3 U231 ( .A(n237), .Y(n360) );
  NAND2X2 U232 ( .A(a[5]), .B(n326), .Y(n237) );
  CLKINVX3 U233 ( .A(n350), .Y(n1) );
  NOR2X4 U234 ( .A(a[2]), .B(n133), .Y(n329) );
  BUFX3 U235 ( .A(n348), .Y(n3) );
  NOR2X4 U236 ( .A(a[7]), .B(n201), .Y(n298) );
  CLKINVX3 U237 ( .A(a[1]), .Y(n5) );
  CLKINVX3 U238 ( .A(n311), .Y(n346) );
  NAND2X2 U239 ( .A(n278), .B(n326), .Y(n311) );
  BUFX3 U240 ( .A(n351), .Y(n4) );
  AOI21XL U241 ( .A0(n313), .A1(n312), .B0(n311), .Y(n319) );
  AOI21XL U242 ( .A0(n309), .A1(n308), .B0(n336), .Y(n310) );
  AOI21XL U243 ( .A0(n360), .A1(n307), .B0(n306), .Y(n324) );
  AOI21XL U244 ( .A0(n305), .A1(n304), .B0(n303), .Y(n306) );
  AOI21XL U245 ( .A0(n4), .A1(n308), .B0(n3), .Y(n294) );
  AOI21XL U246 ( .A0(n213), .A1(n308), .B0(n328), .Y(n216) );
  AOI21XL U247 ( .A0(n270), .A1(n353), .B0(n311), .Y(n183) );
  AOI21XL U248 ( .A0(n329), .A1(n226), .B0(n158), .Y(n159) );
  AOI21XL U249 ( .A0(n136), .A1(n352), .B0(n311), .Y(n137) );
  AOI21XL U250 ( .A0(n240), .A1(n249), .B0(n328), .Y(n85) );
  AOI21XL U251 ( .A0(n209), .A1(n320), .B0(n346), .Y(n74) );
  AOI21XL U252 ( .A0(n54), .A1(n53), .B0(n361), .Y(n61) );
  AOI21XL U253 ( .A0(n240), .A1(n82), .B0(n316), .Y(n51) );
  AOI21XL U254 ( .A0(n360), .A1(n290), .B0(n26), .Y(n27) );
  AOI21XL U255 ( .A0(n146), .A1(n353), .B0(n336), .Y(n18) );
  AOI21XL U256 ( .A0(n2), .A1(n251), .B0(n52), .Y(n14) );
  AOI21XL U257 ( .A0(n313), .A1(n200), .B0(n336), .Y(n52) );
  AOI21XL U258 ( .A0(n269), .A1(n268), .B0(n267), .Y(n280) );
  AOI21XL U259 ( .A0(n254), .A1(n3), .B0(n253), .Y(n262) );
  AOI21XL U260 ( .A0(n346), .A1(n347), .B0(n242), .Y(n243) );
  NOR2X1 U261 ( .A(n276), .B(n133), .Y(n348) );
  NOR2X1 U262 ( .A(n267), .B(n201), .Y(n351) );
  INVX1 U263 ( .A(a[7]), .Y(n267) );
  OAI21XL U264 ( .A0(n224), .A1(n341), .B0(n223), .Y(d[2]) );
  OAI21XL U265 ( .A0(n175), .A1(n361), .B0(n174), .Y(d[3]) );
  OAI21XL U266 ( .A0(n95), .A1(n361), .B0(n94), .Y(d[5]) );
  OAI21XL U267 ( .A0(n64), .A1(n299), .B0(n63), .Y(d[6]) );
  OAI21XL U268 ( .A0(n34), .A1(n361), .B0(n33), .Y(d[7]) );
  OAI21XL U269 ( .A0(n131), .A1(n299), .B0(n130), .Y(d[4]) );
  OAI21XL U270 ( .A0(n289), .A1(n321), .B0(n288), .Y(d[1]) );
  NAND2X1 U271 ( .A(a[7]), .B(a[5]), .Y(n133) );
  NOR2X1 U272 ( .A(n5), .B(n246), .Y(n214) );
  NAND2X1 U273 ( .A(a[4]), .B(n35), .Y(n269) );
  NOR2X1 U274 ( .A(a[4]), .B(n5), .Y(n273) );
  OAI21XL U275 ( .A0(n273), .A1(n229), .B0(n3), .Y(n7) );
  NOR2X1 U276 ( .A(a[7]), .B(a[2]), .Y(n340) );
  INVX1 U277 ( .A(n246), .Y(n252) );
  OAI21XL U278 ( .A0(n70), .A1(n340), .B0(n135), .Y(n6) );
  NAND3X1 U279 ( .A(n99), .B(n7), .C(n6), .Y(n12) );
  INVX1 U280 ( .A(n70), .Y(n115) );
  NOR2X1 U281 ( .A(n264), .B(n5), .Y(n325) );
  NAND3X1 U282 ( .A(n10), .B(n9), .C(n8), .Y(n11) );
  AOI211X1 U283 ( .A0(n329), .A1(n214), .B0(n12), .C0(n11), .Y(n34) );
  INVX1 U284 ( .A(a[6]), .Y(n20) );
  NOR2X1 U285 ( .A(a[0]), .B(n20), .Y(n129) );
  INVX1 U286 ( .A(n264), .Y(n309) );
  INVX1 U287 ( .A(n24), .Y(n327) );
  NAND2X1 U288 ( .A(n264), .B(n5), .Y(n349) );
  INVX1 U289 ( .A(n191), .Y(n200) );
  INVX1 U290 ( .A(n4), .Y(n336) );
  NAND2X1 U291 ( .A(n35), .B(n202), .Y(n107) );
  NAND2X1 U292 ( .A(n24), .B(n249), .Y(n266) );
  NAND4X1 U293 ( .A(n16), .B(n15), .C(n14), .D(n13), .Y(n32) );
  NAND2X1 U294 ( .A(a[3]), .B(n5), .Y(n270) );
  INVX1 U295 ( .A(n107), .Y(n41) );
  NOR2X1 U296 ( .A(n199), .B(n273), .Y(n165) );
  INVX1 U297 ( .A(n313), .Y(n271) );
  INVX1 U298 ( .A(n295), .Y(n213) );
  NOR2X1 U299 ( .A(a[1]), .B(n213), .Y(n228) );
  INVX1 U300 ( .A(n228), .Y(n239) );
  NAND2X1 U301 ( .A(n5), .B(n309), .Y(n144) );
  NOR2BX1 U302 ( .AN(n144), .B(n185), .Y(n96) );
  INVX1 U303 ( .A(n199), .Y(n146) );
  NAND2X1 U304 ( .A(a[0]), .B(n20), .Y(n299) );
  INVX1 U305 ( .A(n230), .Y(n256) );
  NAND2X1 U306 ( .A(n200), .B(n349), .Y(n121) );
  NAND2X1 U307 ( .A(n309), .B(n86), .Y(n290) );
  INVX1 U308 ( .A(n3), .Y(n303) );
  NAND2X1 U309 ( .A(n239), .B(n353), .Y(n105) );
  OAI21XL U310 ( .A0(n303), .A1(n105), .B0(n25), .Y(n26) );
  NOR2X1 U311 ( .A(a[6]), .B(a[0]), .Y(n93) );
  INVX1 U312 ( .A(n185), .Y(n113) );
  INVX1 U313 ( .A(n229), .Y(n304) );
  NAND2X1 U314 ( .A(n113), .B(n304), .Y(n104) );
  OAI21XL U315 ( .A0(n273), .A1(n164), .B0(n3), .Y(n36) );
  NAND4BXL U316 ( .AN(n250), .B(n38), .C(n37), .D(n36), .Y(n39) );
  NOR2X1 U317 ( .A(n145), .B(n332), .Y(n337) );
  INVX1 U318 ( .A(n273), .Y(n111) );
  INVX1 U319 ( .A(n308), .Y(n149) );
  NAND4X1 U320 ( .A(n48), .B(n47), .C(n46), .D(n45), .Y(n62) );
  INVX1 U321 ( .A(n214), .Y(n240) );
  INVX1 U322 ( .A(n332), .Y(n82) );
  INVX1 U323 ( .A(n329), .Y(n316) );
  OAI21XL U324 ( .A0(a[4]), .A1(n350), .B0(n49), .Y(n50) );
  NAND2X1 U325 ( .A(n313), .B(n256), .Y(n293) );
  NOR2X1 U326 ( .A(n355), .B(n293), .Y(n167) );
  OAI21XL U327 ( .A0(n325), .A1(n229), .B0(n298), .Y(n59) );
  OAI21XL U328 ( .A0(n120), .A1(n303), .B0(n55), .Y(n56) );
  NAND2X1 U329 ( .A(n270), .B(n312), .Y(n227) );
  INVX1 U330 ( .A(n190), .Y(n198) );
  NAND2X1 U331 ( .A(n3), .B(n313), .Y(n180) );
  NOR2X1 U332 ( .A(n350), .B(n313), .Y(n143) );
  NOR2X1 U333 ( .A(n278), .B(n276), .Y(n333) );
  OAI21XL U334 ( .A0(n353), .A1(n328), .B0(n75), .Y(n79) );
  INVX1 U335 ( .A(n76), .Y(n208) );
  OAI21XL U336 ( .A0(n225), .A1(n316), .B0(n77), .Y(n78) );
  NAND2X1 U337 ( .A(n346), .B(n213), .Y(n97) );
  INVX1 U338 ( .A(n129), .Y(n321) );
  NAND2X1 U339 ( .A(n111), .B(n270), .Y(n163) );
  OAI21XL U340 ( .A0(n120), .A1(n311), .B0(n83), .Y(n84) );
  NOR2X1 U341 ( .A(n149), .B(n320), .Y(n156) );
  NAND4X1 U342 ( .A(n100), .B(n99), .C(n98), .D(n97), .Y(n101) );
  AOI211X1 U343 ( .A0(n1), .A1(n156), .B0(n102), .C0(n101), .Y(n131) );
  OAI21XL U344 ( .A0(n252), .A1(n350), .B0(n180), .Y(n106) );
  NOR2X1 U345 ( .A(n107), .B(n5), .Y(n356) );
  OAI21XL U346 ( .A0(n190), .A1(n356), .B0(n329), .Y(n108) );
  NAND4BXL U347 ( .AN(n112), .B(n110), .C(n109), .D(n108), .Y(n128) );
  OAI21XL U348 ( .A0(n115), .A1(n197), .B0(n114), .Y(n116) );
  NAND2X1 U349 ( .A(n298), .B(n230), .Y(n247) );
  INVX1 U350 ( .A(n120), .Y(n207) );
  INVX1 U351 ( .A(n121), .Y(n192) );
  OAI21XL U352 ( .A0(n198), .A1(n238), .B0(n237), .Y(n122) );
  OAI21XL U353 ( .A0(a[1]), .A1(n136), .B0(n308), .Y(n132) );
  NOR2X1 U354 ( .A(n328), .B(n146), .Y(n358) );
  OAI21XL U355 ( .A0(n311), .A1(n304), .B0(n147), .Y(n148) );
  OAI21XL U356 ( .A0(n330), .A1(n149), .B0(n329), .Y(n150) );
  NAND4X1 U357 ( .A(n153), .B(n152), .C(n151), .D(n150), .Y(n173) );
  OAI21XL U358 ( .A0(n213), .A1(n255), .B0(n157), .Y(n158) );
  AOI211X1 U359 ( .A0(n287), .A1(n173), .B0(n172), .C0(n171), .Y(n174) );
  OAI21XL U360 ( .A0(n292), .A1(n276), .B0(n193), .Y(n194) );
  OAI21XL U361 ( .A0(n204), .A1(n208), .B0(n203), .Y(n205) );
  OAI21XL U362 ( .A0(n320), .A1(n356), .B0(n3), .Y(n217) );
  NOR2X1 U363 ( .A(n225), .B(n336), .Y(n236) );
  OAI21XL U364 ( .A0(n228), .A1(n273), .B0(n346), .Y(n232) );
  OAI21XL U365 ( .A0(n230), .A1(n229), .B0(n360), .Y(n231) );
  NAND4X1 U366 ( .A(n234), .B(n233), .C(n232), .D(n231), .Y(n235) );
  AOI211X1 U367 ( .A0(n337), .A1(n298), .B0(n236), .C0(n235), .Y(n289) );
  OAI21XL U368 ( .A0(n239), .A1(n238), .B0(n237), .Y(n245) );
  OAI21XL U369 ( .A0(n330), .A1(n316), .B0(n241), .Y(n242) );
  OAI21XL U370 ( .A0(n350), .A1(n347), .B0(n243), .Y(n244) );
  NOR2X1 U371 ( .A(n355), .B(n304), .Y(n314) );
  OAI21XL U372 ( .A0(n273), .A1(n272), .B0(n340), .Y(n274) );
  OAI21XL U373 ( .A0(n280), .A1(n279), .B0(n278), .Y(n281) );
  OAI21XL U374 ( .A0(n317), .A1(n316), .B0(n315), .Y(n318) );
  OAI21XL U375 ( .A0(n337), .A1(n336), .B0(n335), .Y(n338) );
  OAI21XL U376 ( .A0(n356), .A1(n355), .B0(n354), .Y(n357) );
endmodule


module aes_sbox_3 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368;

  INVX1 U1 ( .A(n99), .Y(n341) );
  OAI22X1 U2 ( .A0(n102), .A1(n237), .B0(n165), .B1(n303), .Y(n1) );
  AOI222X1 U3 ( .A0(n185), .A1(n10), .B0(n107), .B1(n298), .C0(n272), .C1(n329), .Y(n2) );
  NAND3X1 U4 ( .A(n103), .B(n104), .C(n2), .Y(n3) );
  AOI211X1 U5 ( .A0(n7), .A1(n156), .B0(n1), .C0(n3), .Y(n131) );
  NOR2X1 U6 ( .A(n196), .B(n105), .Y(n4) );
  AOI211X1 U7 ( .A0(n106), .A1(n10), .B0(n112), .C0(n4), .Y(n5) );
  OAI21XL U8 ( .A0(n190), .A1(n356), .B0(n329), .Y(n6) );
  NAND3X1 U9 ( .A(n110), .B(n5), .C(n6), .Y(n128) );
  NOR2BX1 U10 ( .AN(n349), .B(n311), .Y(n250) );
  AOI211XL U11 ( .A0(n287), .A1(n286), .B0(n285), .C0(n284), .Y(n288) );
  AOI31XL U12 ( .A0(n263), .A1(n262), .A2(n261), .B0(n341), .Y(n285) );
  AOI211X1 U13 ( .A0(n287), .A1(n222), .B0(n221), .C0(n220), .Y(n223) );
  NAND2XL U14 ( .A(n239), .B(n268), .Y(n339) );
  NOR2XL U15 ( .A(n328), .B(n146), .Y(n358) );
  NOR2X1 U16 ( .A(n199), .B(n273), .Y(n165) );
  INVX1 U17 ( .A(n325), .Y(n268) );
  NOR2X1 U18 ( .A(a[2]), .B(n278), .Y(n76) );
  CLKINVX3 U19 ( .A(a[5]), .Y(n278) );
  AOI31XL U20 ( .A0(n35), .A1(n34), .A2(n33), .B0(n341), .Y(n36) );
  AOI31XL U21 ( .A0(n125), .A1(n124), .A2(n123), .B0(n341), .Y(n126) );
  AOI211X1 U22 ( .A0(n7), .A1(n308), .B0(n183), .C0(n182), .Y(n224) );
  AOI21XL U23 ( .A0(n340), .A1(n339), .B0(n338), .Y(n342) );
  AOI2BB2XL U24 ( .B0(n360), .B1(n291), .A0N(n350), .A1N(n290), .Y(n302) );
  INVXL U25 ( .A(n260), .Y(n291) );
  NOR2XL U26 ( .A(n228), .B(n327), .Y(n260) );
  NAND2XL U27 ( .A(n113), .B(n88), .Y(n162) );
  INVXL U28 ( .A(n154), .Y(n312) );
  AOI32XL U29 ( .A0(n113), .A1(a[7]), .A2(n269), .B0(n163), .B1(n267), .Y(n197) );
  NAND2XL U30 ( .A(n313), .B(n240), .Y(n347) );
  NOR2X1 U31 ( .A(a[1]), .B(n295), .Y(n320) );
  NOR2XL U32 ( .A(n325), .B(n135), .Y(n265) );
  NOR2X1 U33 ( .A(n295), .B(n11), .Y(n154) );
  AOI2BB2XL U34 ( .B0(n360), .B1(n164), .A0N(n303), .A1N(n163), .Y(n169) );
  NAND2XL U35 ( .A(n144), .B(n30), .Y(n155) );
  NAND2XL U36 ( .A(a[1]), .B(n295), .Y(n92) );
  NAND2XL U37 ( .A(n198), .B(n277), .Y(n345) );
  INVX1 U38 ( .A(n298), .Y(n355) );
  CLKINVX3 U39 ( .A(n328), .Y(n8) );
  NAND2XL U40 ( .A(n330), .B(n11), .Y(n249) );
  NOR2XL U41 ( .A(n11), .B(n269), .Y(n191) );
  NOR2X1 U42 ( .A(a[1]), .B(n109), .Y(n332) );
  CLKINVX3 U43 ( .A(n269), .Y(n330) );
  NOR2XL U44 ( .A(a[1]), .B(n246), .Y(n190) );
  INVXL U45 ( .A(n270), .Y(n334) );
  NAND2X1 U46 ( .A(a[1]), .B(n41), .Y(n353) );
  NAND2X1 U47 ( .A(a[6]), .B(a[0]), .Y(n361) );
  INVX1 U48 ( .A(a[3]), .Y(n41) );
  AOI211XL U49 ( .A0(n129), .A1(n38), .B0(n37), .C0(n36), .Y(n39) );
  AOI211XL U50 ( .A0(n129), .A1(n128), .B0(n127), .C0(n126), .Y(n130) );
  AOI211XL U51 ( .A0(n129), .A1(n68), .B0(n67), .C0(n66), .Y(n69) );
  AOI31XL U52 ( .A0(n29), .A1(n28), .A2(n27), .B0(n299), .Y(n37) );
  OAI211XL U53 ( .A0(n249), .A1(n355), .B0(n248), .C0(n247), .Y(n286) );
  AOI211XL U54 ( .A0(n329), .A1(n260), .B0(n259), .C0(n258), .Y(n261) );
  OR4X2 U55 ( .A(n368), .B(n367), .C(n366), .D(n365), .Y(d[0]) );
  AOI211XL U56 ( .A0(n99), .A1(n98), .B0(n97), .C0(n96), .Y(n100) );
  AOI31XL U57 ( .A0(n95), .A1(n94), .A2(n93), .B0(n299), .Y(n96) );
  AOI31XL U58 ( .A0(n65), .A1(n64), .A2(n63), .B0(n341), .Y(n66) );
  AOI31XL U59 ( .A0(n212), .A1(n211), .A2(n210), .B0(n361), .Y(n221) );
  AOI211XL U60 ( .A0(n192), .A1(n10), .B0(n143), .C0(n142), .Y(n175) );
  OAI211XL U61 ( .A0(n197), .A1(n196), .B0(n195), .C0(n194), .Y(n222) );
  AOI31XL U62 ( .A0(n161), .A1(n160), .A2(n159), .B0(n321), .Y(n172) );
  AOI31XL U63 ( .A0(n170), .A1(n169), .A2(n168), .B0(n341), .Y(n171) );
  OAI22XL U64 ( .A0(n257), .A1(n350), .B0(n256), .B1(n255), .Y(n258) );
  AOI31XL U65 ( .A0(n246), .A1(n256), .A2(n245), .B0(n244), .Y(n248) );
  AOI22XL U66 ( .A0(n257), .A1(n298), .B0(n268), .B1(n108), .Y(n110) );
  AOI31XL U67 ( .A0(n344), .A1(n343), .A2(n342), .B0(n341), .Y(n366) );
  AOI31XL U68 ( .A0(n302), .A1(n301), .A2(n300), .B0(n299), .Y(n368) );
  OAI211XL U69 ( .A0(n80), .A1(n121), .B0(n79), .C0(n78), .Y(n98) );
  AOI211XL U70 ( .A0(n260), .A1(n360), .B0(n25), .C0(n24), .Y(n27) );
  OAI211XL U71 ( .A0(n350), .A1(n268), .B0(n141), .C0(n140), .Y(n142) );
  AOI211XL U72 ( .A0(n10), .A1(n339), .B0(n358), .C0(n148), .Y(n151) );
  AOI211XL U73 ( .A0(n329), .A1(n162), .B0(n91), .C0(n90), .Y(n94) );
  AOI211XL U74 ( .A0(a[7]), .A1(n339), .B0(n102), .C0(n115), .Y(n25) );
  AOI211XL U75 ( .A0(n298), .A1(n107), .B0(n46), .C0(n45), .Y(n70) );
  AOI211XL U76 ( .A0(n9), .A1(n92), .B0(n57), .C0(n56), .Y(n60) );
  AOI211XL U77 ( .A0(n326), .A1(n188), .B0(n58), .C0(n167), .Y(n59) );
  AOI211XL U78 ( .A0(n250), .A1(n240), .B0(n178), .C0(n62), .Y(n63) );
  AOI211XL U79 ( .A0(n8), .A1(n291), .B0(n167), .C0(n166), .Y(n168) );
  INVXL U80 ( .A(n107), .Y(n257) );
  AOI31XL U81 ( .A0(n118), .A1(n117), .A2(n247), .B0(n361), .Y(n127) );
  AOI211XL U82 ( .A0(n346), .A1(n268), .B0(n143), .C0(n119), .Y(n125) );
  AOI22XL U83 ( .A0(n8), .A1(n207), .B0(n192), .B1(n122), .Y(n123) );
  AOI21X1 U84 ( .A0(n360), .A1(n227), .B0(n75), .Y(n101) );
  AOI211XL U85 ( .A0(n329), .A1(n198), .B0(n77), .C0(n143), .Y(n78) );
  AOI31XL U86 ( .A0(n87), .A1(n86), .A2(n103), .B0(n321), .Y(n97) );
  AOI31XL U87 ( .A0(n324), .A1(n323), .A2(n322), .B0(n321), .Y(n367) );
  AOI31XL U88 ( .A0(n364), .A1(n363), .A2(n362), .B0(n361), .Y(n365) );
  AOI211XL U89 ( .A0(n7), .A1(n207), .B0(n206), .C0(n205), .Y(n211) );
  AOI211XL U90 ( .A0(n189), .A1(n188), .B0(n187), .C0(n186), .Y(n195) );
  AOI31XL U91 ( .A0(n219), .A1(n218), .A2(n217), .B0(n321), .Y(n220) );
  OAI211XL U92 ( .A0(n337), .A1(n237), .B0(n181), .C0(n180), .Y(n182) );
  AOI31XL U93 ( .A0(n283), .A1(n282), .A2(n281), .B0(n361), .Y(n284) );
  AOI22XL U94 ( .A0(n8), .A1(n227), .B0(n9), .B1(n226), .Y(n234) );
  AOI211XL U95 ( .A0(n360), .A1(n359), .B0(n358), .C0(n357), .Y(n362) );
  AOI211XL U96 ( .A0(n329), .A1(n266), .B0(n216), .C0(n215), .Y(n218) );
  AOI221XL U97 ( .A0(n346), .A1(n330), .B0(n9), .B1(n269), .C0(n116), .Y(n117)
         );
  AOI211XL U98 ( .A0(n320), .A1(n7), .B0(n319), .C0(n318), .Y(n322) );
  AOI211XL U99 ( .A0(n350), .A1(n303), .B0(n185), .C0(n264), .Y(n186) );
  AOI211XL U100 ( .A0(n8), .A1(n139), .B0(n138), .C0(n137), .Y(n140) );
  AOI211XL U101 ( .A0(n298), .A1(n179), .B0(n178), .C0(n177), .Y(n181) );
  AOI2BB2XL U102 ( .B0(n264), .B1(n360), .A0N(n350), .A1N(n265), .Y(n283) );
  AOI211XL U103 ( .A0(n10), .A1(n251), .B0(n250), .C0(n314), .Y(n263) );
  AOI211XL U104 ( .A0(n298), .A1(n290), .B0(n85), .C0(n84), .Y(n86) );
  OAI211XL U105 ( .A0(n252), .A1(n336), .B0(n74), .C0(n73), .Y(n75) );
  AOI2BB2XL U106 ( .B0(n10), .B1(n337), .A0N(n350), .A1N(n179), .Y(n54) );
  NAND2XL U107 ( .A(n239), .B(n277), .Y(n188) );
  AOI22XL U108 ( .A0(n7), .A1(n230), .B0(n252), .B1(n329), .Y(n233) );
  NOR3XL U109 ( .A(n325), .B(n252), .C(n328), .Y(n253) );
  AOI22XL U110 ( .A0(n9), .A1(n192), .B0(n360), .B1(n154), .Y(n161) );
  AOI211XL U111 ( .A0(a[2]), .A1(n134), .B0(n317), .C0(n133), .Y(n138) );
  OAI22XL U112 ( .A0(n356), .A1(n354), .B0(n176), .B1(n184), .Y(n177) );
  AOI22XL U113 ( .A0(n192), .A1(n276), .B0(n237), .B1(n316), .Y(n193) );
  AOI22XL U114 ( .A0(a[1]), .A1(n10), .B0(n7), .B1(n334), .Y(n219) );
  AOI22XL U115 ( .A0(a[3]), .A1(n10), .B0(n7), .B1(n349), .Y(n363) );
  AOI31XL U116 ( .A0(n8), .A1(n353), .A2(n352), .B0(n310), .Y(n323) );
  AOI211XL U117 ( .A0(n298), .A1(n352), .B0(n297), .C0(n296), .Y(n300) );
  AOI2BB2XL U118 ( .B0(n8), .B1(n293), .A0N(n316), .A1N(n292), .Y(n301) );
  AOI22XL U119 ( .A0(n9), .A1(n50), .B0(n346), .B1(n290), .Y(n51) );
  AOI22XL U120 ( .A0(n228), .A1(n329), .B0(n298), .B1(n105), .Y(n53) );
  AOI22XL U121 ( .A0(n7), .A1(n106), .B0(n326), .B1(n176), .Y(n44) );
  OAI22XL U122 ( .A0(n41), .A1(n328), .B0(n201), .B1(n155), .Y(n46) );
  AOI22XL U123 ( .A0(n7), .A1(n293), .B0(n259), .B1(n268), .Y(n89) );
  AOI22XL U124 ( .A0(n102), .A1(n7), .B0(n10), .B1(n305), .Y(n87) );
  AOI22XL U125 ( .A0(n7), .A1(n307), .B0(n10), .B1(n48), .Y(n35) );
  AOI22XL U126 ( .A0(n165), .A1(n8), .B0(n23), .B1(n268), .Y(n28) );
  AOI22XL U127 ( .A0(n9), .A1(n134), .B0(n360), .B1(n266), .Y(n19) );
  NAND2XL U128 ( .A(n268), .B(n349), .Y(n251) );
  AOI22XL U129 ( .A0(n7), .A1(n295), .B0(n298), .B1(n327), .Y(n21) );
  AOI22XL U130 ( .A0(n7), .A1(n30), .B0(n346), .B1(n320), .Y(n15) );
  AOI2BB2XL U131 ( .B0(n10), .B1(n92), .A0N(n237), .A1N(n106), .Y(n61) );
  NOR2XL U132 ( .A(n228), .B(n154), .Y(n120) );
  NOR2XL U133 ( .A(n185), .B(n104), .Y(n178) );
  AOI22XL U134 ( .A0(n7), .A1(n214), .B0(n329), .B1(n268), .Y(n64) );
  AOI22XL U135 ( .A0(n330), .A1(n9), .B0(n298), .B1(n139), .Y(n74) );
  INVXL U136 ( .A(n156), .Y(n226) );
  AOI22XL U137 ( .A0(n7), .A1(n290), .B0(n346), .B1(n269), .Y(n157) );
  AOI22XL U138 ( .A0(n10), .A1(n162), .B0(n329), .B1(n179), .Y(n170) );
  NAND3XL U139 ( .A(n9), .B(n144), .C(n92), .Y(n93) );
  NOR2XL U140 ( .A(n213), .B(n237), .Y(n259) );
  AOI22XL U141 ( .A0(n298), .A1(n146), .B0(n10), .B1(n163), .Y(n95) );
  AOI22XL U142 ( .A0(n76), .A1(n154), .B0(n10), .B1(n266), .Y(n79) );
  AOI211XL U143 ( .A0(n8), .A1(n271), .B0(n72), .C0(n297), .Y(n73) );
  NAND2XL U144 ( .A(n113), .B(n246), .Y(n139) );
  AOI22XL U145 ( .A0(n9), .A1(n49), .B0(n346), .B1(n71), .Y(n29) );
  NOR2XL U146 ( .A(n154), .B(n332), .Y(n134) );
  AOI22XL U147 ( .A0(n298), .A1(n154), .B0(n10), .B1(n265), .Y(n14) );
  NAND2XL U148 ( .A(n8), .B(n269), .Y(n104) );
  AOI22XL U149 ( .A0(n8), .A1(n102), .B0(n346), .B1(n11), .Y(n55) );
  AOI22XL U150 ( .A0(n8), .A1(n49), .B0(n360), .B1(n48), .Y(n52) );
  INVXL U151 ( .A(n92), .Y(n176) );
  AOI22XL U152 ( .A0(a[3]), .A1(n346), .B0(n8), .B1(n202), .Y(n204) );
  AOI22XL U153 ( .A0(n199), .A1(n333), .B0(n329), .B1(n345), .Y(n212) );
  INVXL U154 ( .A(n184), .Y(n187) );
  OAI211XL U155 ( .A0(n277), .A1(n276), .B0(n275), .C0(n274), .Y(n279) );
  AOI22XL U156 ( .A0(n9), .A1(n266), .B0(n329), .B1(n265), .Y(n282) );
  AOI22XL U157 ( .A0(n8), .A1(n292), .B0(n334), .B1(n10), .Y(n241) );
  NAND2XL U158 ( .A(n353), .B(n352), .Y(n359) );
  AOI22XL U159 ( .A0(n9), .A1(n347), .B0(n346), .B1(n345), .Y(n364) );
  AOI22XL U160 ( .A0(n330), .A1(n329), .B0(n8), .B1(n327), .Y(n343) );
  INVXL U161 ( .A(n314), .Y(n315) );
  NOR2XL U162 ( .A(n295), .B(n294), .Y(n296) );
  AOI22XL U163 ( .A0(n9), .A1(n230), .B0(n10), .B1(n225), .Y(n203) );
  AOI22XL U164 ( .A0(n189), .A1(n320), .B0(n8), .B1(n265), .Y(n114) );
  NOR2XL U165 ( .A(n165), .B(n311), .Y(n166) );
  AOI22XL U166 ( .A0(n271), .A1(n10), .B0(n8), .B1(n155), .Y(n160) );
  OAI2BB1XL U167 ( .A0N(n214), .A1N(n326), .B0(n247), .Y(n215) );
  NAND2XL U168 ( .A(n109), .B(n256), .Y(n307) );
  AOI22XL U169 ( .A0(n8), .A1(n121), .B0(n329), .B1(n155), .Y(n34) );
  NAND2XL U170 ( .A(n313), .B(n200), .Y(n50) );
  NAND2XL U171 ( .A(n10), .B(n249), .Y(n184) );
  AOI22XL U172 ( .A0(n230), .A1(n209), .B0(n360), .B1(n313), .Y(n16) );
  AOI22XL U173 ( .A0(n10), .A1(n353), .B0(n112), .B1(n111), .Y(n118) );
  AND2X2 U174 ( .A(n305), .B(n88), .Y(n225) );
  AOI31XL U175 ( .A0(n355), .A1(n237), .A2(n180), .B0(n330), .Y(n77) );
  AOI22XL U176 ( .A0(n298), .A1(n132), .B0(n360), .B1(n308), .Y(n141) );
  NOR2XL U177 ( .A(n185), .B(n272), .Y(n317) );
  INVXL U178 ( .A(n135), .Y(n352) );
  AOI22XL U179 ( .A0(n271), .A1(n360), .B0(n340), .B1(n332), .Y(n147) );
  NOR3XL U180 ( .A(n185), .B(n264), .C(n311), .Y(n297) );
  AOI22XL U181 ( .A0(a[1]), .A1(n298), .B0(n9), .B1(n144), .Y(n153) );
  AOI211XL U182 ( .A0(a[7]), .A1(n71), .B0(n191), .C0(n115), .Y(n72) );
  NOR2XL U183 ( .A(n47), .B(n149), .Y(n105) );
  OAI22XL U184 ( .A0(n327), .A1(n237), .B0(n201), .B1(n200), .Y(n206) );
  OAI22XL U185 ( .A0(n355), .A1(n198), .B0(n308), .B1(n316), .Y(n119) );
  AOI22XL U186 ( .A0(n230), .A1(n10), .B0(n340), .B1(n356), .Y(n124) );
  AOI22XL U187 ( .A0(n190), .A1(n360), .B0(n329), .B1(n109), .Y(n43) );
  NOR2XL U188 ( .A(n271), .B(n355), .Y(n23) );
  NOR2XL U189 ( .A(n295), .B(n230), .Y(n49) );
  AOI22XL U190 ( .A0(a[4]), .A1(n298), .B0(n346), .B1(n308), .Y(n31) );
  NAND3XL U191 ( .A(n209), .B(n246), .C(n208), .Y(n210) );
  AOI22XL U192 ( .A0(n334), .A1(n333), .B0(n332), .B1(n331), .Y(n335) );
  NAND3XL U193 ( .A(n9), .B(a[3]), .C(n208), .Y(n83) );
  NOR2XL U194 ( .A(n191), .B(n190), .Y(n292) );
  NOR2XL U195 ( .A(a[1]), .B(n330), .Y(n272) );
  AOI22XL U196 ( .A0(n145), .A1(n333), .B0(n254), .B1(n331), .Y(n152) );
  AOI22XL U197 ( .A0(n326), .A1(n325), .B0(n9), .B1(n11), .Y(n344) );
  NOR2XL U198 ( .A(n237), .B(n332), .Y(n112) );
  NAND2XL U199 ( .A(n308), .B(n270), .Y(n71) );
  AOI22XL U200 ( .A0(n191), .A1(n209), .B0(n329), .B1(n309), .Y(n22) );
  NOR2XL U201 ( .A(a[1]), .B(n252), .Y(n135) );
  NAND2XL U202 ( .A(n313), .B(n305), .Y(n48) );
  OR2X2 U203 ( .A(a[7]), .B(n115), .Y(n350) );
  NOR2XL U204 ( .A(n47), .B(a[1]), .Y(n199) );
  NAND2XL U205 ( .A(n111), .B(n349), .Y(n179) );
  AOI22XL U206 ( .A0(n271), .A1(n326), .B0(n331), .B1(n270), .Y(n275) );
  NAND3XL U207 ( .A(n333), .B(n82), .C(n246), .Y(n81) );
  INVXL U208 ( .A(n333), .Y(n238) );
  NAND2XL U209 ( .A(n329), .B(n313), .Y(n354) );
  INVXL U210 ( .A(n299), .Y(n287) );
  INVXL U211 ( .A(n201), .Y(n189) );
  INVXL U212 ( .A(n196), .Y(n209) );
  NAND2XL U213 ( .A(a[1]), .B(n264), .Y(n305) );
  OR2X2 U214 ( .A(n267), .B(n196), .Y(n328) );
  NAND2XL U215 ( .A(a[2]), .B(n278), .Y(n196) );
  NOR2XL U216 ( .A(a[1]), .B(n202), .Y(n164) );
  AOI22XL U217 ( .A0(a[1]), .A1(a[7]), .B0(n267), .B1(n11), .Y(n82) );
  NAND2XL U218 ( .A(n267), .B(n278), .Y(n255) );
  NOR2XL U219 ( .A(n267), .B(n276), .Y(n331) );
  INVXL U220 ( .A(n277), .Y(n254) );
  AOI22XL U221 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n276), .Y(n136) );
  NOR2XL U222 ( .A(a[3]), .B(a[1]), .Y(n229) );
  NAND2XL U223 ( .A(a[4]), .B(a[1]), .Y(n277) );
  INVX2 U224 ( .A(a[2]), .Y(n276) );
  INVX2 U225 ( .A(a[4]), .Y(n202) );
  NAND2XL U226 ( .A(a[3]), .B(a[1]), .Y(n30) );
  NAND2X2 U227 ( .A(n278), .B(n276), .Y(n201) );
  NOR2X2 U228 ( .A(n41), .B(n202), .Y(n264) );
  NOR2X2 U229 ( .A(n47), .B(n11), .Y(n185) );
  NAND2X2 U230 ( .A(a[1]), .B(n246), .Y(n308) );
  NAND2X2 U231 ( .A(a[3]), .B(n202), .Y(n246) );
  NOR2X2 U232 ( .A(n276), .B(a[7]), .Y(n326) );
  NOR2X2 U233 ( .A(n252), .B(n330), .Y(n295) );
  NOR2X2 U234 ( .A(n330), .B(n11), .Y(n230) );
  NAND2X2 U235 ( .A(n202), .B(n11), .Y(n313) );
  CLKINVX3 U236 ( .A(n237), .Y(n360) );
  NAND2X2 U237 ( .A(a[5]), .B(n326), .Y(n237) );
  CLKINVX3 U238 ( .A(n350), .Y(n7) );
  NOR2X4 U239 ( .A(a[2]), .B(n133), .Y(n329) );
  BUFX3 U240 ( .A(n348), .Y(n9) );
  NOR2X4 U241 ( .A(a[7]), .B(n201), .Y(n298) );
  CLKINVX3 U242 ( .A(a[1]), .Y(n11) );
  CLKINVX3 U243 ( .A(n311), .Y(n346) );
  NAND2X2 U244 ( .A(n278), .B(n326), .Y(n311) );
  BUFX3 U245 ( .A(n351), .Y(n10) );
  AOI21XL U246 ( .A0(n313), .A1(n312), .B0(n311), .Y(n319) );
  AOI21XL U247 ( .A0(n309), .A1(n308), .B0(n336), .Y(n310) );
  AOI21XL U248 ( .A0(n360), .A1(n307), .B0(n306), .Y(n324) );
  AOI21XL U249 ( .A0(n305), .A1(n304), .B0(n303), .Y(n306) );
  AOI21XL U250 ( .A0(n10), .A1(n308), .B0(n9), .Y(n294) );
  AOI21XL U251 ( .A0(n213), .A1(n308), .B0(n328), .Y(n216) );
  AOI21XL U252 ( .A0(n270), .A1(n353), .B0(n311), .Y(n183) );
  AOI21XL U253 ( .A0(n329), .A1(n226), .B0(n158), .Y(n159) );
  AOI21XL U254 ( .A0(n136), .A1(n352), .B0(n311), .Y(n137) );
  AOI21XL U255 ( .A0(n240), .A1(n249), .B0(n328), .Y(n91) );
  AOI21XL U256 ( .A0(n209), .A1(n320), .B0(n346), .Y(n80) );
  AOI21XL U257 ( .A0(n60), .A1(n59), .B0(n361), .Y(n67) );
  AOI21XL U258 ( .A0(n240), .A1(n88), .B0(n316), .Y(n57) );
  AOI21XL U259 ( .A0(n360), .A1(n290), .B0(n32), .Y(n33) );
  AOI21XL U260 ( .A0(n146), .A1(n353), .B0(n336), .Y(n24) );
  AOI21XL U261 ( .A0(n8), .A1(n251), .B0(n58), .Y(n20) );
  AOI21XL U262 ( .A0(n313), .A1(n200), .B0(n336), .Y(n58) );
  AOI21XL U263 ( .A0(n269), .A1(n268), .B0(n267), .Y(n280) );
  AOI21XL U264 ( .A0(n254), .A1(n9), .B0(n253), .Y(n262) );
  AOI21XL U265 ( .A0(n346), .A1(n347), .B0(n242), .Y(n243) );
  NOR2X1 U266 ( .A(n276), .B(n133), .Y(n348) );
  NOR2X1 U267 ( .A(n267), .B(n201), .Y(n351) );
  INVX1 U268 ( .A(a[7]), .Y(n267) );
  OAI21XL U269 ( .A0(n224), .A1(n341), .B0(n223), .Y(d[2]) );
  OAI21XL U270 ( .A0(n175), .A1(n361), .B0(n174), .Y(d[3]) );
  OAI21XL U271 ( .A0(n101), .A1(n361), .B0(n100), .Y(d[5]) );
  OAI21XL U272 ( .A0(n70), .A1(n299), .B0(n69), .Y(d[6]) );
  OAI21XL U273 ( .A0(n40), .A1(n361), .B0(n39), .Y(d[7]) );
  OAI21XL U274 ( .A0(n131), .A1(n299), .B0(n130), .Y(d[4]) );
  OAI21XL U275 ( .A0(n289), .A1(n321), .B0(n288), .Y(d[1]) );
  NAND2X1 U276 ( .A(a[7]), .B(a[5]), .Y(n133) );
  NOR2X1 U277 ( .A(n11), .B(n246), .Y(n214) );
  NAND2X1 U278 ( .A(a[4]), .B(n41), .Y(n269) );
  NOR2X1 U279 ( .A(a[4]), .B(n11), .Y(n273) );
  OAI21XL U280 ( .A0(n273), .A1(n229), .B0(n9), .Y(n13) );
  NOR2X1 U281 ( .A(a[7]), .B(a[2]), .Y(n340) );
  INVX1 U282 ( .A(n246), .Y(n252) );
  OAI21XL U283 ( .A0(n76), .A1(n340), .B0(n135), .Y(n12) );
  NAND3X1 U284 ( .A(n104), .B(n13), .C(n12), .Y(n18) );
  INVX1 U285 ( .A(n76), .Y(n115) );
  NOR2X1 U286 ( .A(n264), .B(n11), .Y(n325) );
  NAND3X1 U287 ( .A(n16), .B(n15), .C(n14), .Y(n17) );
  AOI211X1 U288 ( .A0(n329), .A1(n214), .B0(n18), .C0(n17), .Y(n40) );
  INVX1 U289 ( .A(a[6]), .Y(n26) );
  NOR2X1 U290 ( .A(a[0]), .B(n26), .Y(n129) );
  INVX1 U291 ( .A(n264), .Y(n309) );
  INVX1 U292 ( .A(n30), .Y(n327) );
  NAND2X1 U293 ( .A(n264), .B(n11), .Y(n349) );
  INVX1 U294 ( .A(n191), .Y(n200) );
  INVX1 U295 ( .A(n10), .Y(n336) );
  NAND2X1 U296 ( .A(n41), .B(n202), .Y(n109) );
  NAND2X1 U297 ( .A(n30), .B(n249), .Y(n266) );
  NAND4X1 U298 ( .A(n22), .B(n21), .C(n20), .D(n19), .Y(n38) );
  NAND2X1 U299 ( .A(a[3]), .B(n11), .Y(n270) );
  INVX1 U300 ( .A(n109), .Y(n47) );
  INVX1 U301 ( .A(n313), .Y(n271) );
  INVX1 U302 ( .A(n295), .Y(n213) );
  NOR2X1 U303 ( .A(a[1]), .B(n213), .Y(n228) );
  INVX1 U304 ( .A(n228), .Y(n239) );
  NAND2X1 U305 ( .A(n11), .B(n309), .Y(n144) );
  NOR2BX1 U306 ( .AN(n144), .B(n185), .Y(n102) );
  INVX1 U307 ( .A(n199), .Y(n146) );
  NAND2X1 U308 ( .A(a[0]), .B(n26), .Y(n299) );
  INVX1 U309 ( .A(n230), .Y(n256) );
  NAND2X1 U310 ( .A(n200), .B(n349), .Y(n121) );
  NAND2X1 U311 ( .A(n309), .B(n92), .Y(n290) );
  INVX1 U312 ( .A(n9), .Y(n303) );
  NAND2X1 U313 ( .A(n239), .B(n353), .Y(n107) );
  OAI21XL U314 ( .A0(n303), .A1(n107), .B0(n31), .Y(n32) );
  NOR2X1 U315 ( .A(a[6]), .B(a[0]), .Y(n99) );
  INVX1 U316 ( .A(n185), .Y(n113) );
  INVX1 U317 ( .A(n229), .Y(n304) );
  NAND2X1 U318 ( .A(n113), .B(n304), .Y(n106) );
  OAI21XL U319 ( .A0(n273), .A1(n164), .B0(n9), .Y(n42) );
  NAND4BXL U320 ( .AN(n250), .B(n44), .C(n43), .D(n42), .Y(n45) );
  INVX1 U321 ( .A(n353), .Y(n145) );
  NOR2X1 U322 ( .A(n145), .B(n332), .Y(n337) );
  INVX1 U323 ( .A(n273), .Y(n111) );
  INVX1 U324 ( .A(n308), .Y(n149) );
  NAND4X1 U325 ( .A(n54), .B(n53), .C(n52), .D(n51), .Y(n68) );
  INVX1 U326 ( .A(n214), .Y(n240) );
  INVX1 U327 ( .A(n332), .Y(n88) );
  INVX1 U328 ( .A(n329), .Y(n316) );
  OAI21XL U329 ( .A0(a[4]), .A1(n350), .B0(n55), .Y(n56) );
  NAND2X1 U330 ( .A(n313), .B(n256), .Y(n293) );
  NOR2X1 U331 ( .A(n355), .B(n293), .Y(n167) );
  OAI21XL U332 ( .A0(n325), .A1(n229), .B0(n298), .Y(n65) );
  OAI21XL U333 ( .A0(n120), .A1(n303), .B0(n61), .Y(n62) );
  NAND2X1 U334 ( .A(n270), .B(n312), .Y(n227) );
  INVX1 U335 ( .A(n190), .Y(n198) );
  NAND2X1 U336 ( .A(n9), .B(n313), .Y(n180) );
  NOR2X1 U337 ( .A(n350), .B(n313), .Y(n143) );
  NOR2X1 U338 ( .A(n278), .B(n276), .Y(n333) );
  OAI21XL U339 ( .A0(n353), .A1(n328), .B0(n81), .Y(n85) );
  INVX1 U340 ( .A(n82), .Y(n208) );
  OAI21XL U341 ( .A0(n225), .A1(n316), .B0(n83), .Y(n84) );
  NAND2X1 U342 ( .A(n346), .B(n213), .Y(n103) );
  INVX1 U343 ( .A(n129), .Y(n321) );
  NAND2X1 U344 ( .A(n111), .B(n270), .Y(n163) );
  OAI21XL U345 ( .A0(n120), .A1(n311), .B0(n89), .Y(n90) );
  NOR2X1 U346 ( .A(n149), .B(n320), .Y(n156) );
  OAI21XL U347 ( .A0(n252), .A1(n350), .B0(n180), .Y(n108) );
  NOR2X1 U348 ( .A(n109), .B(n11), .Y(n356) );
  OAI21XL U349 ( .A0(n115), .A1(n197), .B0(n114), .Y(n116) );
  NAND2X1 U350 ( .A(n298), .B(n230), .Y(n247) );
  INVX1 U351 ( .A(n120), .Y(n207) );
  INVX1 U352 ( .A(n121), .Y(n192) );
  OAI21XL U353 ( .A0(n198), .A1(n238), .B0(n237), .Y(n122) );
  OAI21XL U354 ( .A0(a[1]), .A1(n136), .B0(n308), .Y(n132) );
  OAI21XL U355 ( .A0(n311), .A1(n304), .B0(n147), .Y(n148) );
  OAI21XL U356 ( .A0(n330), .A1(n149), .B0(n329), .Y(n150) );
  NAND4X1 U357 ( .A(n153), .B(n152), .C(n151), .D(n150), .Y(n173) );
  OAI21XL U358 ( .A0(n213), .A1(n255), .B0(n157), .Y(n158) );
  AOI211X1 U359 ( .A0(n287), .A1(n173), .B0(n172), .C0(n171), .Y(n174) );
  OAI21XL U360 ( .A0(n292), .A1(n276), .B0(n193), .Y(n194) );
  OAI21XL U361 ( .A0(n204), .A1(n208), .B0(n203), .Y(n205) );
  OAI21XL U362 ( .A0(n320), .A1(n356), .B0(n9), .Y(n217) );
  NOR2X1 U363 ( .A(n225), .B(n336), .Y(n236) );
  OAI21XL U364 ( .A0(n228), .A1(n273), .B0(n346), .Y(n232) );
  OAI21XL U365 ( .A0(n230), .A1(n229), .B0(n360), .Y(n231) );
  NAND4X1 U366 ( .A(n234), .B(n233), .C(n232), .D(n231), .Y(n235) );
  AOI211X1 U367 ( .A0(n337), .A1(n298), .B0(n236), .C0(n235), .Y(n289) );
  OAI21XL U368 ( .A0(n239), .A1(n238), .B0(n237), .Y(n245) );
  OAI21XL U369 ( .A0(n330), .A1(n316), .B0(n241), .Y(n242) );
  OAI21XL U370 ( .A0(n350), .A1(n347), .B0(n243), .Y(n244) );
  NOR2X1 U371 ( .A(n355), .B(n304), .Y(n314) );
  OAI21XL U372 ( .A0(n273), .A1(n272), .B0(n340), .Y(n274) );
  OAI21XL U373 ( .A0(n280), .A1(n279), .B0(n278), .Y(n281) );
  OAI21XL U374 ( .A0(n317), .A1(n316), .B0(n315), .Y(n318) );
  OAI21XL U375 ( .A0(n337), .A1(n336), .B0(n335), .Y(n338) );
  OAI21XL U376 ( .A0(n356), .A1(n355), .B0(n354), .Y(n357) );
endmodule


module aes_key_expand_128 ( clk, kld, key, wo_0, wo_1, wo_2, wo_3 );
  input [127:0] key;
  output [31:0] wo_0;
  output [31:0] wo_1;
  output [31:0] wo_2;
  output [31:0] wo_3;
  input clk, kld;
  wire   N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, n1, n2, n3, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n29, n30, n31, n32, n33, n34, n35, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n61, n62, n63, n64, n65, n66, n67,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96, n97,
         n98, n99, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n125, n126, n127, n128, n258, n259, n260, n261, n262,
         n263, n264, n265, n4, n28, n36, n60, n68, n92, n100, n124, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311;
  wire   [31:0] subword;
  wire   [31:0] rcon;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23;

  aes_sbox_3 u0 ( .a(wo_3[23:16]), .d(subword[31:24]) );
  aes_sbox_2 u1 ( .a(wo_3[15:8]), .d(subword[23:16]) );
  aes_sbox_1 u2 ( .a(wo_3[7:0]), .d(subword[15:8]) );
  aes_sbox_0 u3 ( .a(wo_3[31:24]), .d(subword[7:0]) );
  aes_rcon r0 ( .clk(clk), .kld(kld), .out({rcon[31:24], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23}) );
  DFFHQX1 \w_reg[2][0]  ( .D(n127), .CK(clk), .Q(wo_2[0]) );
  DFFHQX1 \w_reg[2][1]  ( .D(n123), .CK(clk), .Q(wo_2[1]) );
  DFFHQX1 \w_reg[2][2]  ( .D(n119), .CK(clk), .Q(wo_2[2]) );
  DFFHQX1 \w_reg[2][3]  ( .D(n115), .CK(clk), .Q(wo_2[3]) );
  DFFHQX1 \w_reg[2][8]  ( .D(n95), .CK(clk), .Q(wo_2[8]) );
  DFFHQX1 \w_reg[1][8]  ( .D(n94), .CK(clk), .Q(wo_1[8]) );
  DFFHQX1 \w_reg[2][9]  ( .D(n91), .CK(clk), .Q(wo_2[9]) );
  DFFHQX1 \w_reg[1][9]  ( .D(n90), .CK(clk), .Q(wo_1[9]) );
  DFFHQX1 \w_reg[2][10]  ( .D(n87), .CK(clk), .Q(wo_2[10]) );
  DFFHQX1 \w_reg[1][10]  ( .D(n86), .CK(clk), .Q(wo_1[10]) );
  DFFHQX1 \w_reg[2][11]  ( .D(n83), .CK(clk), .Q(wo_2[11]) );
  DFFHQX1 \w_reg[1][11]  ( .D(n82), .CK(clk), .Q(wo_1[11]) );
  DFFHQX1 \w_reg[2][12]  ( .D(n79), .CK(clk), .Q(wo_2[12]) );
  DFFHQX1 \w_reg[1][12]  ( .D(n78), .CK(clk), .Q(wo_1[12]) );
  DFFHQX1 \w_reg[2][13]  ( .D(n75), .CK(clk), .Q(wo_2[13]) );
  DFFHQX1 \w_reg[1][13]  ( .D(n74), .CK(clk), .Q(wo_1[13]) );
  DFFHQX1 \w_reg[2][14]  ( .D(n71), .CK(clk), .Q(wo_2[14]) );
  DFFHQX1 \w_reg[1][14]  ( .D(n70), .CK(clk), .Q(wo_1[14]) );
  DFFHQX1 \w_reg[2][16]  ( .D(n63), .CK(clk), .Q(wo_2[16]) );
  DFFHQX1 \w_reg[1][16]  ( .D(n62), .CK(clk), .Q(wo_1[16]) );
  DFFHQX1 \w_reg[2][17]  ( .D(n59), .CK(clk), .Q(wo_2[17]) );
  DFFHQX1 \w_reg[1][17]  ( .D(n58), .CK(clk), .Q(wo_1[17]) );
  DFFHQX1 \w_reg[2][18]  ( .D(n55), .CK(clk), .Q(wo_2[18]) );
  DFFHQX1 \w_reg[1][18]  ( .D(n54), .CK(clk), .Q(wo_1[18]) );
  DFFHQX1 \w_reg[2][19]  ( .D(n51), .CK(clk), .Q(wo_2[19]) );
  DFFHQX1 \w_reg[1][19]  ( .D(n50), .CK(clk), .Q(wo_1[19]) );
  DFFHQX1 \w_reg[2][20]  ( .D(n47), .CK(clk), .Q(wo_2[20]) );
  DFFHQX1 \w_reg[1][20]  ( .D(n46), .CK(clk), .Q(wo_1[20]) );
  DFFHQX1 \w_reg[2][21]  ( .D(n43), .CK(clk), .Q(wo_2[21]) );
  DFFHQX1 \w_reg[1][21]  ( .D(n42), .CK(clk), .Q(wo_1[21]) );
  DFFHQX1 \w_reg[2][22]  ( .D(n39), .CK(clk), .Q(wo_2[22]) );
  DFFHQX1 \w_reg[1][22]  ( .D(n38), .CK(clk), .Q(wo_1[22]) );
  DFFHQX1 \w_reg[2][24]  ( .D(n31), .CK(clk), .Q(wo_2[24]) );
  DFFHQX1 \w_reg[1][24]  ( .D(n30), .CK(clk), .Q(wo_1[24]) );
  DFFHQX1 \w_reg[2][25]  ( .D(n27), .CK(clk), .Q(wo_2[25]) );
  DFFHQX1 \w_reg[1][25]  ( .D(n26), .CK(clk), .Q(wo_1[25]) );
  DFFHQX1 \w_reg[2][26]  ( .D(n23), .CK(clk), .Q(wo_2[26]) );
  DFFHQX1 \w_reg[1][26]  ( .D(n22), .CK(clk), .Q(wo_1[26]) );
  DFFHQX1 \w_reg[2][27]  ( .D(n19), .CK(clk), .Q(wo_2[27]) );
  DFFHQX1 \w_reg[1][27]  ( .D(n18), .CK(clk), .Q(wo_1[27]) );
  DFFHQX1 \w_reg[2][28]  ( .D(n15), .CK(clk), .Q(wo_2[28]) );
  DFFHQX1 \w_reg[1][28]  ( .D(n14), .CK(clk), .Q(wo_1[28]) );
  DFFHQX1 \w_reg[2][29]  ( .D(n11), .CK(clk), .Q(wo_2[29]) );
  DFFHQX1 \w_reg[1][29]  ( .D(n10), .CK(clk), .Q(wo_1[29]) );
  DFFHQX1 \w_reg[2][30]  ( .D(n7), .CK(clk), .Q(wo_2[30]) );
  DFFHQX1 \w_reg[1][30]  ( .D(n6), .CK(clk), .Q(wo_1[30]) );
  DFFHQX1 \w_reg[1][0]  ( .D(n126), .CK(clk), .Q(wo_1[0]) );
  DFFHQX1 \w_reg[1][1]  ( .D(n122), .CK(clk), .Q(wo_1[1]) );
  DFFHQX1 \w_reg[1][2]  ( .D(n118), .CK(clk), .Q(wo_1[2]) );
  DFFHQX1 \w_reg[1][3]  ( .D(n114), .CK(clk), .Q(wo_1[3]) );
  DFFHQX1 \w_reg[2][4]  ( .D(n111), .CK(clk), .Q(wo_2[4]) );
  DFFHQX1 \w_reg[1][4]  ( .D(n110), .CK(clk), .Q(wo_1[4]) );
  DFFHQX1 \w_reg[2][5]  ( .D(n107), .CK(clk), .Q(wo_2[5]) );
  DFFHQX1 \w_reg[1][5]  ( .D(n106), .CK(clk), .Q(wo_1[5]) );
  DFFHQX1 \w_reg[2][6]  ( .D(n103), .CK(clk), .Q(wo_2[6]) );
  DFFHQX1 \w_reg[1][6]  ( .D(n102), .CK(clk), .Q(wo_1[6]) );
  DFFHQX1 \w_reg[2][7]  ( .D(n99), .CK(clk), .Q(wo_2[7]) );
  DFFHQX1 \w_reg[1][7]  ( .D(n98), .CK(clk), .Q(wo_1[7]) );
  DFFHQX1 \w_reg[2][31]  ( .D(n3), .CK(clk), .Q(wo_2[31]) );
  DFFHQX1 \w_reg[1][31]  ( .D(n2), .CK(clk), .Q(wo_1[31]) );
  DFFHQX1 \w_reg[2][23]  ( .D(n35), .CK(clk), .Q(wo_2[23]) );
  DFFHQX1 \w_reg[1][23]  ( .D(n34), .CK(clk), .Q(wo_1[23]) );
  DFFHQX1 \w_reg[2][15]  ( .D(n67), .CK(clk), .Q(wo_2[15]) );
  DFFHQX1 \w_reg[1][15]  ( .D(n66), .CK(clk), .Q(wo_1[15]) );
  DFFHQX1 \w_reg[0][8]  ( .D(n93), .CK(clk), .Q(wo_0[8]) );
  DFFHQX1 \w_reg[0][9]  ( .D(n89), .CK(clk), .Q(wo_0[9]) );
  DFFHQX1 \w_reg[0][10]  ( .D(n85), .CK(clk), .Q(wo_0[10]) );
  DFFHQX1 \w_reg[0][11]  ( .D(n81), .CK(clk), .Q(wo_0[11]) );
  DFFHQX1 \w_reg[0][12]  ( .D(n77), .CK(clk), .Q(wo_0[12]) );
  DFFHQX1 \w_reg[0][13]  ( .D(n73), .CK(clk), .Q(wo_0[13]) );
  DFFHQX1 \w_reg[0][14]  ( .D(n69), .CK(clk), .Q(wo_0[14]) );
  DFFHQX1 \w_reg[0][16]  ( .D(n61), .CK(clk), .Q(wo_0[16]) );
  DFFHQX1 \w_reg[0][17]  ( .D(n57), .CK(clk), .Q(wo_0[17]) );
  DFFHQX1 \w_reg[0][18]  ( .D(n53), .CK(clk), .Q(wo_0[18]) );
  DFFHQX1 \w_reg[0][19]  ( .D(n49), .CK(clk), .Q(wo_0[19]) );
  DFFHQX1 \w_reg[0][20]  ( .D(n45), .CK(clk), .Q(wo_0[20]) );
  DFFHQX1 \w_reg[0][21]  ( .D(n41), .CK(clk), .Q(wo_0[21]) );
  DFFHQX1 \w_reg[0][22]  ( .D(n37), .CK(clk), .Q(wo_0[22]) );
  DFFHQX1 \w_reg[0][24]  ( .D(n29), .CK(clk), .Q(wo_0[24]) );
  DFFHQX1 \w_reg[0][25]  ( .D(n25), .CK(clk), .Q(wo_0[25]) );
  DFFHQX1 \w_reg[0][26]  ( .D(n21), .CK(clk), .Q(wo_0[26]) );
  DFFHQX1 \w_reg[0][27]  ( .D(n17), .CK(clk), .Q(wo_0[27]) );
  DFFHQX1 \w_reg[0][28]  ( .D(n13), .CK(clk), .Q(wo_0[28]) );
  DFFHQX1 \w_reg[0][29]  ( .D(n9), .CK(clk), .Q(wo_0[29]) );
  DFFHQX1 \w_reg[0][30]  ( .D(n5), .CK(clk), .Q(wo_0[30]) );
  DFFHQX1 \w_reg[0][0]  ( .D(n125), .CK(clk), .Q(wo_0[0]) );
  DFFHQX1 \w_reg[0][1]  ( .D(n121), .CK(clk), .Q(wo_0[1]) );
  DFFHQX1 \w_reg[0][2]  ( .D(n117), .CK(clk), .Q(wo_0[2]) );
  DFFHQX1 \w_reg[0][3]  ( .D(n113), .CK(clk), .Q(wo_0[3]) );
  DFFHQX1 \w_reg[0][4]  ( .D(n109), .CK(clk), .Q(wo_0[4]) );
  DFFHQX1 \w_reg[0][5]  ( .D(n105), .CK(clk), .Q(wo_0[5]) );
  DFFHQX1 \w_reg[0][6]  ( .D(n101), .CK(clk), .Q(wo_0[6]) );
  DFFHQX1 \w_reg[0][7]  ( .D(n97), .CK(clk), .Q(wo_0[7]) );
  DFFHQX1 \w_reg[0][31]  ( .D(n1), .CK(clk), .Q(wo_0[31]) );
  DFFHQX1 \w_reg[0][23]  ( .D(n33), .CK(clk), .Q(wo_0[23]) );
  DFFHQX1 \w_reg[0][15]  ( .D(n65), .CK(clk), .Q(wo_0[15]) );
  DFFHQX1 \w_reg[3][14]  ( .D(n72), .CK(clk), .Q(wo_3[14]) );
  DFFHQX1 \w_reg[3][22]  ( .D(n40), .CK(clk), .Q(wo_3[22]) );
  DFFHQX1 \w_reg[3][30]  ( .D(n8), .CK(clk), .Q(wo_3[30]) );
  DFFHQX1 \w_reg[3][6]  ( .D(n104), .CK(clk), .Q(wo_3[6]) );
  DFFHQX1 \w_reg[3][8]  ( .D(n96), .CK(clk), .Q(wo_3[8]) );
  DFFHQX1 \w_reg[3][16]  ( .D(n64), .CK(clk), .Q(wo_3[16]) );
  DFFHQX1 \w_reg[3][24]  ( .D(n32), .CK(clk), .Q(wo_3[24]) );
  DFFHQX1 \w_reg[3][0]  ( .D(n128), .CK(clk), .Q(wo_3[0]) );
  DFFHQX1 \w_reg[3][13]  ( .D(n76), .CK(clk), .Q(wo_3[13]) );
  DFFHQX1 \w_reg[3][21]  ( .D(n44), .CK(clk), .Q(wo_3[21]) );
  DFFHQX1 \w_reg[3][29]  ( .D(n12), .CK(clk), .Q(wo_3[29]) );
  DFFHQX1 \w_reg[3][5]  ( .D(n108), .CK(clk), .Q(wo_3[5]) );
  DFFHQX1 \w_reg[3][10]  ( .D(n88), .CK(clk), .Q(wo_3[10]) );
  DFFHQX1 \w_reg[3][18]  ( .D(n56), .CK(clk), .Q(wo_3[18]) );
  DFFHQX1 \w_reg[3][26]  ( .D(n24), .CK(clk), .Q(wo_3[26]) );
  DFFHQX1 \w_reg[3][2]  ( .D(n120), .CK(clk), .Q(wo_3[2]) );
  DFFHQX1 \w_reg[3][12]  ( .D(n80), .CK(clk), .Q(wo_3[12]) );
  DFFHQX1 \w_reg[3][20]  ( .D(n48), .CK(clk), .Q(wo_3[20]) );
  DFFHQX1 \w_reg[3][28]  ( .D(n16), .CK(clk), .Q(wo_3[28]) );
  DFFHQX1 \w_reg[3][4]  ( .D(n112), .CK(clk), .Q(wo_3[4]) );
  DFFHQX1 \w_reg[3][11]  ( .D(n84), .CK(clk), .Q(wo_3[11]) );
  DFFHQX1 \w_reg[3][19]  ( .D(n52), .CK(clk), .Q(wo_3[19]) );
  DFFHQX1 \w_reg[3][27]  ( .D(n20), .CK(clk), .Q(wo_3[27]) );
  DFFHQX1 \w_reg[3][3]  ( .D(n116), .CK(clk), .Q(wo_3[3]) );
  XOR2X1 U404 ( .A(wo_0[24]), .B(subword[24]), .Y(n265) );
  XOR2X1 U372 ( .A(wo_0[8]), .B(subword[8]), .Y(N33) );
  XOR2X1 U356 ( .A(wo_0[0]), .B(subword[0]), .Y(N41) );
  XOR2X1 U388 ( .A(wo_0[16]), .B(subword[16]), .Y(N25) );
  XOR2X1 U360 ( .A(wo_0[2]), .B(subword[2]), .Y(N39) );
  XOR2X1 U384 ( .A(wo_0[14]), .B(subword[14]), .Y(N27) );
  XOR2X1 U398 ( .A(wo_0[21]), .B(subword[21]), .Y(N20) );
  XOR2X1 U408 ( .A(wo_0[26]), .B(subword[26]), .Y(n263) );
  XOR2X1 U416 ( .A(wo_0[30]), .B(subword[30]), .Y(n259) );
  XOR2X1 U324 ( .A(wo_1[0]), .B(N41), .Y(N107) );
  XOR2X1 U410 ( .A(wo_0[27]), .B(subword[27]), .Y(n262) );
  XOR2X1 U400 ( .A(wo_0[22]), .B(subword[22]), .Y(N19) );
  XOR2X1 U376 ( .A(wo_0[10]), .B(subword[10]), .Y(N31) );
  XOR2X1 U382 ( .A(wo_0[13]), .B(subword[13]), .Y(N28) );
  XOR2X1 U405 ( .A(rcon[24]), .B(n265), .Y(N17) );
  XOR2X1 U378 ( .A(wo_0[11]), .B(subword[11]), .Y(N30) );
  XOR2X1 U362 ( .A(wo_0[3]), .B(subword[3]), .Y(N38) );
  XOR2X1 U414 ( .A(wo_0[29]), .B(subword[29]), .Y(n260) );
  XOR2X1 U332 ( .A(wo_1[8]), .B(N33), .Y(N99) );
  XOR2X1 U392 ( .A(wo_0[18]), .B(subword[18]), .Y(N23) );
  XOR2X1 U340 ( .A(wo_1[16]), .B(N25), .Y(N91) );
  XOR2X1 U394 ( .A(wo_0[19]), .B(subword[19]), .Y(N22) );
  XOR2X1 U366 ( .A(wo_0[5]), .B(subword[5]), .Y(N36) );
  XOR2X1 U368 ( .A(wo_0[6]), .B(subword[6]), .Y(N35) );
  XOR2X1 U308 ( .A(wo_2[16]), .B(N91), .Y(N157) );
  XOR2X1 U396 ( .A(wo_0[20]), .B(subword[20]), .Y(N21) );
  XOR2X1 U415 ( .A(rcon[29]), .B(n260), .Y(N12) );
  XOR2X1 U412 ( .A(wo_0[28]), .B(subword[28]), .Y(n261) );
  XOR2X1 U402 ( .A(wo_0[23]), .B(subword[23]), .Y(N18) );
  XOR2X1 U334 ( .A(wo_1[10]), .B(N31), .Y(N97) );
  XOR2X1 U300 ( .A(wo_2[8]), .B(N99), .Y(N165) );
  XOR2X1 U326 ( .A(wo_1[2]), .B(N39), .Y(N105) );
  XOR2X1 U292 ( .A(wo_2[0]), .B(N107), .Y(N173) );
  XOR2X1 U411 ( .A(rcon[27]), .B(n262), .Y(N14) );
  XOR2X1 U380 ( .A(wo_0[12]), .B(subword[12]), .Y(N29) );
  XOR2X1 U417 ( .A(rcon[30]), .B(n259), .Y(N11) );
  XOR2X1 U345 ( .A(wo_1[21]), .B(N20), .Y(N86) );
  XOR2X1 U343 ( .A(wo_1[19]), .B(N22), .Y(N88) );
  XOR2X1 U409 ( .A(rcon[26]), .B(n263), .Y(N15) );
  XOR2X1 U330 ( .A(wo_1[6]), .B(N35), .Y(N101) );
  XOR2X1 U338 ( .A(wo_1[14]), .B(N27), .Y(N93) );
  XOR2X1 U342 ( .A(wo_1[18]), .B(N23), .Y(N89) );
  XOR2X1 U348 ( .A(wo_1[24]), .B(N17), .Y(N83) );
  XOR2X1 U335 ( .A(wo_1[11]), .B(N30), .Y(N96) );
  XOR2X1 U337 ( .A(wo_1[13]), .B(N28), .Y(N94) );
  XOR2X1 U327 ( .A(wo_1[3]), .B(N38), .Y(N104) );
  XOR2X1 U418 ( .A(wo_0[31]), .B(subword[31]), .Y(n258) );
  XOR2X1 U329 ( .A(wo_1[5]), .B(N36), .Y(N102) );
  XOR2X1 U386 ( .A(wo_0[15]), .B(subword[15]), .Y(N26) );
  XOR2X1 U346 ( .A(wo_1[22]), .B(N19), .Y(N85) );
  XOR2X1 U370 ( .A(wo_0[7]), .B(subword[7]), .Y(N34) );
  XOR2X1 U364 ( .A(wo_0[4]), .B(subword[4]), .Y(N37) );
  XOR2X1 U310 ( .A(wo_2[18]), .B(N89), .Y(N155) );
  XOR2X1 U419 ( .A(rcon[31]), .B(n258), .Y(N10) );
  XOR2X1 U311 ( .A(wo_2[19]), .B(N88), .Y(N154) );
  XOR2X1 U390 ( .A(wo_0[17]), .B(subword[17]), .Y(N24) );
  XOR2X1 U298 ( .A(wo_2[6]), .B(N101), .Y(N167) );
  XOR2X1 U306 ( .A(wo_2[14]), .B(N93), .Y(N159) );
  XOR2X1 U354 ( .A(wo_1[30]), .B(N11), .Y(N77) );
  XOR2X1 U328 ( .A(wo_1[4]), .B(N37), .Y(N103) );
  XOR2X1 U344 ( .A(wo_1[20]), .B(N21), .Y(N87) );
  XOR2X1 U297 ( .A(wo_2[5]), .B(N102), .Y(N168) );
  XOR2X1 U339 ( .A(wo_1[15]), .B(N26), .Y(N92) );
  XOR2X1 U313 ( .A(wo_2[21]), .B(N86), .Y(N152) );
  XOR2X1 U358 ( .A(wo_0[1]), .B(subword[1]), .Y(N40) );
  XOR2X1 U303 ( .A(wo_2[11]), .B(N96), .Y(N162) );
  XOR2X1 U295 ( .A(wo_2[3]), .B(N104), .Y(N170) );
  XOR2X1 U302 ( .A(wo_2[10]), .B(N97), .Y(N163) );
  XOR2X1 U353 ( .A(wo_1[29]), .B(N12), .Y(N78) );
  XOR2X1 U406 ( .A(wo_0[25]), .B(subword[25]), .Y(n264) );
  XOR2X1 U413 ( .A(rcon[28]), .B(n261), .Y(N13) );
  XOR2X1 U336 ( .A(wo_1[12]), .B(N29), .Y(N95) );
  XOR2X1 U374 ( .A(wo_0[9]), .B(subword[9]), .Y(N32) );
  XOR2X1 U347 ( .A(wo_1[23]), .B(N18), .Y(N84) );
  XOR2X1 U316 ( .A(wo_2[24]), .B(N83), .Y(N149) );
  XOR2X1 U294 ( .A(wo_2[2]), .B(N105), .Y(N171) );
  XOR2X1 U350 ( .A(wo_1[26]), .B(N15), .Y(N81) );
  XOR2X1 U331 ( .A(wo_1[7]), .B(N34), .Y(N100) );
  XOR2X1 U351 ( .A(wo_1[27]), .B(N14), .Y(N80) );
  XOR2X1 U305 ( .A(wo_2[13]), .B(N94), .Y(N160) );
  XOR2X1 U314 ( .A(wo_2[22]), .B(N85), .Y(N151) );
  XOR2X1 U325 ( .A(wo_1[1]), .B(N40), .Y(N106) );
  XOR2X1 U296 ( .A(wo_2[4]), .B(N103), .Y(N169) );
  XOR2X1 U319 ( .A(wo_2[27]), .B(N80), .Y(N146) );
  XOR2X1 U322 ( .A(wo_2[30]), .B(N77), .Y(N143) );
  XOR2X1 U299 ( .A(wo_2[7]), .B(N100), .Y(N166) );
  XOR2X1 U352 ( .A(wo_1[28]), .B(N13), .Y(N79) );
  XOR2X1 U307 ( .A(wo_2[15]), .B(N92), .Y(N158) );
  XOR2X1 U304 ( .A(wo_2[12]), .B(N95), .Y(N161) );
  XOR2X1 U312 ( .A(wo_2[20]), .B(N87), .Y(N153) );
  XOR2X1 U315 ( .A(wo_2[23]), .B(N84), .Y(N150) );
  XOR2X1 U321 ( .A(wo_2[29]), .B(N78), .Y(N144) );
  XOR2X1 U341 ( .A(wo_1[17]), .B(N24), .Y(N90) );
  XOR2X1 U318 ( .A(wo_2[26]), .B(N81), .Y(N147) );
  XOR2X1 U333 ( .A(wo_1[9]), .B(N32), .Y(N98) );
  XOR2X1 U407 ( .A(rcon[25]), .B(n264), .Y(N16) );
  XOR2X1 U355 ( .A(wo_1[31]), .B(N10), .Y(N76) );
  XOR2X1 U309 ( .A(wo_2[17]), .B(N90), .Y(N156) );
  XOR2X1 U349 ( .A(wo_1[25]), .B(N16), .Y(N82) );
  XOR2X1 U293 ( .A(wo_2[1]), .B(N106), .Y(N172) );
  XOR2X1 U320 ( .A(wo_2[28]), .B(N79), .Y(N145) );
  XOR2X1 U323 ( .A(wo_2[31]), .B(N76), .Y(N142) );
  XOR2X1 U301 ( .A(wo_2[9]), .B(N98), .Y(N164) );
  XOR2X1 U317 ( .A(wo_2[25]), .B(N82), .Y(N148) );
  DFFX2 \w_reg[3][17]  ( .D(n255), .CK(clk), .QN(wo_3[17]) );
  DFFX2 \w_reg[3][1]  ( .D(n203), .CK(clk), .QN(wo_3[1]) );
  DFFX2 \w_reg[3][9]  ( .D(n229), .CK(clk), .QN(wo_3[9]) );
  DFFX2 \w_reg[3][23]  ( .D(n282), .CK(clk), .QN(wo_3[23]) );
  DFFX2 \w_reg[3][7]  ( .D(n222), .CK(clk), .QN(wo_3[7]) );
  DFFX2 \w_reg[3][15]  ( .D(n248), .CK(clk), .QN(wo_3[15]) );
  DFFX2 \w_reg[3][31]  ( .D(n308), .CK(clk), .QN(wo_3[31]) );
  DFFX2 \w_reg[3][25]  ( .D(n289), .CK(clk), .QN(wo_3[25]) );
  NAND2X1 U3 ( .A(wo_3[11]), .B(N162), .Y(n4) );
  OAI211X1 U4 ( .A0(wo_3[11]), .A1(N162), .B0(n192), .C0(n4), .Y(n28) );
  OAI2BB1X1 U5 ( .A0N(key[11]), .A1N(kld), .B0(n28), .Y(n84) );
  OAI21XL U6 ( .A0(wo_3[25]), .A1(N148), .B0(n199), .Y(n36) );
  AOI21X1 U7 ( .A0(wo_3[25]), .A1(N148), .B0(n36), .Y(n60) );
  AOI21X1 U8 ( .A0(key[25]), .A1(kld), .B0(n60), .Y(n289) );
  NAND2X1 U9 ( .A(wo_3[27]), .B(N146), .Y(n68) );
  OAI211X1 U10 ( .A0(wo_3[27]), .A1(N146), .B0(n198), .C0(n68), .Y(n92) );
  OAI2BB1X1 U11 ( .A0N(key[27]), .A1N(kld), .B0(n92), .Y(n20) );
  NAND2X1 U12 ( .A(wo_3[28]), .B(N145), .Y(n100) );
  OAI211X1 U13 ( .A0(wo_3[28]), .A1(N145), .B0(n196), .C0(n100), .Y(n124) );
  OAI2BB1X1 U14 ( .A0N(key[28]), .A1N(kld), .B0(n124), .Y(n16) );
  NAND2X1 U15 ( .A(wo_3[12]), .B(N161), .Y(n129) );
  OAI211X1 U16 ( .A0(wo_3[12]), .A1(N161), .B0(n192), .C0(n129), .Y(n130) );
  OAI2BB1X1 U17 ( .A0N(key[12]), .A1N(kld), .B0(n130), .Y(n80) );
  OAI21XL U18 ( .A0(wo_3[31]), .A1(N142), .B0(n191), .Y(n131) );
  AOI21X1 U19 ( .A0(wo_3[31]), .A1(N142), .B0(n131), .Y(n132) );
  AOI21X1 U20 ( .A0(key[31]), .A1(kld), .B0(n132), .Y(n308) );
  OAI21XL U21 ( .A0(wo_3[15]), .A1(N158), .B0(n194), .Y(n133) );
  AOI21X1 U22 ( .A0(wo_3[15]), .A1(N158), .B0(n133), .Y(n134) );
  AOI21X1 U23 ( .A0(key[15]), .A1(kld), .B0(n134), .Y(n248) );
  OAI21XL U24 ( .A0(wo_3[23]), .A1(N150), .B0(n197), .Y(n135) );
  AOI21X1 U25 ( .A0(wo_3[23]), .A1(N150), .B0(n135), .Y(n136) );
  AOI21X1 U26 ( .A0(key[23]), .A1(kld), .B0(n136), .Y(n282) );
  OAI21XL U27 ( .A0(wo_3[17]), .A1(N156), .B0(n195), .Y(n137) );
  AOI21X1 U28 ( .A0(wo_3[17]), .A1(N156), .B0(n137), .Y(n138) );
  AOI21X1 U29 ( .A0(key[17]), .A1(kld), .B0(n138), .Y(n255) );
  NAND2X1 U30 ( .A(wo_3[3]), .B(N170), .Y(n139) );
  OAI211X1 U31 ( .A0(wo_3[3]), .A1(N170), .B0(n186), .C0(n139), .Y(n140) );
  OAI2BB1X1 U32 ( .A0N(key[3]), .A1N(kld), .B0(n140), .Y(n116) );
  NAND2X1 U33 ( .A(wo_3[19]), .B(N154), .Y(n141) );
  OAI211X1 U34 ( .A0(wo_3[19]), .A1(N154), .B0(n198), .C0(n141), .Y(n142) );
  OAI2BB1X1 U35 ( .A0N(key[19]), .A1N(kld), .B0(n142), .Y(n52) );
  NAND2X1 U36 ( .A(wo_3[4]), .B(N169), .Y(n143) );
  OAI211X1 U37 ( .A0(wo_3[4]), .A1(N169), .B0(n187), .C0(n143), .Y(n144) );
  OAI2BB1X1 U38 ( .A0N(key[4]), .A1N(kld), .B0(n144), .Y(n112) );
  NAND2X1 U39 ( .A(wo_3[20]), .B(N153), .Y(n145) );
  OAI211X1 U40 ( .A0(wo_3[20]), .A1(N153), .B0(n196), .C0(n145), .Y(n146) );
  OAI2BB1X1 U41 ( .A0N(key[20]), .A1N(kld), .B0(n146), .Y(n48) );
  NAND2X1 U42 ( .A(wo_3[5]), .B(N168), .Y(n147) );
  OAI211X1 U43 ( .A0(wo_3[5]), .A1(N168), .B0(n188), .C0(n147), .Y(n148) );
  OAI2BB1X1 U44 ( .A0N(key[5]), .A1N(kld), .B0(n148), .Y(n108) );
  NAND2X1 U45 ( .A(wo_3[16]), .B(N157), .Y(n149) );
  OAI211X1 U46 ( .A0(wo_3[16]), .A1(N157), .B0(n192), .C0(n149), .Y(n150) );
  OAI2BB1X1 U47 ( .A0N(key[16]), .A1N(kld), .B0(n150), .Y(n64) );
  NAND2X1 U48 ( .A(wo_3[8]), .B(N165), .Y(n151) );
  OAI211X1 U49 ( .A0(wo_3[8]), .A1(N165), .B0(n190), .C0(n151), .Y(n152) );
  OAI2BB1X1 U50 ( .A0N(key[8]), .A1N(kld), .B0(n152), .Y(n96) );
  NAND2X1 U51 ( .A(wo_3[30]), .B(N143), .Y(n153) );
  OAI211X1 U52 ( .A0(wo_3[30]), .A1(N143), .B0(n199), .C0(n153), .Y(n154) );
  OAI2BB1X1 U53 ( .A0N(key[30]), .A1N(kld), .B0(n154), .Y(n8) );
  OAI21XL U54 ( .A0(wo_3[7]), .A1(N166), .B0(n189), .Y(n155) );
  AOI21X1 U55 ( .A0(wo_3[7]), .A1(N166), .B0(n155), .Y(n156) );
  AOI21X1 U56 ( .A0(key[7]), .A1(kld), .B0(n156), .Y(n222) );
  OAI21XL U57 ( .A0(wo_3[9]), .A1(N164), .B0(n190), .Y(n157) );
  AOI21X1 U58 ( .A0(wo_3[9]), .A1(N164), .B0(n157), .Y(n158) );
  AOI21X1 U59 ( .A0(key[9]), .A1(kld), .B0(n158), .Y(n229) );
  OAI21XL U60 ( .A0(wo_3[1]), .A1(N172), .B0(n185), .Y(n159) );
  AOI21X1 U61 ( .A0(wo_3[1]), .A1(N172), .B0(n159), .Y(n160) );
  AOI21X1 U62 ( .A0(key[1]), .A1(kld), .B0(n160), .Y(n203) );
  NAND2X1 U63 ( .A(wo_3[2]), .B(N171), .Y(n161) );
  OAI211X1 U64 ( .A0(wo_3[2]), .A1(N171), .B0(n186), .C0(n161), .Y(n162) );
  OAI2BB1X1 U65 ( .A0N(key[2]), .A1N(kld), .B0(n162), .Y(n120) );
  NAND2X1 U66 ( .A(wo_3[26]), .B(N147), .Y(n163) );
  OAI211X1 U67 ( .A0(wo_3[26]), .A1(N147), .B0(n198), .C0(n163), .Y(n164) );
  OAI2BB1X1 U68 ( .A0N(key[26]), .A1N(kld), .B0(n164), .Y(n24) );
  NAND2X1 U69 ( .A(wo_3[18]), .B(N155), .Y(n165) );
  OAI211X1 U70 ( .A0(wo_3[18]), .A1(N155), .B0(n195), .C0(n165), .Y(n166) );
  OAI2BB1X1 U71 ( .A0N(key[18]), .A1N(kld), .B0(n166), .Y(n56) );
  NAND2X1 U72 ( .A(wo_3[10]), .B(N163), .Y(n167) );
  OAI211X1 U73 ( .A0(wo_3[10]), .A1(N163), .B0(n191), .C0(n167), .Y(n168) );
  OAI2BB1X1 U74 ( .A0N(key[10]), .A1N(kld), .B0(n168), .Y(n88) );
  NAND2X1 U75 ( .A(wo_3[29]), .B(N144), .Y(n169) );
  OAI211X1 U76 ( .A0(wo_3[29]), .A1(N144), .B0(n199), .C0(n169), .Y(n170) );
  OAI2BB1X1 U77 ( .A0N(key[29]), .A1N(kld), .B0(n170), .Y(n12) );
  NAND2X1 U78 ( .A(wo_3[21]), .B(N152), .Y(n171) );
  OAI211X1 U79 ( .A0(wo_3[21]), .A1(N152), .B0(n196), .C0(n171), .Y(n172) );
  OAI2BB1X1 U80 ( .A0N(key[21]), .A1N(kld), .B0(n172), .Y(n44) );
  NAND2X1 U81 ( .A(wo_3[13]), .B(N160), .Y(n173) );
  OAI211X1 U82 ( .A0(wo_3[13]), .A1(N160), .B0(n193), .C0(n173), .Y(n174) );
  OAI2BB1X1 U83 ( .A0N(key[13]), .A1N(kld), .B0(n174), .Y(n76) );
  NAND2X1 U84 ( .A(wo_3[0]), .B(N173), .Y(n175) );
  OAI211X1 U85 ( .A0(wo_3[0]), .A1(N173), .B0(n187), .C0(n175), .Y(n176) );
  OAI2BB1X1 U86 ( .A0N(key[0]), .A1N(kld), .B0(n176), .Y(n128) );
  NAND2X1 U87 ( .A(wo_3[24]), .B(N149), .Y(n177) );
  OAI211X1 U88 ( .A0(wo_3[24]), .A1(N149), .B0(n197), .C0(n177), .Y(n178) );
  OAI2BB1X1 U89 ( .A0N(key[24]), .A1N(kld), .B0(n178), .Y(n32) );
  NAND2X1 U90 ( .A(wo_3[6]), .B(N167), .Y(n179) );
  OAI211X1 U91 ( .A0(wo_3[6]), .A1(N167), .B0(n188), .C0(n179), .Y(n180) );
  OAI2BB1X1 U92 ( .A0N(key[6]), .A1N(kld), .B0(n180), .Y(n104) );
  NAND2X1 U93 ( .A(wo_3[22]), .B(N151), .Y(n181) );
  OAI211X1 U94 ( .A0(wo_3[22]), .A1(N151), .B0(n192), .C0(n181), .Y(n182) );
  OAI2BB1X1 U95 ( .A0N(key[22]), .A1N(kld), .B0(n182), .Y(n40) );
  NAND2X1 U96 ( .A(wo_3[14]), .B(N159), .Y(n183) );
  OAI211X1 U97 ( .A0(wo_3[14]), .A1(N159), .B0(n194), .C0(n183), .Y(n184) );
  OAI2BB1X1 U98 ( .A0N(key[14]), .A1N(kld), .B0(n184), .Y(n72) );
  INVX1 U99 ( .A(kld), .Y(n196) );
  INVX1 U100 ( .A(kld), .Y(n194) );
  INVX1 U101 ( .A(kld), .Y(n188) );
  INVX1 U102 ( .A(kld), .Y(n186) );
  INVX1 U103 ( .A(kld), .Y(n195) );
  INVX1 U104 ( .A(kld), .Y(n190) );
  INVX1 U105 ( .A(kld), .Y(n191) );
  INVX1 U106 ( .A(kld), .Y(n189) );
  INVX1 U107 ( .A(kld), .Y(n185) );
  INVX1 U108 ( .A(kld), .Y(n187) );
  AOI22XL U109 ( .A0(kld), .A1(key[79]), .B0(N92), .B1(n193), .Y(n250) );
  AOI22XL U110 ( .A0(kld), .A1(key[68]), .B0(N103), .B1(n187), .Y(n214) );
  AOI22XL U111 ( .A0(kld), .A1(key[87]), .B0(N84), .B1(n197), .Y(n284) );
  AOI22XL U112 ( .A0(kld), .A1(key[93]), .B0(N78), .B1(n199), .Y(n303) );
  AOI22XL U113 ( .A0(kld), .A1(key[94]), .B0(N77), .B1(n193), .Y(n306) );
  AOI22XL U114 ( .A0(kld), .A1(key[83]), .B0(N88), .B1(n192), .Y(n271) );
  AOI22XL U115 ( .A0(kld), .A1(key[88]), .B0(N83), .B1(n192), .Y(n287) );
  INVX2 U116 ( .A(kld), .Y(n198) );
  INVX2 U117 ( .A(kld), .Y(n193) );
  INVX1 U118 ( .A(kld), .Y(n199) );
  INVX2 U119 ( .A(kld), .Y(n192) );
  INVX1 U120 ( .A(kld), .Y(n197) );
  AOI22XL U121 ( .A0(kld), .A1(key[81]), .B0(N90), .B1(n195), .Y(n257) );
  AOI22XL U122 ( .A0(kld), .A1(key[95]), .B0(N76), .B1(n189), .Y(n310) );
  AOI22XL U123 ( .A0(kld), .A1(key[73]), .B0(N98), .B1(n191), .Y(n231) );
  AOI22XL U124 ( .A0(kld), .A1(key[92]), .B0(N79), .B1(n186), .Y(n300) );
  AOI22XL U125 ( .A0(kld), .A1(key[65]), .B0(N106), .B1(n185), .Y(n205) );
  AOI22XL U126 ( .A0(kld), .A1(key[91]), .B0(N80), .B1(n195), .Y(n297) );
  AOI22XL U127 ( .A0(kld), .A1(key[71]), .B0(N100), .B1(n189), .Y(n224) );
  AOI22XL U128 ( .A0(kld), .A1(key[84]), .B0(N87), .B1(n196), .Y(n274) );
  AOI22XL U129 ( .A0(kld), .A1(key[76]), .B0(N95), .B1(n193), .Y(n240) );
  AOI22XL U130 ( .A0(kld), .A1(key[90]), .B0(N81), .B1(n198), .Y(n294) );
  AOI22XL U131 ( .A0(kld), .A1(key[85]), .B0(N86), .B1(n191), .Y(n277) );
  AOI22XL U132 ( .A0(kld), .A1(key[75]), .B0(N96), .B1(n192), .Y(n237) );
  AOI22XL U133 ( .A0(kld), .A1(key[66]), .B0(N105), .B1(n186), .Y(n208) );
  AOI22XL U134 ( .A0(kld), .A1(key[67]), .B0(N104), .B1(n187), .Y(n211) );
  AOI22XL U135 ( .A0(kld), .A1(key[86]), .B0(N85), .B1(n198), .Y(n280) );
  AOI22XL U136 ( .A0(kld), .A1(key[78]), .B0(N93), .B1(n194), .Y(n246) );
  AOI22XL U137 ( .A0(kld), .A1(key[69]), .B0(N102), .B1(n188), .Y(n217) );
  AOI22XL U138 ( .A0(kld), .A1(key[77]), .B0(N94), .B1(n193), .Y(n243) );
  AOI22XL U139 ( .A0(kld), .A1(key[74]), .B0(N97), .B1(n191), .Y(n234) );
  AOI22XL U140 ( .A0(kld), .A1(key[70]), .B0(N101), .B1(n189), .Y(n220) );
  AOI22XL U141 ( .A0(kld), .A1(key[82]), .B0(N89), .B1(n198), .Y(n268) );
  AOI22XL U142 ( .A0(kld), .A1(key[80]), .B0(N91), .B1(n192), .Y(n253) );
  AOI22XL U143 ( .A0(kld), .A1(key[64]), .B0(N107), .B1(n185), .Y(n201) );
  AOI22XL U144 ( .A0(kld), .A1(key[72]), .B0(N99), .B1(n190), .Y(n227) );
  INVXL U145 ( .A(n290), .Y(n27) );
  INVXL U146 ( .A(n230), .Y(n91) );
  INVXL U147 ( .A(n204), .Y(n123) );
  INVXL U148 ( .A(n291), .Y(n26) );
  INVXL U149 ( .A(n299), .Y(n15) );
  INVXL U150 ( .A(n309), .Y(n3) );
  INVXL U151 ( .A(n256), .Y(n59) );
  INVXL U152 ( .A(n239), .Y(n79) );
  INVXL U153 ( .A(n300), .Y(n14) );
  INVXL U154 ( .A(n302), .Y(n11) );
  INVXL U155 ( .A(n283), .Y(n35) );
  INVXL U156 ( .A(n273), .Y(n47) );
  INVXL U157 ( .A(n249), .Y(n67) );
  INVXL U158 ( .A(n293), .Y(n23) );
  INVXL U159 ( .A(n223), .Y(n99) );
  INVXL U160 ( .A(n205), .Y(n122) );
  INVXL U161 ( .A(n231), .Y(n90) );
  INVXL U162 ( .A(n296), .Y(n19) );
  INVXL U163 ( .A(n305), .Y(n7) );
  AOI22XL U164 ( .A0(kld), .A1(key[89]), .B0(N82), .B1(n197), .Y(n291) );
  INVXL U165 ( .A(n257), .Y(n58) );
  INVXL U166 ( .A(n292), .Y(n25) );
  INVXL U167 ( .A(n310), .Y(n2) );
  INVXL U168 ( .A(n213), .Y(n111) );
  INVXL U169 ( .A(n232), .Y(n89) );
  INVXL U170 ( .A(n311), .Y(n1) );
  INVXL U171 ( .A(n216), .Y(n107) );
  INVXL U172 ( .A(n214), .Y(n110) );
  INVXL U173 ( .A(n219), .Y(n103) );
  INVXL U174 ( .A(n306), .Y(n6) );
  INVXL U175 ( .A(n294), .Y(n22) );
  INVXL U176 ( .A(n207), .Y(n119) );
  INVXL U177 ( .A(n297), .Y(n18) );
  INVXL U178 ( .A(n224), .Y(n98) );
  INVXL U179 ( .A(n301), .Y(n13) );
  INVXL U180 ( .A(n303), .Y(n10) );
  INVXL U181 ( .A(n210), .Y(n115) );
  INVXL U182 ( .A(n276), .Y(n43) );
  INVXL U183 ( .A(n279), .Y(n39) );
  INVXL U184 ( .A(n242), .Y(n75) );
  INVXL U185 ( .A(n274), .Y(n46) );
  INVXL U186 ( .A(n284), .Y(n34) );
  INVXL U187 ( .A(n240), .Y(n78) );
  INVXL U188 ( .A(n250), .Y(n66) );
  INVXL U189 ( .A(n270), .Y(n51) );
  INVXL U190 ( .A(n236), .Y(n83) );
  INVXL U191 ( .A(n267), .Y(n55) );
  INVXL U192 ( .A(n206), .Y(n121) );
  INVXL U193 ( .A(n286), .Y(n31) );
  INVXL U194 ( .A(n245), .Y(n71) );
  INVXL U195 ( .A(n233), .Y(n87) );
  AOI22XL U196 ( .A0(kld), .A1(key[121]), .B0(N16), .B1(n189), .Y(n292) );
  INVXL U197 ( .A(n266), .Y(n57) );
  INVXL U198 ( .A(n220), .Y(n102) );
  INVXL U199 ( .A(n287), .Y(n30) );
  AOI22XL U200 ( .A0(kld), .A1(key[105]), .B0(N32), .B1(n191), .Y(n232) );
  INVXL U201 ( .A(n295), .Y(n21) );
  INVXL U202 ( .A(n217), .Y(n106) );
  AOI22XL U203 ( .A0(kld), .A1(key[127]), .B0(N10), .B1(n188), .Y(n311) );
  INVXL U204 ( .A(n234), .Y(n86) );
  INVXL U205 ( .A(n252), .Y(n63) );
  AOI22XL U206 ( .A0(kld), .A1(key[113]), .B0(N24), .B1(n195), .Y(n266) );
  INVXL U207 ( .A(n277), .Y(n42) );
  INVXL U208 ( .A(n280), .Y(n38) );
  INVXL U209 ( .A(n304), .Y(n9) );
  INVXL U210 ( .A(n275), .Y(n45) );
  INVXL U211 ( .A(n285), .Y(n33) );
  INVXL U212 ( .A(n241), .Y(n77) );
  INVXL U213 ( .A(n246), .Y(n70) );
  AOI22XL U214 ( .A0(kld), .A1(key[124]), .B0(N13), .B1(n190), .Y(n301) );
  INVXL U215 ( .A(n225), .Y(n97) );
  INVXL U216 ( .A(n251), .Y(n65) );
  INVXL U217 ( .A(n271), .Y(n50) );
  INVXL U218 ( .A(n237), .Y(n82) );
  INVXL U219 ( .A(n298), .Y(n17) );
  INVXL U220 ( .A(n226), .Y(n95) );
  INVXL U221 ( .A(n268), .Y(n54) );
  INVXL U222 ( .A(n307), .Y(n5) );
  INVXL U223 ( .A(n243), .Y(n74) );
  INVXL U224 ( .A(n208), .Y(n118) );
  AOI22XL U225 ( .A0(kld), .A1(key[97]), .B0(N40), .B1(n185), .Y(n206) );
  INVXL U226 ( .A(n200), .Y(n127) );
  INVXL U227 ( .A(n211), .Y(n114) );
  INVXL U228 ( .A(n215), .Y(n109) );
  INVXL U229 ( .A(n244), .Y(n73) );
  AOI22XL U230 ( .A0(kld), .A1(key[122]), .B0(N15), .B1(n198), .Y(n295) );
  AOI22XL U231 ( .A0(kld), .A1(key[103]), .B0(N34), .B1(n189), .Y(n225) );
  INVXL U232 ( .A(n209), .Y(n117) );
  AOI22XL U233 ( .A0(kld), .A1(key[123]), .B0(N14), .B1(n198), .Y(n298) );
  INVXL U234 ( .A(n227), .Y(n94) );
  INVXL U235 ( .A(n281), .Y(n37) );
  AOI22XL U236 ( .A0(kld), .A1(key[119]), .B0(N18), .B1(n197), .Y(n285) );
  AOI22XL U237 ( .A0(kld), .A1(key[108]), .B0(N29), .B1(n193), .Y(n241) );
  AOI22XL U238 ( .A0(kld), .A1(key[125]), .B0(N12), .B1(n199), .Y(n304) );
  INVXL U239 ( .A(n212), .Y(n113) );
  INVXL U240 ( .A(n235), .Y(n85) );
  INVXL U241 ( .A(n238), .Y(n81) );
  INVXL U242 ( .A(n288), .Y(n29) );
  AOI22XL U243 ( .A0(kld), .A1(key[100]), .B0(N37), .B1(n187), .Y(n215) );
  INVXL U244 ( .A(n201), .Y(n126) );
  AOI22XL U245 ( .A0(kld), .A1(key[111]), .B0(N26), .B1(n198), .Y(n251) );
  INVXL U246 ( .A(n278), .Y(n41) );
  AOI22XL U247 ( .A0(kld), .A1(key[126]), .B0(N11), .B1(n193), .Y(n307) );
  INVXL U248 ( .A(n247), .Y(n69) );
  INVXL U249 ( .A(n253), .Y(n62) );
  AOI22XL U250 ( .A0(kld), .A1(key[116]), .B0(N21), .B1(n196), .Y(n275) );
  INVXL U251 ( .A(n218), .Y(n105) );
  INVXL U252 ( .A(n269), .Y(n53) );
  INVXL U253 ( .A(n221), .Y(n101) );
  INVXL U254 ( .A(n272), .Y(n49) );
  AOI22XL U255 ( .A0(kld), .A1(key[106]), .B0(N31), .B1(n191), .Y(n235) );
  AOI22XL U256 ( .A0(kld), .A1(key[114]), .B0(N23), .B1(n193), .Y(n269) );
  AOI22XL U257 ( .A0(kld), .A1(key[118]), .B0(N19), .B1(n187), .Y(n281) );
  AOI22XL U258 ( .A0(kld), .A1(key[107]), .B0(N30), .B1(n192), .Y(n238) );
  AOI22XL U259 ( .A0(kld), .A1(key[101]), .B0(N36), .B1(n188), .Y(n218) );
  AOI22XL U260 ( .A0(kld), .A1(key[109]), .B0(N28), .B1(n193), .Y(n244) );
  AOI22XL U261 ( .A0(kld), .A1(key[120]), .B0(N17), .B1(n192), .Y(n288) );
  AOI22XL U262 ( .A0(kld), .A1(key[110]), .B0(N27), .B1(n194), .Y(n247) );
  INVXL U263 ( .A(n254), .Y(n61) );
  AOI22XL U264 ( .A0(kld), .A1(key[99]), .B0(N38), .B1(n187), .Y(n212) );
  INVXL U265 ( .A(n202), .Y(n125) );
  AOI22XL U266 ( .A0(kld), .A1(key[98]), .B0(N39), .B1(n186), .Y(n209) );
  AOI22XL U267 ( .A0(kld), .A1(key[117]), .B0(N20), .B1(n185), .Y(n278) );
  AOI22XL U268 ( .A0(kld), .A1(key[102]), .B0(N35), .B1(n189), .Y(n221) );
  INVXL U269 ( .A(n228), .Y(n93) );
  AOI22XL U270 ( .A0(kld), .A1(key[115]), .B0(N22), .B1(n192), .Y(n272) );
  AOI22XL U271 ( .A0(kld), .A1(key[112]), .B0(N25), .B1(n193), .Y(n254) );
  AOI22XL U272 ( .A0(kld), .A1(key[96]), .B0(N41), .B1(n185), .Y(n202) );
  AOI22XL U273 ( .A0(kld), .A1(key[104]), .B0(N33), .B1(n190), .Y(n228) );
  AOI22X1 U274 ( .A0(kld), .A1(key[32]), .B0(N173), .B1(n185), .Y(n200) );
  AOI22X1 U275 ( .A0(kld), .A1(key[33]), .B0(N172), .B1(n185), .Y(n204) );
  AOI22X1 U276 ( .A0(kld), .A1(key[34]), .B0(N171), .B1(n186), .Y(n207) );
  AOI22X1 U277 ( .A0(kld), .A1(key[35]), .B0(N170), .B1(n186), .Y(n210) );
  AOI22X1 U278 ( .A0(kld), .A1(key[36]), .B0(N169), .B1(n187), .Y(n213) );
  AOI22X1 U279 ( .A0(kld), .A1(key[37]), .B0(N168), .B1(n188), .Y(n216) );
  AOI22X1 U280 ( .A0(kld), .A1(key[38]), .B0(N167), .B1(n188), .Y(n219) );
  AOI22X1 U281 ( .A0(kld), .A1(key[39]), .B0(N166), .B1(n189), .Y(n223) );
  AOI22X1 U282 ( .A0(kld), .A1(key[40]), .B0(N165), .B1(n190), .Y(n226) );
  AOI22X1 U283 ( .A0(kld), .A1(key[41]), .B0(N164), .B1(n190), .Y(n230) );
  AOI22X1 U284 ( .A0(kld), .A1(key[42]), .B0(N163), .B1(n191), .Y(n233) );
  AOI22X1 U285 ( .A0(kld), .A1(key[43]), .B0(N162), .B1(n192), .Y(n236) );
  AOI22X1 U286 ( .A0(kld), .A1(key[44]), .B0(N161), .B1(n192), .Y(n239) );
  AOI22X1 U287 ( .A0(kld), .A1(key[45]), .B0(N160), .B1(n193), .Y(n242) );
  AOI22X1 U288 ( .A0(kld), .A1(key[46]), .B0(N159), .B1(n194), .Y(n245) );
  AOI22X1 U289 ( .A0(kld), .A1(key[47]), .B0(N158), .B1(n194), .Y(n249) );
  AOI22X1 U290 ( .A0(kld), .A1(key[48]), .B0(N157), .B1(n193), .Y(n252) );
  AOI22X1 U291 ( .A0(kld), .A1(key[49]), .B0(N156), .B1(n195), .Y(n256) );
  AOI22X1 U357 ( .A0(kld), .A1(key[50]), .B0(N155), .B1(n195), .Y(n267) );
  AOI22X1 U359 ( .A0(kld), .A1(key[51]), .B0(N154), .B1(n193), .Y(n270) );
  AOI22X1 U361 ( .A0(kld), .A1(key[52]), .B0(N153), .B1(n196), .Y(n273) );
  AOI22X1 U363 ( .A0(kld), .A1(key[53]), .B0(N152), .B1(n196), .Y(n276) );
  AOI22X1 U365 ( .A0(kld), .A1(key[54]), .B0(N151), .B1(n198), .Y(n279) );
  AOI22X1 U367 ( .A0(kld), .A1(key[55]), .B0(N150), .B1(n197), .Y(n283) );
  AOI22X1 U369 ( .A0(kld), .A1(key[56]), .B0(N149), .B1(n197), .Y(n286) );
  AOI22X1 U371 ( .A0(kld), .A1(key[57]), .B0(N148), .B1(n194), .Y(n290) );
  AOI22X1 U373 ( .A0(kld), .A1(key[58]), .B0(N147), .B1(n198), .Y(n293) );
  AOI22X1 U375 ( .A0(kld), .A1(key[59]), .B0(N146), .B1(n198), .Y(n296) );
  AOI22X1 U377 ( .A0(kld), .A1(key[60]), .B0(N145), .B1(n193), .Y(n299) );
  AOI22X1 U379 ( .A0(kld), .A1(key[61]), .B0(N144), .B1(n199), .Y(n302) );
  AOI22X1 U381 ( .A0(kld), .A1(key[62]), .B0(N143), .B1(n199), .Y(n305) );
  AOI22X1 U383 ( .A0(kld), .A1(key[63]), .B0(N142), .B1(n198), .Y(n309) );
endmodule


module aes_sbox_19 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  AOI21XL U4 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  AOI211XL U5 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  INVX1 U6 ( .A(n116), .Y(n203) );
  NOR2X1 U7 ( .A(n248), .B(n142), .Y(n357) );
  INVX1 U8 ( .A(n195), .Y(n142) );
  NAND2X1 U9 ( .A(n194), .B(n274), .Y(n344) );
  INVX1 U10 ( .A(n324), .Y(n265) );
  AOI31XL U11 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI21XL U12 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  AOI2BB2XL U13 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  NAND2XL U14 ( .A(n235), .B(n265), .Y(n338) );
  INVXL U15 ( .A(n257), .Y(n289) );
  NOR2XL U16 ( .A(n224), .B(n326), .Y(n257) );
  NAND2XL U17 ( .A(n109), .B(n78), .Y(n158) );
  AOI22XL U18 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NAND2XL U19 ( .A(n140), .B(n20), .Y(n151) );
  NOR2XL U20 ( .A(n181), .B(n95), .Y(n174) );
  NOR2X1 U21 ( .A(n293), .B(n323), .Y(n150) );
  NOR2X1 U22 ( .A(a[1]), .B(n293), .Y(n318) );
  NAND2XL U23 ( .A(a[1]), .B(n293), .Y(n82) );
  NOR2XL U24 ( .A(n324), .B(n131), .Y(n262) );
  INVXL U25 ( .A(n352), .Y(n141) );
  INVXL U26 ( .A(n267), .Y(n333) );
  NOR2X1 U27 ( .A(a[1]), .B(n103), .Y(n331) );
  NOR2XL U28 ( .A(a[1]), .B(n242), .Y(n186) );
  NOR2X4 U29 ( .A(n264), .B(n197), .Y(n350) );
  NAND2X1 U30 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI211XL U31 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  OR4X2 U32 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U33 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI211XL U34 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  AOI31XL U35 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI31XL U36 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI211XL U37 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U38 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  OAI211XL U39 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U40 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U41 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI31XL U42 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI31XL U43 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI31XL U44 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  OAI22XL U45 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  OAI211XL U46 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI211XL U47 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI22XL U48 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  AOI211XL U49 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI31XL U50 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U51 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U52 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI211XL U53 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OAI211XL U54 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI211XL U55 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI31XL U56 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI22XL U57 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI22XL U58 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI31XL U59 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  NAND2XL U60 ( .A(n296), .B(n101), .Y(n94) );
  OAI211XL U61 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  AOI211XL U62 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  INVXL U63 ( .A(n101), .Y(n254) );
  AOI31XL U64 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  OAI211XL U65 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U66 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  AOI211XL U67 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U68 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U69 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI22XL U70 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI22XL U71 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  AOI31XL U72 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI31XL U73 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI22XL U74 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI211XL U75 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  OAI211XL U76 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  NOR2XL U77 ( .A(n150), .B(n331), .Y(n130) );
  AOI31XL U78 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  NOR2XL U79 ( .A(n224), .B(n150), .Y(n116) );
  AOI22XL U80 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  AOI211XL U81 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  NAND2XL U82 ( .A(n235), .B(n274), .Y(n184) );
  AOI221XL U83 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  INVXL U84 ( .A(n150), .Y(n310) );
  AOI211XL U85 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI22XL U86 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI22XL U87 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI211XL U88 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI2BB2XL U89 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U90 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI211XL U91 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI22XL U92 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI22XL U93 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI22XL U94 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI211XL U95 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  INVXL U96 ( .A(n152), .Y(n222) );
  AOI31XL U97 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI22XL U98 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  OAI22XL U99 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI22XL U100 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI211XL U101 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI22XL U102 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI2BB2XL U103 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI211XL U104 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI2BB2XL U105 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI22XL U106 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  NAND2XL U107 ( .A(n265), .B(n348), .Y(n247) );
  AOI211XL U108 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  INVXL U109 ( .A(n312), .Y(n313) );
  NOR2XL U110 ( .A(n293), .B(n292), .Y(n294) );
  NAND2XL U111 ( .A(n103), .B(n253), .Y(n305) );
  NAND2XL U112 ( .A(n352), .B(n351), .Y(n358) );
  AOI22XL U113 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  NOR2XL U114 ( .A(n209), .B(n233), .Y(n256) );
  AOI211XL U115 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI22XL U116 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  AOI22XL U117 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI2BB2XL U118 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  OAI22XL U119 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI22XL U120 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI22XL U121 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  AOI22XL U122 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  NAND2XL U123 ( .A(n109), .B(n242), .Y(n135) );
  AOI22XL U124 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  OAI2BB1XL U125 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  NOR2XL U126 ( .A(n161), .B(n309), .Y(n162) );
  AOI22XL U127 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  INVXL U128 ( .A(n82), .Y(n172) );
  AOI32XL U129 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  AOI22XL U130 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  INVXL U131 ( .A(n180), .Y(n183) );
  AOI211XL U132 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  OAI22XL U133 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  NAND3XL U134 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  OAI211XL U135 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U136 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI2BB2XL U137 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  AOI22XL U138 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  AOI22XL U139 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  NAND2XL U140 ( .A(n311), .B(n196), .Y(n40) );
  AOI211XL U141 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  AOI22XL U142 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  AND2X2 U143 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U144 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  OAI22XL U145 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI22XL U146 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  AOI22XL U147 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  AOI22XL U148 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  NOR3XL U149 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  NOR3XL U150 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI22XL U151 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  AOI2BB2XL U152 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI31XL U153 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI22XL U154 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AOI22XL U155 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  NOR2XL U156 ( .A(n268), .B(n354), .Y(n13) );
  OAI22XL U157 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  NOR2XL U158 ( .A(n181), .B(n269), .Y(n315) );
  AOI22XL U159 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  NAND2XL U160 ( .A(n350), .B(n245), .Y(n180) );
  AOI22XL U161 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  INVXL U162 ( .A(n131), .Y(n351) );
  NOR2XL U163 ( .A(n37), .B(n145), .Y(n99) );
  NOR2XL U164 ( .A(n293), .B(n226), .Y(n39) );
  AOI22XL U165 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AOI22XL U166 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  AOI22XL U167 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI22XL U168 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  AOI22XL U169 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  NAND2XL U170 ( .A(n311), .B(n236), .Y(n346) );
  AOI22XL U171 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  NOR2XL U172 ( .A(n233), .B(n331), .Y(n108) );
  NOR2XL U173 ( .A(a[1]), .B(n329), .Y(n269) );
  NAND2XL U174 ( .A(n306), .B(n267), .Y(n61) );
  AOI22XL U175 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NAND3XL U176 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  NAND2XL U177 ( .A(n311), .B(n303), .Y(n38) );
  AOI22XL U178 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  NAND2XL U179 ( .A(n329), .B(n323), .Y(n245) );
  NAND2XL U180 ( .A(n107), .B(n348), .Y(n175) );
  AOI22XL U181 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NOR2XL U182 ( .A(n37), .B(a[1]), .Y(n195) );
  AOI22XL U183 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  NOR2XL U184 ( .A(n187), .B(n186), .Y(n290) );
  NOR2XL U185 ( .A(a[1]), .B(n249), .Y(n131) );
  NAND3XL U186 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  AOI22XL U187 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  INVXL U188 ( .A(n297), .Y(n284) );
  INVXL U189 ( .A(n332), .Y(n234) );
  NAND2XL U190 ( .A(a[1]), .B(n261), .Y(n303) );
  NAND2XL U191 ( .A(n328), .B(n311), .Y(n353) );
  INVXL U192 ( .A(n197), .Y(n185) );
  NAND3XL U193 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  NAND2XL U194 ( .A(n264), .B(n275), .Y(n252) );
  INVXL U195 ( .A(n274), .Y(n251) );
  AOI22XL U196 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  AOI22XL U197 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U198 ( .A(a[1]), .B(n198), .Y(n160) );
  NOR2XL U199 ( .A(n264), .B(n273), .Y(n330) );
  NOR2XL U200 ( .A(a[3]), .B(a[1]), .Y(n225) );
  NAND2XL U201 ( .A(a[3]), .B(a[1]), .Y(n20) );
  NAND2XL U202 ( .A(a[4]), .B(a[1]), .Y(n274) );
  INVX2 U203 ( .A(a[7]), .Y(n264) );
  CLKINVX3 U204 ( .A(n266), .Y(n329) );
  NAND2X2 U205 ( .A(a[4]), .B(n31), .Y(n266) );
  OAI21X1 U206 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U207 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U208 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U209 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U210 ( .A(a[5]), .Y(n275) );
  NOR2X2 U211 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U212 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U213 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U214 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U215 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U216 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U217 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U218 ( .A(n233), .Y(n359) );
  NAND2X2 U219 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U220 ( .A(n349), .Y(n288) );
  NOR2X4 U221 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U222 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U223 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U224 ( .A(n347), .Y(n1) );
  CLKINVX3 U225 ( .A(a[2]), .Y(n273) );
  OAI21X1 U226 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U227 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U228 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U229 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U230 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U231 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31X4 U232 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  CLKINVX3 U233 ( .A(n309), .Y(n345) );
  NAND2X2 U234 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U235 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U236 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U237 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U238 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U239 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U240 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U241 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U242 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U243 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U244 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U245 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U246 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U247 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U248 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U249 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U250 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U251 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U252 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U253 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U254 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U255 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U256 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U257 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U258 ( .A(a[1]), .Y(n323) );
  NAND2X1 U259 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U260 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U261 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U262 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U263 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U264 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U265 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U266 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U267 ( .A(n242), .Y(n249) );
  OAI21XL U268 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U269 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U270 ( .A(n192), .Y(n205) );
  INVX1 U271 ( .A(n66), .Y(n111) );
  NOR2X1 U272 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U273 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U274 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U275 ( .A(a[6]), .B(a[0]), .Y(n360) );
  INVX1 U276 ( .A(a[6]), .Y(n16) );
  NOR2X1 U277 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U278 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U279 ( .A(n261), .Y(n307) );
  INVX1 U280 ( .A(n20), .Y(n326) );
  NAND2X1 U281 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U282 ( .A(n187), .Y(n196) );
  INVX1 U283 ( .A(n350), .Y(n335) );
  NAND2X1 U284 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U285 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U286 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U287 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U288 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U289 ( .A(n103), .Y(n37) );
  NOR2X1 U290 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U291 ( .A(n311), .Y(n268) );
  INVX1 U292 ( .A(n293), .Y(n209) );
  NOR2X1 U293 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U294 ( .A(n224), .Y(n235) );
  NAND2X1 U295 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U296 ( .AN(n140), .B(n181), .Y(n92) );
  NAND2X1 U297 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U298 ( .A(n226), .Y(n253) );
  NAND2X1 U299 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U300 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U301 ( .A(n1), .Y(n301) );
  NAND2X1 U302 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U303 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U304 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U305 ( .A(n89), .Y(n340) );
  AOI211X1 U306 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U307 ( .A(n327), .Y(n248) );
  INVX1 U308 ( .A(n181), .Y(n109) );
  INVX1 U309 ( .A(n225), .Y(n302) );
  NAND2X1 U310 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U311 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U312 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U313 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U314 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U315 ( .A(n270), .Y(n107) );
  INVX1 U316 ( .A(n306), .Y(n145) );
  NAND4X1 U317 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U318 ( .A(n210), .Y(n236) );
  INVX1 U319 ( .A(n331), .Y(n78) );
  INVX1 U320 ( .A(n328), .Y(n314) );
  OAI21XL U321 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U322 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U323 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U324 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_4 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  NAND2XL U4 ( .A(n235), .B(n265), .Y(n338) );
  INVXL U5 ( .A(n116), .Y(n203) );
  INVX1 U6 ( .A(n324), .Y(n265) );
  INVXL U7 ( .A(n192), .Y(n205) );
  INVX2 U8 ( .A(a[4]), .Y(n198) );
  AOI31XL U9 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI21XL U10 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  AOI2BB2XL U11 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI211XL U12 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI211XL U13 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  INVXL U14 ( .A(n257), .Y(n289) );
  NOR2XL U15 ( .A(n224), .B(n326), .Y(n257) );
  NOR2XL U16 ( .A(n248), .B(n142), .Y(n357) );
  AOI22XL U17 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  AOI32XL U18 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(n193) );
  NAND2XL U19 ( .A(n109), .B(n78), .Y(n158) );
  NOR2XL U20 ( .A(n181), .B(n95), .Y(n174) );
  NOR2X1 U21 ( .A(n293), .B(n323), .Y(n150) );
  NAND2XL U22 ( .A(n140), .B(n20), .Y(n151) );
  NAND2XL U23 ( .A(a[1]), .B(n293), .Y(n82) );
  NOR2XL U24 ( .A(n324), .B(n131), .Y(n262) );
  NOR2X1 U25 ( .A(a[1]), .B(n293), .Y(n318) );
  NAND2XL U26 ( .A(n194), .B(n274), .Y(n344) );
  NAND2XL U27 ( .A(n329), .B(n323), .Y(n245) );
  NAND2XL U28 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U29 ( .A(a[1]), .B(n103), .Y(n331) );
  CLKINVX3 U30 ( .A(n266), .Y(n329) );
  INVXL U31 ( .A(n267), .Y(n333) );
  INVXL U32 ( .A(n352), .Y(n141) );
  NOR2XL U33 ( .A(n323), .B(n266), .Y(n187) );
  NOR2X4 U34 ( .A(n264), .B(n197), .Y(n350) );
  NOR2XL U35 ( .A(a[1]), .B(n242), .Y(n186) );
  NAND2X1 U36 ( .A(a[1]), .B(n31), .Y(n352) );
  INVX1 U37 ( .A(n89), .Y(n340) );
  AOI31XL U38 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  OR4X2 U39 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U40 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U41 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  AOI211XL U42 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI31XL U43 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI31XL U44 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U45 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI31XL U46 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31XL U47 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U48 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  OAI211XL U49 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI211XL U50 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI211XL U51 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI211XL U52 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U53 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI21X1 U54 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  AOI211XL U55 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI31XL U56 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  AOI31XL U57 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  OAI211XL U58 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI22XL U59 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI22XL U60 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  AOI211XL U61 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI31XL U62 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI31XL U63 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  OAI22XL U64 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI22XL U65 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  OAI211XL U66 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI31XL U67 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  INVXL U68 ( .A(n101), .Y(n254) );
  AOI31XL U69 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  AOI211XL U70 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  NAND2XL U71 ( .A(n296), .B(n101), .Y(n94) );
  AOI31XL U72 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  OAI211XL U73 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  AOI211XL U74 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U75 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U76 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI22XL U77 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U78 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  OAI211XL U79 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U80 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI31XL U81 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  INVXL U82 ( .A(n150), .Y(n310) );
  AOI211XL U83 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  AOI22XL U84 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI211XL U85 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI22XL U86 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  NOR2XL U87 ( .A(n150), .B(n331), .Y(n130) );
  AOI221XL U88 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI31XL U89 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  NAND2XL U90 ( .A(n235), .B(n274), .Y(n184) );
  NOR2XL U91 ( .A(n224), .B(n150), .Y(n116) );
  AOI31XL U92 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  AOI22XL U93 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  OAI211XL U94 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  AOI211XL U95 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI31XL U96 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  INVXL U97 ( .A(n152), .Y(n222) );
  AOI211XL U98 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI2BB2XL U99 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  NAND2XL U100 ( .A(n265), .B(n348), .Y(n247) );
  AOI22XL U101 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI211XL U102 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI22XL U103 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI22XL U104 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI22XL U105 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI2BB2XL U106 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U107 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI211XL U108 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI22XL U109 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI211XL U110 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI22XL U111 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI211XL U112 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI2BB2XL U113 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI22XL U114 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI22XL U115 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  OAI22XL U116 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI22XL U117 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  NAND2XL U118 ( .A(n352), .B(n351), .Y(n358) );
  AOI22XL U119 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  INVXL U120 ( .A(n312), .Y(n313) );
  NAND2XL U121 ( .A(n103), .B(n253), .Y(n305) );
  NOR2XL U122 ( .A(n293), .B(n292), .Y(n294) );
  OAI211XL U123 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U124 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI22XL U125 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  OAI22XL U126 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  NAND3XL U127 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  AOI22XL U128 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  AOI22XL U129 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI211XL U130 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI22XL U131 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  AOI22XL U132 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI2BB2XL U133 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  OAI22XL U134 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI22XL U135 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  AOI22XL U136 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  AOI22XL U137 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  AOI2BB2XL U138 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  NOR2XL U139 ( .A(n209), .B(n233), .Y(n256) );
  OAI2BB1XL U140 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  AOI22XL U141 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  AOI22XL U142 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  AOI211XL U143 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  INVXL U144 ( .A(n180), .Y(n183) );
  INVXL U145 ( .A(n82), .Y(n172) );
  NOR2XL U146 ( .A(n161), .B(n309), .Y(n162) );
  AOI22XL U147 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  NAND2XL U148 ( .A(n109), .B(n242), .Y(n135) );
  OAI22XL U149 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  NAND2XL U150 ( .A(n350), .B(n245), .Y(n180) );
  AOI22XL U151 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  AOI22XL U152 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI22XL U153 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  AOI22XL U154 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  AOI2BB2XL U155 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U156 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  AOI22XL U157 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  NOR2XL U158 ( .A(n181), .B(n269), .Y(n315) );
  NOR2XL U159 ( .A(n293), .B(n226), .Y(n39) );
  NAND2XL U160 ( .A(n311), .B(n196), .Y(n40) );
  NOR3XL U161 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI22XL U162 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  AOI211XL U163 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  AOI31XL U164 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  NOR3XL U165 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  NOR2XL U166 ( .A(n37), .B(n145), .Y(n99) );
  AOI22XL U167 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  OAI22XL U168 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U169 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AOI22XL U170 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  NOR2XL U171 ( .A(n268), .B(n354), .Y(n13) );
  INVXL U172 ( .A(n131), .Y(n351) );
  AOI22XL U173 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  AOI22XL U174 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AOI22XL U175 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  AOI22XL U176 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  NAND2XL U177 ( .A(n311), .B(n236), .Y(n346) );
  AND2X2 U178 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U179 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  NAND3XL U180 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NAND2XL U181 ( .A(n306), .B(n267), .Y(n61) );
  AOI22XL U182 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NAND2XL U183 ( .A(n107), .B(n348), .Y(n175) );
  NAND3XL U184 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  NAND2XL U185 ( .A(n311), .B(n303), .Y(n38) );
  NOR2XL U186 ( .A(n37), .B(a[1]), .Y(n195) );
  NOR2XL U187 ( .A(n187), .B(n186), .Y(n290) );
  NOR2XL U188 ( .A(a[1]), .B(n249), .Y(n131) );
  AOI22XL U189 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  AOI22XL U190 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  AOI22XL U191 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NOR2XL U192 ( .A(a[1]), .B(n329), .Y(n269) );
  AOI22XL U193 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  AOI22XL U194 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  NOR2XL U195 ( .A(n233), .B(n331), .Y(n108) );
  INVXL U196 ( .A(n297), .Y(n284) );
  INVXL U197 ( .A(n332), .Y(n234) );
  NAND2XL U198 ( .A(n328), .B(n311), .Y(n353) );
  NAND2XL U199 ( .A(a[1]), .B(n261), .Y(n303) );
  INVXL U200 ( .A(n197), .Y(n185) );
  NAND3XL U201 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  NOR2XL U202 ( .A(n264), .B(n273), .Y(n330) );
  AOI22XL U203 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U204 ( .A(a[1]), .B(n198), .Y(n160) );
  NAND2XL U205 ( .A(n264), .B(n275), .Y(n252) );
  INVXL U206 ( .A(n274), .Y(n251) );
  AOI22XL U207 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  INVX2 U208 ( .A(a[7]), .Y(n264) );
  NAND2XL U209 ( .A(a[4]), .B(a[1]), .Y(n274) );
  NAND2XL U210 ( .A(a[3]), .B(a[1]), .Y(n20) );
  NOR2XL U211 ( .A(a[3]), .B(a[1]), .Y(n225) );
  OAI21X1 U212 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U213 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  OAI21X1 U214 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U215 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U216 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U217 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U218 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U219 ( .A(a[5]), .Y(n275) );
  NOR2X2 U220 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U221 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U222 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U223 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U224 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U225 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U226 ( .A(n233), .Y(n359) );
  NAND2X2 U227 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U228 ( .A(n349), .Y(n288) );
  NOR2X4 U229 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U230 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U231 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U232 ( .A(n347), .Y(n1) );
  CLKINVX3 U233 ( .A(a[2]), .Y(n273) );
  NOR2X4 U234 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U235 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  NAND2X2 U236 ( .A(a[6]), .B(a[0]), .Y(n360) );
  CLKINVX3 U237 ( .A(n309), .Y(n345) );
  NAND2X2 U238 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U239 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U240 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U241 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U242 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U243 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U244 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U245 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U246 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U247 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U248 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U249 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U250 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U251 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U252 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U253 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U254 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U255 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U256 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U257 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U258 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  AOI21XL U259 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U260 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  NOR2X1 U261 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U262 ( .A(a[1]), .Y(n323) );
  NAND2X1 U263 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U264 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U265 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U266 ( .A(a[4]), .B(n31), .Y(n266) );
  NOR2X1 U267 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U268 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U269 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U270 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U271 ( .A(n242), .Y(n249) );
  OAI21XL U272 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U273 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U274 ( .A(n66), .Y(n111) );
  NOR2X1 U275 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U276 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U277 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  INVX1 U278 ( .A(a[6]), .Y(n16) );
  NOR2X1 U279 ( .A(a[0]), .B(n16), .Y(n125) );
  INVX1 U280 ( .A(n261), .Y(n307) );
  INVX1 U281 ( .A(n20), .Y(n326) );
  NAND2X1 U282 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U283 ( .A(n187), .Y(n196) );
  INVX1 U284 ( .A(n350), .Y(n335) );
  NAND2X1 U285 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U286 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U287 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U288 ( .A(a[3]), .B(n323), .Y(n267) );
  INVX1 U289 ( .A(n103), .Y(n37) );
  NOR2X1 U290 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U291 ( .A(n311), .Y(n268) );
  INVX1 U292 ( .A(n293), .Y(n209) );
  NOR2X1 U293 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U294 ( .A(n224), .Y(n235) );
  NAND2X1 U295 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U296 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U297 ( .A(n195), .Y(n142) );
  NAND2X1 U298 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U299 ( .A(n226), .Y(n253) );
  NAND2X1 U300 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U301 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U302 ( .A(n1), .Y(n301) );
  NAND2X1 U303 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U304 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U305 ( .A(a[6]), .B(a[0]), .Y(n89) );
  AOI211X1 U306 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U307 ( .A(n327), .Y(n248) );
  INVX1 U308 ( .A(n181), .Y(n109) );
  INVX1 U309 ( .A(n225), .Y(n302) );
  NAND2X1 U310 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U311 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U312 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U313 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U314 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U315 ( .A(n270), .Y(n107) );
  INVX1 U316 ( .A(n306), .Y(n145) );
  NAND4X1 U317 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U318 ( .A(n210), .Y(n236) );
  INVX1 U319 ( .A(n331), .Y(n78) );
  INVX1 U320 ( .A(n328), .Y(n314) );
  OAI21XL U321 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U322 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U323 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U324 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_5 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  OAI21XL U4 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  INVXL U5 ( .A(n116), .Y(n203) );
  NAND2XL U6 ( .A(n235), .B(n265), .Y(n338) );
  NAND2XL U7 ( .A(n327), .B(n266), .Y(n95) );
  INVXL U8 ( .A(n192), .Y(n205) );
  INVX2 U9 ( .A(a[4]), .Y(n198) );
  AOI31XL U10 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI2BB2XL U11 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI21XL U12 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  AOI211XL U13 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI211XL U14 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  INVXL U15 ( .A(n257), .Y(n289) );
  NOR2XL U16 ( .A(n224), .B(n326), .Y(n257) );
  AOI32XL U17 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(n193) );
  NOR2XL U18 ( .A(n248), .B(n142), .Y(n357) );
  NAND2XL U19 ( .A(n109), .B(n78), .Y(n158) );
  NOR2X1 U20 ( .A(n268), .B(n354), .Y(n13) );
  NAND2XL U21 ( .A(n140), .B(n20), .Y(n151) );
  NAND2XL U22 ( .A(a[1]), .B(n293), .Y(n82) );
  NOR2XL U23 ( .A(n181), .B(n95), .Y(n174) );
  NOR2XL U24 ( .A(n324), .B(n131), .Y(n262) );
  NOR2X1 U25 ( .A(n293), .B(n323), .Y(n150) );
  NAND2XL U26 ( .A(n194), .B(n274), .Y(n344) );
  NOR2X1 U27 ( .A(a[1]), .B(n293), .Y(n318) );
  NAND2XL U28 ( .A(n329), .B(n323), .Y(n245) );
  INVX2 U29 ( .A(n324), .Y(n265) );
  CLKINVX3 U30 ( .A(n266), .Y(n329) );
  NOR2X1 U31 ( .A(a[1]), .B(n103), .Y(n331) );
  NOR2XL U32 ( .A(n323), .B(n266), .Y(n187) );
  NOR2X4 U33 ( .A(n264), .B(n197), .Y(n350) );
  NOR2XL U34 ( .A(a[1]), .B(n242), .Y(n186) );
  INVXL U35 ( .A(n267), .Y(n333) );
  INVXL U36 ( .A(n352), .Y(n141) );
  INVX1 U37 ( .A(n89), .Y(n340) );
  NAND2X1 U38 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI31XL U39 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  OR4X2 U40 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U41 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U42 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI211XL U43 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  AOI31XL U44 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U45 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U46 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI31XL U47 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI31XL U48 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI211XL U49 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U50 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  OAI211XL U51 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI21X1 U52 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  AOI22XL U53 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI211XL U54 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI211XL U55 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI31XL U56 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  OAI22XL U57 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI31XL U58 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  OAI211XL U59 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI22XL U60 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  OAI211XL U61 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI31XL U62 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U63 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI31XL U64 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  AOI22XL U65 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI211XL U66 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI211XL U67 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI31XL U68 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  NAND2XL U69 ( .A(n296), .B(n101), .Y(n94) );
  INVXL U70 ( .A(n101), .Y(n254) );
  AOI211XL U71 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  AOI31XL U72 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  AOI22XL U73 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  OAI211XL U74 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI31XL U75 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  AOI211XL U76 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI211XL U77 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U78 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U79 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  OAI211XL U80 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  OAI211XL U81 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  INVXL U82 ( .A(n150), .Y(n310) );
  AOI22XL U83 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  AOI211XL U84 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI22XL U85 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  AOI31XL U86 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI31XL U87 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  NOR2XL U88 ( .A(n150), .B(n331), .Y(n130) );
  NAND2XL U89 ( .A(n235), .B(n274), .Y(n184) );
  AOI211XL U90 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  NOR2XL U91 ( .A(n224), .B(n150), .Y(n116) );
  AOI221XL U92 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI22XL U93 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI211XL U94 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  AOI31XL U95 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI2BB2XL U96 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U97 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI22XL U98 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI211XL U99 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI22XL U100 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI22XL U101 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  INVXL U102 ( .A(n152), .Y(n222) );
  AOI22XL U103 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI211XL U104 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  NAND2XL U105 ( .A(n265), .B(n348), .Y(n247) );
  AOI22XL U106 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI31XL U107 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI211XL U108 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI2BB2XL U109 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  OAI22XL U110 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI22XL U111 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI211XL U112 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI22XL U113 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI2BB2XL U114 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI211XL U115 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI22XL U116 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI211XL U117 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI22XL U118 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI22XL U119 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  AOI22XL U120 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  INVXL U121 ( .A(n312), .Y(n313) );
  NOR2XL U122 ( .A(n293), .B(n292), .Y(n294) );
  NAND2XL U123 ( .A(n352), .B(n351), .Y(n358) );
  AOI22XL U124 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  AOI22XL U125 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI2BB2XL U126 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  AOI2BB2XL U127 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U128 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI22XL U129 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  OAI211XL U130 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U131 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  AOI22XL U132 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  OAI2BB1XL U133 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  AOI22XL U134 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  NAND2XL U135 ( .A(n103), .B(n253), .Y(n305) );
  INVXL U136 ( .A(n82), .Y(n172) );
  INVXL U137 ( .A(n180), .Y(n183) );
  AOI211XL U138 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  OAI22XL U139 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  OAI22XL U140 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  AOI22XL U141 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  NOR2XL U142 ( .A(n161), .B(n309), .Y(n162) );
  AOI211XL U143 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  NAND2XL U144 ( .A(n109), .B(n242), .Y(n135) );
  AOI22XL U145 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  AOI22XL U146 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  AOI22XL U147 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  NOR2XL U148 ( .A(n209), .B(n233), .Y(n256) );
  NAND3XL U149 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  NOR2XL U150 ( .A(n293), .B(n226), .Y(n39) );
  AOI31XL U151 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI22XL U152 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  AOI22XL U153 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  AND2X2 U154 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U155 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  NOR2XL U156 ( .A(n181), .B(n269), .Y(n315) );
  INVXL U157 ( .A(n131), .Y(n351) );
  AOI22XL U158 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  AOI22XL U159 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI22XL U160 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  AOI2BB2XL U161 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U162 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AOI22XL U163 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  AOI22XL U164 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  NAND2XL U165 ( .A(n311), .B(n196), .Y(n40) );
  NAND2XL U166 ( .A(n350), .B(n245), .Y(n180) );
  OAI22XL U167 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U168 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AOI22XL U169 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  AOI22XL U170 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  AOI22XL U171 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  OAI22XL U172 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  NAND2XL U173 ( .A(n311), .B(n236), .Y(n346) );
  AOI22XL U174 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  NOR3XL U175 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  AOI211XL U176 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  NOR3XL U177 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  NOR2XL U178 ( .A(n37), .B(n145), .Y(n99) );
  AOI22XL U179 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  AOI22XL U180 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  AOI22XL U181 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  NOR2XL U182 ( .A(n37), .B(a[1]), .Y(n195) );
  NOR2XL U183 ( .A(a[1]), .B(n249), .Y(n131) );
  NAND3XL U184 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  AOI22XL U185 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  NOR2XL U186 ( .A(n187), .B(n186), .Y(n290) );
  NAND2XL U187 ( .A(n311), .B(n303), .Y(n38) );
  AOI22XL U188 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  NAND2XL U189 ( .A(n306), .B(n267), .Y(n61) );
  AOI22XL U190 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NAND2XL U191 ( .A(n107), .B(n348), .Y(n175) );
  NAND3XL U192 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NOR2XL U193 ( .A(n233), .B(n331), .Y(n108) );
  AOI22XL U194 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NOR2XL U195 ( .A(a[1]), .B(n329), .Y(n269) );
  NAND2XL U196 ( .A(a[1]), .B(n261), .Y(n303) );
  INVXL U197 ( .A(n297), .Y(n284) );
  NAND3XL U198 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  INVXL U199 ( .A(n332), .Y(n234) );
  INVXL U200 ( .A(n197), .Y(n185) );
  NAND2XL U201 ( .A(n328), .B(n311), .Y(n353) );
  AOI22XL U202 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  NOR2XL U203 ( .A(a[1]), .B(n198), .Y(n160) );
  NAND2XL U204 ( .A(n264), .B(n275), .Y(n252) );
  NOR2XL U205 ( .A(n264), .B(n273), .Y(n330) );
  INVXL U206 ( .A(n274), .Y(n251) );
  AOI22XL U207 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NAND2XL U208 ( .A(a[3]), .B(a[1]), .Y(n20) );
  INVX2 U209 ( .A(a[7]), .Y(n264) );
  INVX1 U210 ( .A(a[6]), .Y(n16) );
  NOR2XL U211 ( .A(a[3]), .B(a[1]), .Y(n225) );
  NAND2XL U212 ( .A(a[4]), .B(a[1]), .Y(n274) );
  OAI21X1 U213 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  OAI21X1 U214 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U215 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U216 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U217 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U218 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U219 ( .A(a[5]), .Y(n275) );
  NOR2X2 U220 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U221 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U222 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U223 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U224 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U225 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U226 ( .A(n233), .Y(n359) );
  NAND2X2 U227 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U228 ( .A(n349), .Y(n288) );
  NOR2X4 U229 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U230 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U231 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U232 ( .A(n347), .Y(n1) );
  CLKINVX3 U233 ( .A(a[2]), .Y(n273) );
  NOR2X4 U234 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U235 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  NAND2X2 U236 ( .A(a[6]), .B(a[0]), .Y(n360) );
  CLKINVX3 U237 ( .A(n309), .Y(n345) );
  NAND2X2 U238 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U239 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U240 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U241 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U242 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U243 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U244 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U245 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U246 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U247 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U248 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U249 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U250 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U251 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U252 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U253 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U254 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U255 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U256 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U257 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U258 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  AOI21XL U259 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U260 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  NOR2X1 U261 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U262 ( .A(a[1]), .Y(n323) );
  NAND2X1 U263 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U264 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U265 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U266 ( .A(a[4]), .B(n31), .Y(n266) );
  NOR2X1 U267 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U268 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U269 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U270 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U271 ( .A(n242), .Y(n249) );
  OAI21XL U272 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U273 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U274 ( .A(n66), .Y(n111) );
  NOR2X1 U275 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U276 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U277 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NOR2X1 U278 ( .A(a[0]), .B(n16), .Y(n125) );
  INVX1 U279 ( .A(n261), .Y(n307) );
  INVX1 U280 ( .A(n20), .Y(n326) );
  NAND2X1 U281 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U282 ( .A(n187), .Y(n196) );
  INVX1 U283 ( .A(n350), .Y(n335) );
  NAND2X1 U284 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U285 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U286 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U287 ( .A(a[3]), .B(n323), .Y(n267) );
  INVX1 U288 ( .A(n103), .Y(n37) );
  NOR2X1 U289 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U290 ( .A(n311), .Y(n268) );
  AOI22X1 U291 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  INVX1 U292 ( .A(n293), .Y(n209) );
  NOR2X1 U293 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U294 ( .A(n224), .Y(n235) );
  NAND2X1 U295 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U296 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U297 ( .A(n195), .Y(n142) );
  NAND2X1 U298 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U299 ( .A(n226), .Y(n253) );
  NAND2X1 U300 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U301 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U302 ( .A(n1), .Y(n301) );
  NAND2X1 U303 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U304 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U305 ( .A(a[6]), .B(a[0]), .Y(n89) );
  AOI211X1 U306 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U307 ( .A(n327), .Y(n248) );
  INVX1 U308 ( .A(n181), .Y(n109) );
  INVX1 U309 ( .A(n225), .Y(n302) );
  NAND2X1 U310 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U311 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U312 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U313 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U314 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U315 ( .A(n270), .Y(n107) );
  INVX1 U316 ( .A(n306), .Y(n145) );
  NAND4X1 U317 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U318 ( .A(n210), .Y(n236) );
  INVX1 U319 ( .A(n331), .Y(n78) );
  INVX1 U320 ( .A(n328), .Y(n314) );
  OAI21XL U321 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U322 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U323 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U324 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_6 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  OAI21XL U4 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  NOR2XL U5 ( .A(n268), .B(n354), .Y(n13) );
  INVX1 U6 ( .A(n324), .Y(n265) );
  AOI31XL U7 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI21XL U8 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  AOI2BB2XL U9 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI211XL U10 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  AOI211XL U11 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  INVXL U12 ( .A(n257), .Y(n289) );
  NAND2XL U13 ( .A(n235), .B(n265), .Y(n338) );
  NOR2XL U14 ( .A(n224), .B(n326), .Y(n257) );
  INVXL U15 ( .A(n150), .Y(n310) );
  NAND2XL U16 ( .A(n109), .B(n78), .Y(n158) );
  AOI32XL U17 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(n193) );
  AOI22XL U18 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NOR2XL U19 ( .A(n248), .B(n142), .Y(n357) );
  NOR2XL U20 ( .A(n324), .B(n131), .Y(n262) );
  NAND2XL U21 ( .A(n140), .B(n20), .Y(n151) );
  NAND2XL U22 ( .A(n194), .B(n274), .Y(n344) );
  NOR2XL U23 ( .A(n181), .B(n95), .Y(n174) );
  NOR2X1 U24 ( .A(n293), .B(n323), .Y(n150) );
  NOR2X1 U25 ( .A(a[1]), .B(n293), .Y(n318) );
  NAND2XL U26 ( .A(a[1]), .B(n293), .Y(n82) );
  NAND2XL U27 ( .A(n327), .B(n266), .Y(n95) );
  NAND2XL U28 ( .A(n329), .B(n323), .Y(n245) );
  CLKINVX3 U29 ( .A(n266), .Y(n329) );
  INVXL U30 ( .A(n352), .Y(n141) );
  NOR2XL U31 ( .A(a[1]), .B(n242), .Y(n186) );
  NOR2XL U32 ( .A(n323), .B(n266), .Y(n187) );
  NOR2X1 U33 ( .A(a[1]), .B(n103), .Y(n331) );
  INVXL U34 ( .A(n267), .Y(n333) );
  NOR2X4 U35 ( .A(n264), .B(n197), .Y(n350) );
  NAND2X1 U36 ( .A(a[1]), .B(n31), .Y(n352) );
  INVX1 U37 ( .A(n89), .Y(n340) );
  OR4X2 U38 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U39 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI31XL U40 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI211XL U41 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U42 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  AOI31XL U43 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31XL U44 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI211XL U45 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U46 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  OAI211XL U47 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U48 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI31XL U49 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U50 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI211XL U51 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI31XL U52 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI22XL U53 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  OAI211XL U54 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI211XL U55 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI211XL U56 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI22XL U57 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI22XL U58 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI21X1 U59 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  AOI211XL U60 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI211XL U61 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI31XL U62 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI31XL U63 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  OAI22XL U64 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI31XL U65 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  OAI211XL U66 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI31XL U67 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  NAND2XL U68 ( .A(n296), .B(n101), .Y(n94) );
  AOI31XL U69 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  INVXL U70 ( .A(n101), .Y(n254) );
  AOI31XL U71 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  OAI211XL U72 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U73 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U74 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U75 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  AOI211XL U76 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  AOI211XL U77 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI22XL U78 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  OAI211XL U79 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  AOI22XL U80 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  AOI211XL U81 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI22XL U82 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  NOR2XL U83 ( .A(n224), .B(n150), .Y(n116) );
  AOI211XL U84 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI221XL U85 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI31XL U86 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  AOI31XL U87 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI22XL U88 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  AOI31XL U89 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  OAI211XL U90 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  NOR2XL U91 ( .A(n150), .B(n331), .Y(n130) );
  AOI211XL U92 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  NAND2XL U93 ( .A(n235), .B(n274), .Y(n184) );
  AOI211XL U94 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI22XL U95 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI22XL U96 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI22XL U97 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI211XL U98 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  NAND2XL U99 ( .A(n265), .B(n348), .Y(n247) );
  AOI2BB2XL U100 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  OAI22XL U101 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI22XL U102 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI22XL U103 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI2BB2XL U104 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI2BB2XL U105 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI211XL U106 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI211XL U107 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI31XL U108 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI22XL U109 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI22XL U110 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI22XL U111 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI211XL U112 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI22XL U113 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI22XL U114 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI211XL U115 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  INVXL U116 ( .A(n152), .Y(n222) );
  INVXL U117 ( .A(n82), .Y(n172) );
  INVXL U118 ( .A(n180), .Y(n183) );
  AOI22XL U119 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  AOI211XL U120 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  AOI22XL U121 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  OAI22XL U122 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  OAI2BB1XL U123 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  NAND3XL U124 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  AOI211XL U125 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI22XL U126 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  NAND2XL U127 ( .A(n109), .B(n242), .Y(n135) );
  AOI22XL U128 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  OAI22XL U129 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI22XL U130 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  AOI22XL U131 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI2BB2XL U132 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U133 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  NOR2XL U134 ( .A(n161), .B(n309), .Y(n162) );
  AOI22XL U135 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  AOI22XL U136 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  AOI22XL U137 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  NAND2XL U138 ( .A(n103), .B(n253), .Y(n305) );
  AOI22XL U139 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  AOI22XL U140 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  INVXL U141 ( .A(n312), .Y(n313) );
  OAI211XL U142 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U143 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  NOR2XL U144 ( .A(n293), .B(n292), .Y(n294) );
  AOI2BB2XL U145 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  NOR2XL U146 ( .A(n209), .B(n233), .Y(n256) );
  NAND2XL U147 ( .A(n352), .B(n351), .Y(n358) );
  AOI22XL U148 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  AOI22XL U149 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  AOI22XL U150 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  NOR2XL U151 ( .A(n293), .B(n226), .Y(n39) );
  AOI22XL U152 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  AOI31XL U153 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI22XL U154 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  AOI211XL U155 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  NAND2XL U156 ( .A(n311), .B(n236), .Y(n346) );
  NAND2XL U157 ( .A(n311), .B(n196), .Y(n40) );
  AOI22XL U158 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  NAND2XL U159 ( .A(n350), .B(n245), .Y(n180) );
  AOI22XL U160 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  NOR3XL U161 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  AOI22XL U162 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  INVXL U163 ( .A(n131), .Y(n351) );
  NOR2XL U164 ( .A(n181), .B(n269), .Y(n315) );
  AOI2BB2XL U165 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U166 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI22XL U167 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  NOR3XL U168 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI22XL U169 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  AOI22XL U170 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  OAI22XL U171 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI22XL U172 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  NOR2XL U173 ( .A(n37), .B(n145), .Y(n99) );
  AND2X2 U174 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U175 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  OAI22XL U176 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U177 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AOI22XL U178 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  AOI22XL U179 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NOR2XL U180 ( .A(n37), .B(a[1]), .Y(n195) );
  NOR2XL U181 ( .A(a[1]), .B(n329), .Y(n269) );
  NAND3XL U182 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NAND2XL U183 ( .A(n311), .B(n303), .Y(n38) );
  NAND2XL U184 ( .A(n107), .B(n348), .Y(n175) );
  NOR2XL U185 ( .A(a[1]), .B(n249), .Y(n131) );
  NAND2XL U186 ( .A(n306), .B(n267), .Y(n61) );
  AOI22XL U187 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  NOR2XL U188 ( .A(n233), .B(n331), .Y(n108) );
  NOR2XL U189 ( .A(n187), .B(n186), .Y(n290) );
  AOI22XL U190 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  AOI22XL U191 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  AOI22XL U192 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  NAND3XL U193 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  NAND2XL U194 ( .A(a[1]), .B(n261), .Y(n303) );
  INVXL U195 ( .A(n297), .Y(n284) );
  NAND2XL U196 ( .A(n328), .B(n311), .Y(n353) );
  INVXL U197 ( .A(n197), .Y(n185) );
  INVXL U198 ( .A(n332), .Y(n234) );
  NAND3XL U199 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  NAND2XL U200 ( .A(n264), .B(n275), .Y(n252) );
  NOR2XL U201 ( .A(n264), .B(n273), .Y(n330) );
  INVXL U202 ( .A(n274), .Y(n251) );
  AOI22XL U203 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  NOR2XL U204 ( .A(a[1]), .B(n198), .Y(n160) );
  AOI22XL U205 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U206 ( .A(a[3]), .B(a[1]), .Y(n225) );
  NAND2XL U207 ( .A(a[4]), .B(a[1]), .Y(n274) );
  NAND2XL U208 ( .A(a[3]), .B(a[1]), .Y(n20) );
  INVX2 U209 ( .A(a[7]), .Y(n264) );
  OAI21X1 U210 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  OAI21X1 U211 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U212 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U213 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U214 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U215 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U216 ( .A(a[5]), .Y(n275) );
  NOR2X2 U217 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U218 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U219 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U220 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U221 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U222 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U223 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U224 ( .A(n233), .Y(n359) );
  NAND2X2 U225 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U226 ( .A(n349), .Y(n288) );
  NOR2X4 U227 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U228 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U229 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U230 ( .A(n347), .Y(n1) );
  CLKINVX3 U231 ( .A(a[2]), .Y(n273) );
  NOR2X4 U232 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U233 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  NAND2X2 U234 ( .A(a[6]), .B(a[0]), .Y(n360) );
  CLKINVX3 U235 ( .A(n309), .Y(n345) );
  NAND2X2 U236 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U237 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U238 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U239 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U240 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U241 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U242 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U243 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U244 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U245 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U246 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U247 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U248 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U249 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U250 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U251 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U252 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U253 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U254 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U255 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U256 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  AOI21XL U257 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U258 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  NOR2X1 U259 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U260 ( .A(a[1]), .Y(n323) );
  NAND2X1 U261 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U262 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U263 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U264 ( .A(a[4]), .B(n31), .Y(n266) );
  NOR2X1 U265 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U266 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U267 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U268 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U269 ( .A(n242), .Y(n249) );
  OAI21XL U270 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U271 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U272 ( .A(n192), .Y(n205) );
  INVX1 U273 ( .A(n66), .Y(n111) );
  NOR2X1 U274 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U275 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U276 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  INVX1 U277 ( .A(a[6]), .Y(n16) );
  NOR2X1 U278 ( .A(a[0]), .B(n16), .Y(n125) );
  INVX1 U279 ( .A(n261), .Y(n307) );
  INVX1 U280 ( .A(n20), .Y(n326) );
  NAND2X1 U281 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U282 ( .A(n187), .Y(n196) );
  INVX1 U283 ( .A(n350), .Y(n335) );
  NAND2X1 U284 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U285 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U286 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U287 ( .A(a[3]), .B(n323), .Y(n267) );
  INVX1 U288 ( .A(n103), .Y(n37) );
  NOR2X1 U289 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U290 ( .A(n311), .Y(n268) );
  INVX1 U291 ( .A(n293), .Y(n209) );
  NOR2X1 U292 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U293 ( .A(n224), .Y(n235) );
  NAND2X1 U294 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U295 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U296 ( .A(n195), .Y(n142) );
  NAND2X1 U297 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U298 ( .A(n226), .Y(n253) );
  NAND2X1 U299 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U300 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U301 ( .A(n1), .Y(n301) );
  NAND2X1 U302 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U303 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U304 ( .A(a[6]), .B(a[0]), .Y(n89) );
  AOI211X1 U305 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U306 ( .A(n327), .Y(n248) );
  INVX1 U307 ( .A(n181), .Y(n109) );
  INVX1 U308 ( .A(n225), .Y(n302) );
  NAND2X1 U309 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U310 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U311 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U312 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U313 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U314 ( .A(n270), .Y(n107) );
  INVX1 U315 ( .A(n306), .Y(n145) );
  NAND4X1 U316 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U317 ( .A(n210), .Y(n236) );
  INVX1 U318 ( .A(n331), .Y(n78) );
  INVX1 U319 ( .A(n328), .Y(n314) );
  OAI21XL U320 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U321 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U322 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U323 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U324 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U325 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U326 ( .A(n186), .Y(n194) );
  NAND2X1 U327 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U328 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U329 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U330 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U331 ( .A(n72), .Y(n204) );
  OAI21XL U332 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U333 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U334 ( .A(n125), .Y(n319) );
  NAND2X1 U335 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U336 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U337 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U338 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U339 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U340 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U341 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U342 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U343 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U344 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U345 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U346 ( .A(n116), .Y(n203) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_7 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  OAI21XL U4 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  INVXL U5 ( .A(n116), .Y(n203) );
  INVX1 U6 ( .A(n324), .Y(n265) );
  INVXL U7 ( .A(n192), .Y(n205) );
  CLKINVX3 U8 ( .A(n266), .Y(n329) );
  AOI31XL U9 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI211XL U10 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI2BB2XL U11 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI21XL U12 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  AOI211XL U13 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  NAND2XL U14 ( .A(n235), .B(n265), .Y(n338) );
  INVXL U15 ( .A(n257), .Y(n289) );
  NOR2XL U16 ( .A(n224), .B(n326), .Y(n257) );
  INVXL U17 ( .A(n150), .Y(n310) );
  AOI22XL U18 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NAND2XL U19 ( .A(n109), .B(n78), .Y(n158) );
  AOI32XL U20 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(n193) );
  NOR2XL U21 ( .A(n248), .B(n142), .Y(n357) );
  NAND2XL U22 ( .A(n140), .B(n20), .Y(n151) );
  NOR2XL U23 ( .A(n181), .B(n95), .Y(n174) );
  NAND2XL U24 ( .A(n194), .B(n274), .Y(n344) );
  NOR2XL U25 ( .A(n324), .B(n131), .Y(n262) );
  NOR2X1 U26 ( .A(a[1]), .B(n293), .Y(n318) );
  NOR2X1 U27 ( .A(n293), .B(n323), .Y(n150) );
  NAND2XL U28 ( .A(a[1]), .B(n293), .Y(n82) );
  NAND2XL U29 ( .A(n329), .B(n323), .Y(n245) );
  NAND2XL U30 ( .A(n327), .B(n266), .Y(n95) );
  NOR2XL U31 ( .A(n323), .B(n266), .Y(n187) );
  NOR2XL U32 ( .A(a[1]), .B(n242), .Y(n186) );
  NOR2X1 U33 ( .A(a[1]), .B(n103), .Y(n331) );
  INVXL U34 ( .A(n267), .Y(n333) );
  INVXL U35 ( .A(n352), .Y(n141) );
  NOR2X4 U36 ( .A(n264), .B(n197), .Y(n350) );
  NAND2X1 U37 ( .A(a[1]), .B(n31), .Y(n352) );
  INVX1 U38 ( .A(n89), .Y(n340) );
  AOI211XL U39 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  OR4X2 U40 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U41 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI31XL U42 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI211XL U43 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  AOI31XL U44 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI31XL U45 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U46 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31XL U47 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI211XL U48 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  OAI211XL U49 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U50 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U51 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI31XL U52 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U53 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI211XL U54 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI22XL U55 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI31XL U56 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  OAI22XL U57 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI211XL U58 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U59 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI21X1 U60 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  OAI211XL U61 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  OAI211XL U62 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI22XL U63 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  AOI31XL U64 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI211XL U65 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI31XL U66 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI22XL U67 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  OAI211XL U68 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U69 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  AOI211XL U70 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U71 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI31XL U72 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  NAND2XL U73 ( .A(n296), .B(n101), .Y(n94) );
  AOI31XL U74 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  INVXL U75 ( .A(n101), .Y(n254) );
  AOI31XL U76 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  AOI211XL U77 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  OAI211XL U78 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  AOI22XL U79 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U80 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  AOI22XL U81 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  NOR2XL U82 ( .A(n150), .B(n331), .Y(n130) );
  AOI22XL U83 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI211XL U84 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  OAI211XL U85 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  AOI22XL U86 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  AOI31XL U87 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI221XL U88 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI31XL U89 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  AOI31XL U90 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI211XL U91 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI211XL U92 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  NAND2XL U93 ( .A(n235), .B(n274), .Y(n184) );
  NOR2XL U94 ( .A(n224), .B(n150), .Y(n116) );
  AOI2BB2XL U95 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI211XL U96 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI22XL U97 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI22XL U98 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI22XL U99 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI22XL U100 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI22XL U101 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI211XL U102 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI211XL U103 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI22XL U104 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI2BB2XL U105 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U106 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI211XL U107 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI2BB2XL U108 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI211XL U109 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI22XL U110 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI31XL U111 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  NAND2XL U112 ( .A(n265), .B(n348), .Y(n247) );
  INVXL U113 ( .A(n152), .Y(n222) );
  AOI211XL U114 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  OAI22XL U115 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI22XL U116 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI22XL U117 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  NAND2XL U118 ( .A(n352), .B(n351), .Y(n358) );
  AOI22XL U119 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  AOI22XL U120 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  AOI22XL U121 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  OAI22XL U122 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  NAND3XL U123 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  AOI22XL U124 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  AOI22XL U125 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI211XL U126 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI22XL U127 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  AOI22XL U128 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI2BB2XL U129 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  OAI22XL U130 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI22XL U131 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  INVXL U132 ( .A(n180), .Y(n183) );
  AOI211XL U133 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  NAND2XL U134 ( .A(n103), .B(n253), .Y(n305) );
  AOI22XL U135 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  NOR2XL U136 ( .A(n293), .B(n292), .Y(n294) );
  AOI22XL U137 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  OAI2BB1XL U138 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  OAI211XL U139 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U140 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI2BB2XL U141 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  NOR2XL U142 ( .A(n209), .B(n233), .Y(n256) );
  AOI22XL U143 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  NOR2XL U144 ( .A(n161), .B(n309), .Y(n162) );
  INVXL U145 ( .A(n312), .Y(n313) );
  AOI22XL U146 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  INVXL U147 ( .A(n82), .Y(n172) );
  NAND2XL U148 ( .A(n109), .B(n242), .Y(n135) );
  AOI22XL U149 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  AOI22XL U150 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  AOI22XL U151 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  NOR2XL U152 ( .A(n268), .B(n354), .Y(n13) );
  NOR2XL U153 ( .A(n37), .B(n145), .Y(n99) );
  AOI22XL U154 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  AOI31XL U155 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI211XL U156 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  NAND2XL U157 ( .A(n311), .B(n196), .Y(n40) );
  NOR2XL U158 ( .A(n293), .B(n226), .Y(n39) );
  AOI22XL U159 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  INVXL U160 ( .A(n131), .Y(n351) );
  AOI22XL U161 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  NAND2XL U162 ( .A(n311), .B(n236), .Y(n346) );
  AOI22XL U163 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  AND2X2 U164 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U165 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AOI22XL U166 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  OAI22XL U167 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  NAND2XL U168 ( .A(n350), .B(n245), .Y(n180) );
  AOI2BB2XL U169 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U170 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI22XL U171 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  AOI22XL U172 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  AOI22XL U173 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  OAI22XL U174 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI22XL U175 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  NOR2XL U176 ( .A(n181), .B(n269), .Y(n315) );
  NOR3XL U177 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI22XL U178 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  NOR3XL U179 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  AOI22XL U180 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  AOI22XL U181 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  AOI22XL U182 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  AOI22XL U183 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NAND2XL U184 ( .A(n107), .B(n348), .Y(n175) );
  NOR2XL U185 ( .A(n37), .B(a[1]), .Y(n195) );
  NAND2XL U186 ( .A(n311), .B(n303), .Y(n38) );
  NOR2XL U187 ( .A(a[1]), .B(n329), .Y(n269) );
  NOR2XL U188 ( .A(a[1]), .B(n249), .Y(n131) );
  AOI22XL U189 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  NAND3XL U190 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NAND2XL U191 ( .A(n306), .B(n267), .Y(n61) );
  NAND3XL U192 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  NOR2XL U193 ( .A(n233), .B(n331), .Y(n108) );
  NOR2XL U194 ( .A(n187), .B(n186), .Y(n290) );
  AOI22XL U195 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NAND3XL U196 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  NAND2XL U197 ( .A(a[1]), .B(n261), .Y(n303) );
  INVXL U198 ( .A(n332), .Y(n234) );
  INVXL U199 ( .A(n297), .Y(n284) );
  NAND2XL U200 ( .A(n328), .B(n311), .Y(n353) );
  INVXL U201 ( .A(n197), .Y(n185) );
  NOR2XL U202 ( .A(a[1]), .B(n198), .Y(n160) );
  AOI22XL U203 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U204 ( .A(n264), .B(n273), .Y(n330) );
  AOI22XL U205 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  NAND2XL U206 ( .A(n264), .B(n275), .Y(n252) );
  INVXL U207 ( .A(n274), .Y(n251) );
  NAND2XL U208 ( .A(a[3]), .B(a[1]), .Y(n20) );
  INVX2 U209 ( .A(a[7]), .Y(n264) );
  NOR2XL U210 ( .A(a[3]), .B(a[1]), .Y(n225) );
  NAND2XL U211 ( .A(a[4]), .B(a[1]), .Y(n274) );
  OAI21X1 U212 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  OAI21X1 U213 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U214 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U215 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U216 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U217 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U218 ( .A(a[5]), .Y(n275) );
  NOR2X2 U219 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U220 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U221 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U222 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U223 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U224 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U225 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U226 ( .A(n233), .Y(n359) );
  NAND2X2 U227 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U228 ( .A(n349), .Y(n288) );
  NOR2X4 U229 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U230 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U231 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U232 ( .A(n347), .Y(n1) );
  CLKINVX3 U233 ( .A(a[2]), .Y(n273) );
  NOR2X4 U234 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U235 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  NAND2X2 U236 ( .A(a[6]), .B(a[0]), .Y(n360) );
  CLKINVX3 U237 ( .A(n309), .Y(n345) );
  NAND2X2 U238 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U239 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U240 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U241 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U242 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U243 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U244 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U245 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U246 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U247 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U248 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U249 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U250 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U251 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U252 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U253 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U254 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U255 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U256 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U257 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U258 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  AOI21XL U259 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U260 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  NOR2X1 U261 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U262 ( .A(a[1]), .Y(n323) );
  NAND2X1 U263 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U264 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U265 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U266 ( .A(a[4]), .B(n31), .Y(n266) );
  NOR2X1 U267 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U268 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U269 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U270 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U271 ( .A(n242), .Y(n249) );
  OAI21XL U272 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U273 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U274 ( .A(n66), .Y(n111) );
  NOR2X1 U275 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U276 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U277 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  INVX1 U278 ( .A(a[6]), .Y(n16) );
  NOR2X1 U279 ( .A(a[0]), .B(n16), .Y(n125) );
  INVX1 U280 ( .A(n261), .Y(n307) );
  INVX1 U281 ( .A(n20), .Y(n326) );
  NAND2X1 U282 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U283 ( .A(n187), .Y(n196) );
  INVX1 U284 ( .A(n350), .Y(n335) );
  NAND2X1 U285 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U286 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U287 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U288 ( .A(a[3]), .B(n323), .Y(n267) );
  INVX1 U289 ( .A(n103), .Y(n37) );
  NOR2X1 U290 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U291 ( .A(n311), .Y(n268) );
  INVX1 U292 ( .A(n293), .Y(n209) );
  NOR2X1 U293 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U294 ( .A(n224), .Y(n235) );
  NAND2X1 U295 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U296 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U297 ( .A(n195), .Y(n142) );
  NAND2X1 U298 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U299 ( .A(n226), .Y(n253) );
  NAND2X1 U300 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U301 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U302 ( .A(n1), .Y(n301) );
  NAND2X1 U303 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U304 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U305 ( .A(a[6]), .B(a[0]), .Y(n89) );
  AOI211X1 U306 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U307 ( .A(n327), .Y(n248) );
  INVX1 U308 ( .A(n181), .Y(n109) );
  INVX1 U309 ( .A(n225), .Y(n302) );
  NAND2X1 U310 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U311 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U312 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U313 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U314 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U315 ( .A(n270), .Y(n107) );
  INVX1 U316 ( .A(n306), .Y(n145) );
  NAND4X1 U317 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U318 ( .A(n210), .Y(n236) );
  INVX1 U319 ( .A(n331), .Y(n78) );
  INVX1 U320 ( .A(n328), .Y(n314) );
  OAI21XL U321 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U322 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U323 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U324 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule

//lmdpl
//module aes_sbox_8 ( a, d, preclkbar );
module aes_sbox_8 ( a, d,clk, rst,  preclkbar,m_in0_U179, m_in1_U179, m_out_U179, precharge_lmdpl);
  input [7:0] a;
  //lmdpl
  input preclkbar,clk, rst, m_in0_U179, m_in1_U179, m_out_U179, precharge_lmdpl;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  AOI211XL U4 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  AOI21XL U5 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  INVX1 U6 ( .A(n116), .Y(n203) );
  NAND2X1 U7 ( .A(n194), .B(n274), .Y(n344) );
  //wddl
  INVX1 U8 ( .A(n324), .Y(n265) );
 // WDDLINV U8 ( .A(n324), .Y(n265), .clkinv(preclkbar) );
  AOI21XL U9 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  AOI2BB2XL U10 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  INVXL U11 ( .A(n257), .Y(n289) );
  NAND2XL U12 ( .A(n235), .B(n265), .Y(n338) );
  NOR2XL U13 ( .A(n224), .B(n326), .Y(n257) );
  INVXL U14 ( .A(n150), .Y(n310) );
  AOI22XL U15 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NOR2XL U16 ( .A(n248), .B(n142), .Y(n357) );
  NAND2XL U17 ( .A(n109), .B(n78), .Y(n158) );
  //wddl
  NOR2XL U18 ( .A(n324), .B(n131), .Y(n262) );
 // WDDLNOR2X U18 ( .A(n324), .B(n131), .Y(n262), .clkinv(preclkbar) );
  NOR2XL U19 ( .A(n181), .B(n95), .Y(n174) );
  //wddl
  NAND2XL U20 ( .A(a[1]), .B(n293), .Y(n82) );
 // WDDLNAND2X U20 ( .A(a[1]), .B(n293), .Y(n82), .clkinv(preclkbar) );
  //wddl
  NOR2X1 U21 ( .A(n293), .B(n323), .Y(n150) );
  //WDDLNOR2X U21 ( .A(n293), .B(n323), .Y(n150), .clkinv(preclkbar) );
  //wddl
  NOR2X1 U22 ( .A(a[1]), .B(n293), .Y(n318) );
  //WDDLNOR2X U22 ( .A(a[1]), .B(n293), .Y(n318), .clkinv(preclkbar) );
  //wddl
  NAND2XL U23 ( .A(n140), .B(n20), .Y(n151) );
  //WDDLNAND2X U23 ( .A(n140), .B(n20), .Y(n151), .clkinv(preclkbar) );
  INVXL U24 ( .A(n352), .Y(n141) );
  INVXL U25 ( .A(n267), .Y(n333) );
  //wddl
  NOR2X1 U26 ( .A(a[1]), .B(n103), .Y(n331) );
  //WDDLNOR2X U26 ( .A(a[1]), .B(n103), .Y(n331), .clkinv(preclkbar) );
  //wddl
  NOR2XL U27 ( .A(a[1]), .B(n242), .Y(n186) );
  //WDDLNOR2X U27 ( .A(a[1]), .B(n242), .Y(n186), .clkinv(preclkbar) );
  NOR2X4 U28 ( .A(n264), .B(n197), .Y(n350) );
  //wddl
  NAND2X1 U29 ( .A(a[1]), .B(n31), .Y(n352) );
  //WDDLNAND2X U29 ( .A(a[1]), .B(n31), .Y(n352), .clkinv(preclkbar) );
  AOI211XL U30 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  OR4X2 U31 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U32 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI31XL U33 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI211XL U34 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U35 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U36 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI31XL U37 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI31XL U38 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U39 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  OAI211XL U40 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U41 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U42 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI211XL U43 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI31XL U44 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  OAI22XL U45 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  OAI211XL U46 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI211XL U47 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI22XL U48 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  AOI31XL U49 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U50 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U51 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI22XL U52 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  OAI211XL U53 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI211XL U54 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI211XL U55 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI31XL U56 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI31XL U57 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI22XL U58 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  NAND2XL U59 ( .A(n296), .B(n101), .Y(n94) );
  AOI211XL U60 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  OAI211XL U61 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  OAI211XL U62 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  INVXL U63 ( .A(n101), .Y(n254) );
  AOI211XL U64 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  AOI31XL U65 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  AOI31XL U66 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  AOI211XL U67 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U68 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI22XL U69 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U70 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  OAI211XL U71 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  AOI22XL U72 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  AOI31XL U73 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI22XL U74 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI211XL U75 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  NOR2XL U76 ( .A(n150), .B(n331), .Y(n130) );
  AOI22XL U77 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  AOI211XL U78 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  AOI31XL U79 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  NAND2XL U80 ( .A(n235), .B(n274), .Y(n184) );
  NOR2XL U81 ( .A(n224), .B(n150), .Y(n116) );
  AOI211XL U82 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI221XL U83 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI31XL U84 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI22XL U85 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI211XL U86 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI211XL U87 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI2BB2XL U88 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI211XL U89 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI22XL U90 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI31XL U91 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI2BB2XL U92 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U93 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI22XL U94 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI22XL U95 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI22XL U96 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  OAI22XL U97 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI22XL U98 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI211XL U99 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI211XL U100 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  INVXL U101 ( .A(n152), .Y(n222) );
  AOI2BB2XL U102 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  NAND2XL U103 ( .A(n265), .B(n348), .Y(n247) );
  AOI211XL U104 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI22XL U105 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI22XL U106 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI22XL U107 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  NOR2XL U108 ( .A(n293), .B(n292), .Y(n294) );
  NAND2XL U109 ( .A(n103), .B(n253), .Y(n305) );
  INVXL U110 ( .A(n312), .Y(n313) );
  AOI22XL U111 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  INVXL U112 ( .A(n180), .Y(n183) );
  AOI211XL U113 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  AOI22XL U114 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  AOI22XL U115 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  OAI2BB1XL U116 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  NOR2XL U117 ( .A(n209), .B(n233), .Y(n256) );
  AOI2BB2XL U118 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  AOI22XL U119 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  OAI211XL U120 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  //wddl
  NAND2XL U121 ( .A(n352), .B(n351), .Y(n358) );
  //WDDLNAND2X U121 ( .A(n352), .B(n351), .Y(n358), .clkinv(preclkbar) );
  AOI32XL U122 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  AOI22XL U123 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  AOI22XL U124 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  OAI22XL U125 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  OAI22XL U126 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  NAND3XL U127 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  AOI22XL U128 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  AOI2BB2XL U129 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U130 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI22XL U131 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI22XL U132 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  AOI211XL U133 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI22XL U134 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  AOI22XL U135 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  NOR2XL U136 ( .A(n161), .B(n309), .Y(n162) );
  NAND2XL U137 ( .A(n109), .B(n242), .Y(n135) );
  INVXL U138 ( .A(n82), .Y(n172) );
  AOI22XL U139 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  NOR3XL U140 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  OAI22XL U141 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U142 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AOI22XL U143 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AND2X2 U144 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U145 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  NAND2XL U146 ( .A(n311), .B(n236), .Y(n346) );
  NOR2XL U147 ( .A(n181), .B(n269), .Y(n315) );
  //wddl
  INVXL U148 ( .A(n131), .Y(n351) );
  //WDDLINV U148 ( .A(n131), .Y(n351), .clkinv(preclkbar) );
  NOR3XL U149 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI22XL U150 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  AOI22XL U151 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  NOR2XL U152 ( .A(n293), .B(n226), .Y(n39) );
  NAND2XL U153 ( .A(n311), .B(n196), .Y(n40) );
  AOI211XL U154 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  AOI31XL U155 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI22XL U156 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  AOI22XL U157 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  NOR2XL U158 ( .A(n268), .B(n354), .Y(n13) );
  AOI22XL U159 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  AOI22XL U160 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  AOI22XL U161 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI2BB2XL U162 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  NAND2XL U163 ( .A(n350), .B(n245), .Y(n180) );
  AOI22XL U164 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  //wddl
  NOR2XL U165 ( .A(n37), .B(n145), .Y(n99) );
  //WDDLNOR2X U165 ( .A(n37), .B(n145), .Y(n99), .clkinv(preclkbar) );
  AOI22XL U166 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  OAI22XL U167 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI22XL U168 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  AOI22XL U169 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  AOI22XL U170 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  AOI22XL U171 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NOR2XL U172 ( .A(n187), .B(n186), .Y(n290) );
  NAND3XL U173 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  //wddl
 // NOR2XL U174 ( .A(a[1]), .B(n329), .Y(n269) );
  nor_lmdpl U174 ( .clk(clk), .rst_n(rst), .precharge(precharge_lmdpl), .in0(a[1]), .in1(n329), .m_in0(m_in0_U179), .m_in1(m_in1_U179), .m_out(m_out_U179), .out(n269));
  //WDDLNOR2X U174 ( .A(a[1]), .B(n329), .Y(n269), .clkinv(preclkbar) );
  AOI22XL U175 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  NAND2XL U176 ( .A(n311), .B(n303), .Y(n38) );
  //wddl
  NAND2XL U177 ( .A(n306), .B(n267), .Y(n61) );
  //WDDLNAND2X U177 ( .A(n306), .B(n267), .Y(n61), .clkinv(preclkbar) );
  //wddl
  //NOR2XL U178 ( .A(a[1]), .B(n249), .Y(n131) );
  nor_lmdpl U178 ( .clk(clk), .rst_n(rst), .precharge(precharge_lmdpl), .in0(a[1]), .in1(n249), .m_in0(m_in0_U179), .m_in1(m_in1_U179), .m_out(m_out_U179), .out(n131));
  //WDDLNOR2X U178 ( .A(a[1]), .B(n249), .Y(n131), .clkinv(preclkbar) );
  //wddl
  //NOR2XL U179 ( .A(n37), .B(a[1]), .Y(n195) );
  nor_lmdpl U179 ( .clk(clk), .rst_n(rst), .precharge(precharge_lmdpl), .in0(n37), .in1(a[1]), .m_in0(m_in0_U179), .m_in1(m_in1_U179), .m_out(m_out_U179), .out(n195));
  //WDDLNOR2X U179 ( .A(n37), .B(a[1]), .Y(n195), .clkinv(preclkbar) );
  //wddl
  NAND2XL U180 ( .A(n107), .B(n348), .Y(n175) );
  //WDDLNAND2X U180 ( .A(n107), .B(n348), .Y(n175), .clkinv(preclkbar) );
  NOR2XL U181 ( .A(n233), .B(n331), .Y(n108) );
  //nor_lmdpl U181 ( .clk(clk), .rst_n(rst), .precharge(precharge_lmdpl), .in0(n233), .in1(n331), .m_in0(m_in0_U179), .m_in1(m_in1_U179), .m_out(m_out_U179), .out(n108));
  NAND3XL U182 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  AOI22XL U183 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  AOI22XL U184 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  AOI22XL U185 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NAND2XL U186 ( .A(n329), .B(n323), .Y(n245) );
  NAND3XL U187 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  //wddl
  NAND2XL U188 ( .A(a[1]), .B(n261), .Y(n303) );
  //WDDLNAND2X U188 ( .A(a[1]), .B(n261), .Y(n303), .clkinv(preclkbar) );
  INVXL U189 ( .A(n332), .Y(n234) );
  INVXL U190 ( .A(n297), .Y(n284) );
  NAND2XL U191 ( .A(n328), .B(n311), .Y(n353) );
  INVXL U192 ( .A(n197), .Y(n185) );
  NOR2XL U193 ( .A(n264), .B(n273), .Y(n330) );
  //wddl
  NOR2XL U194 ( .A(a[1]), .B(n198), .Y(n160) );
  //WDDLNOR2X U194 ( .A(a[1]), .B(n198), .Y(n160), .clkinv(preclkbar) );
  INVXL U195 ( .A(n274), .Y(n251) );
  NAND2XL U196 ( .A(n264), .B(n275), .Y(n252) );
  AOI22XL U197 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  AOI22XL U198 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  //wddl
  NOR2XL U199 ( .A(a[3]), .B(a[1]), .Y(n225) );
  //WDDLNOR2X U199 ( .A(a[3]), .B(a[1]), .Y(n225), .clkinv(preclkbar) );
  //wddl
  NAND2XL U200 ( .A(a[3]), .B(a[1]), .Y(n20) );
  //WDDLNAND2X U200 ( .A(a[3]), .B(a[1]), .Y(n20), .clkinv(preclkbar) );
  //wddl
  NAND2XL U201 ( .A(a[4]), .B(a[1]), .Y(n274) );
  //WDDLNAND2X U201 ( .A(a[4]), .B(a[1]), .Y(n274), .clkinv(preclkbar) );
  INVX2 U202 ( .A(a[7]), .Y(n264) );
  CLKINVX3 U203 ( .A(n266), .Y(n329) );
  NAND2X2 U204 ( .A(a[4]), .B(n31), .Y(n266) );
  NAND2X2 U205 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U206 ( .A(a[5]), .Y(n275) );
  OAI21X1 U207 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U208 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U209 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NOR2X2 U210 ( .A(n31), .B(n198), .Y(n261) );
  //wddl
  NOR2X2 U211 ( .A(n37), .B(n323), .Y(n181) );
  //WDDLNOR2X U211 ( .A(n37), .B(n323), .Y(n181),.clkinv(preclkbar) );
  NOR2X2 U212 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U213 ( .A(n249), .B(n329), .Y(n293) );
  //wddl
  NOR2X2 U214 ( .A(n329), .B(n323), .Y(n226) );
  //WDDLNOR2X U214 ( .A(n329), .B(n323), .Y(n226), .clkinv(preclkbar) );
  //wddl
  NAND2X2 U215 ( .A(n198), .B(n323), .Y(n311) );
  //WDDLNAND2X U215 ( .A(n198), .B(n323), .Y(n311), .clkinv(preclkbar) );
  CLKINVX3 U216 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U217 ( .A(n233), .Y(n359) );
  NAND2X2 U218 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U219 ( .A(n349), .Y(n288) );
  NOR2X4 U220 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U221 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U222 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U223 ( .A(n347), .Y(n1) );
  CLKINVX3 U224 ( .A(a[2]), .Y(n273) );
  OAI21X1 U225 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U226 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U227 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U228 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U229 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U230 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  AOI31X4 U231 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  CLKINVX3 U232 ( .A(n309), .Y(n345) );
  NAND2X2 U233 ( .A(n275), .B(n325), .Y(n309) );
  //wddl
  NAND2X2 U234 ( .A(a[1]), .B(n242), .Y(n306) );
  //WDDLNAND2X U234 ( .A(a[1]), .B(n242), .Y(n306), .clkinv(preclkbar) );
  NAND2X2 U235 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U236 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U237 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U238 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U239 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U240 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U241 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U242 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U243 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U244 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U245 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U246 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U247 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U248 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U249 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U250 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U251 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U252 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U253 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U254 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U255 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U256 ( .A(n273), .B(n129), .Y(n347) );
  //wddl
  //CLKINVX3 U257 ( .A(a[1]), .Y(n323) );
  WDDLINV U257 ( .A(a[1]), .Y(n323), .clkinv(preclkbar) );
  NAND2X1 U258 ( .A(a[7]), .B(a[5]), .Y(n129) );
  //wddl
  NOR2X1 U259 ( .A(n323), .B(n242), .Y(n210) );
  //WDDLNOR2X U259 ( .A(n323), .B(n242), .Y(n210), .clkinv(preclkbar) );
  NAND2X1 U260 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U261 ( .A(n327), .B(n266), .Y(n95) );
  //wddl
  NOR2X1 U262 ( .A(a[4]), .B(n323), .Y(n270) );
  //WDDLNOR2X U262 ( .A(a[4]), .B(n323), .Y(n270), .clkinv(preclkbar) );
  OAI21XL U263 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U264 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U265 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U266 ( .A(n242), .Y(n249) );
  OAI21XL U267 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U268 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U269 ( .A(n192), .Y(n205) );
  INVX1 U270 ( .A(n66), .Y(n111) );
  //wddl
  NOR2X1 U271 ( .A(n261), .B(n323), .Y(n324) );
  //WDDLNOR2X U271 ( .A(n261), .B(n323), .Y(n324), .clkinv(preclkbar) );
  NAND3X1 U272 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U273 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U274 ( .A(a[6]), .B(a[0]), .Y(n360) );
  INVX1 U275 ( .A(a[6]), .Y(n16) );
  NOR2X1 U276 ( .A(a[0]), .B(n16), .Y(n125) );
  //wddl
  NOR2X1 U277 ( .A(n323), .B(n266), .Y(n187) );
  //WDDLNOR2X U277 ( .A(n323), .B(n266), .Y(n187), .clkinv(preclkbar) );
  INVX1 U278 ( .A(n261), .Y(n307) );
  INVX1 U279 ( .A(n20), .Y(n326) );
  //wddl
  NAND2X1 U280 ( .A(n261), .B(n323), .Y(n348) );
  //WDDLNAND2X U280 ( .A(n261), .B(n323), .Y(n348), .clkinv(preclkbar) );
  INVX1 U281 ( .A(n187), .Y(n196) );
  INVX1 U282 ( .A(n350), .Y(n335) );
  NAND2X1 U283 ( .A(n31), .B(n198), .Y(n103) );
  //wddl
  NAND2X1 U284 ( .A(n20), .B(n245), .Y(n263) );
  //WDDLNAND2X U284 ( .A(n20), .B(n245), .Y(n263), .clkinv(preclkbar) );
  NAND4X1 U285 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  //wddl
  NAND2X1 U286 ( .A(a[3]), .B(n323), .Y(n267) );
  //WDDLNAND2X U286 ( .A(a[3]), .B(n323), .Y(n267), .clkinv(preclkbar) );
  AOI22X1 U287 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U288 ( .A(n103), .Y(n37) );
  NOR2X1 U289 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U290 ( .A(n311), .Y(n268) );
  INVX1 U291 ( .A(n293), .Y(n209) );
  //wddl
  NOR2X1 U292 ( .A(a[1]), .B(n209), .Y(n224) );
  //WDDLNOR2X U292 ( .A(a[1]), .B(n209), .Y(n224), .clkinv(preclkbar) );
  INVX1 U293 ( .A(n224), .Y(n235) );
  //wddl
  NAND2X1 U294 ( .A(n323), .B(n307), .Y(n140) );
  //WDDLNAND2X U294 ( .A(n323), .B(n307), .Y(n140), .clkinv(preclkbar) );
  NOR2BX1 U295 ( .AN(n140), .B(n181), .Y(n92) );
 //wddl
  //INVX1 U296 ( .A(n195), .Y(n142) ); 
  WDDLINV U296 ( .A(n195), .Y(n142), .clkinv(preclkbar) );
  NAND2X1 U297 ( .A(a[0]), .B(n16), .Y(n297) );
  //wddl
  INVX1 U298 ( .A(n226), .Y(n253) );
  //WDDLINV U298 ( .A(n226), .Y(n253), .clkinv(preclkbar) );
  NAND2X1 U299 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U300 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U301 ( .A(n1), .Y(n301) );
  NAND2X1 U302 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U303 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U304 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U305 ( .A(n89), .Y(n340) );
  AOI211X1 U306 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U307 ( .A(n327), .Y(n248) );
  //wddl
  INVX1 U308 ( .A(n181), .Y(n109) );
  //WDDLINV U308 ( .A(n181), .Y(n109), .clkinv(preclkbar) );
  INVX1 U309 ( .A(n225), .Y(n302) );
  //wddl
  NAND2X1 U310 ( .A(n109), .B(n302), .Y(n100) );
  //WDDLNAND2X U310 ( .A(n109), .B(n302), .Y(n100), .clkinv(preclkbar) );
  OAI21XL U311 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U312 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U313 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U314 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U315 ( .A(n270), .Y(n107) );
  //wddl
  INVX1 U316 ( .A(n306), .Y(n145) );
  //WDDLINV U316 ( .A(n306), .Y(n145), .clkinv(preclkbar) );
  NAND4X1 U317 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U318 ( .A(n210), .Y(n236) );
  INVX1 U319 ( .A(n331), .Y(n78) );
  INVX1 U320 ( .A(n328), .Y(n314) );
  OAI21XL U321 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U322 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U323 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U324 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  //wddl
  INVX1 U332 ( .A(n72), .Y(n204) );
  //WDDLINV U332 ( .A(n72), .Y(n204), .clkinv(preclkbar) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  //wddl
  //NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  nor_lmdpl U338 ( .clk(clk), .rst_n(rst), .precharge(precharge_lmdpl), .in0(n145), .in1(n318), .m_in0(m_in0_U179), .m_in1(m_in1_U179), .m_out(m_out_U179), .out(n152));
  //WDDLNOR2X U338 ( .A(n145), .B(n318), .Y(n152), .clkinv(preclkbar) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  //wddl
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  //WDDLNOR2X U342 ( .A(n103), .B(n323), .Y(n355), .clkinv(preclkbar) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_9 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U2 ( .AN(n348), .B(n309), .Y(n246) );
  AOI21XL U3 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  AOI211XL U4 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  INVX1 U5 ( .A(n116), .Y(n203) );
  NAND2X1 U6 ( .A(n194), .B(n274), .Y(n344) );
  INVX1 U7 ( .A(n296), .Y(n354) );
  INVX1 U8 ( .A(n324), .Y(n265) );
  AOI21XL U9 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  AOI2BB2XL U10 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  NAND2XL U11 ( .A(n235), .B(n265), .Y(n338) );
  INVXL U12 ( .A(n257), .Y(n289) );
  NOR2XL U13 ( .A(n224), .B(n326), .Y(n257) );
  AOI22XL U14 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NAND2XL U15 ( .A(n109), .B(n78), .Y(n158) );
  NOR2XL U16 ( .A(n248), .B(n142), .Y(n357) );
  NOR2X1 U17 ( .A(n293), .B(n323), .Y(n150) );
  NAND2XL U18 ( .A(a[1]), .B(n293), .Y(n82) );
  NOR2X1 U19 ( .A(a[1]), .B(n293), .Y(n318) );
  NOR2XL U20 ( .A(n324), .B(n131), .Y(n262) );
  NOR2XL U21 ( .A(n181), .B(n95), .Y(n174) );
  NAND2XL U22 ( .A(n140), .B(n20), .Y(n151) );
  INVXL U23 ( .A(n352), .Y(n141) );
  INVXL U24 ( .A(n267), .Y(n333) );
  NOR2X1 U25 ( .A(a[1]), .B(n103), .Y(n331) );
  NOR2XL U26 ( .A(a[1]), .B(n242), .Y(n186) );
  NOR2X4 U27 ( .A(n264), .B(n197), .Y(n350) );
  NAND2X1 U28 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI31XL U29 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI211XL U30 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  OR4X2 U31 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U32 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U33 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI31XL U34 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U35 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI31XL U36 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI211XL U37 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U38 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI31XL U39 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  OAI211XL U40 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U41 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI22XL U42 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  AOI22XL U43 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  OAI211XL U44 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI211XL U45 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  OAI22XL U46 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI31XL U47 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  OAI211XL U48 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI31XL U49 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI211XL U50 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI211XL U51 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI22XL U52 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI211XL U53 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI31XL U54 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U55 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI211XL U56 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI31XL U57 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  OAI211XL U58 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U59 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  AOI31XL U60 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  INVXL U61 ( .A(n101), .Y(n254) );
  AOI211XL U62 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U63 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI22XL U64 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U65 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  NAND2XL U66 ( .A(n296), .B(n101), .Y(n94) );
  OAI211XL U67 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  AOI31XL U68 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  AOI211XL U69 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  NOR2XL U70 ( .A(n224), .B(n150), .Y(n116) );
  NOR2XL U71 ( .A(n150), .B(n331), .Y(n130) );
  INVXL U72 ( .A(n150), .Y(n310) );
  AOI211XL U73 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  AOI22XL U74 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  NAND2XL U75 ( .A(n235), .B(n274), .Y(n184) );
  AOI31XL U76 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI22XL U77 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI211XL U78 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI31XL U79 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI221XL U80 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI22XL U81 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  OAI211XL U82 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  AOI211XL U83 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI31XL U84 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  OAI22XL U85 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI22XL U86 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI22XL U87 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI22XL U88 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI22XL U89 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI2BB2XL U90 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U91 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI22XL U92 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI211XL U93 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI211XL U94 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI22XL U95 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI211XL U96 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI22XL U97 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI22XL U98 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI2BB2XL U99 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  NAND2XL U100 ( .A(n265), .B(n348), .Y(n247) );
  INVXL U101 ( .A(n152), .Y(n222) );
  AOI2BB2XL U102 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI211XL U103 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI31XL U104 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI22XL U105 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI211XL U106 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI211XL U107 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  OAI2BB1XL U108 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  AOI22XL U109 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  AOI22XL U110 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  OAI211XL U111 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U112 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI2BB2XL U113 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  NOR2XL U114 ( .A(n209), .B(n233), .Y(n256) );
  AOI211XL U115 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI22XL U116 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI22XL U117 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  AOI22XL U118 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  NAND3XL U119 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  OAI22XL U120 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  NAND2XL U121 ( .A(n109), .B(n242), .Y(n135) );
  AOI22XL U122 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  AOI22XL U123 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  AOI22XL U124 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  AOI211XL U125 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  INVXL U126 ( .A(n180), .Y(n183) );
  OAI22XL U127 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI2BB2XL U128 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI32XL U129 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  AOI22XL U130 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  INVXL U131 ( .A(n82), .Y(n172) );
  AOI22XL U132 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  NOR2XL U133 ( .A(n161), .B(n309), .Y(n162) );
  NOR2XL U134 ( .A(n293), .B(n292), .Y(n294) );
  NAND2XL U135 ( .A(n103), .B(n253), .Y(n305) );
  AOI22XL U136 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  INVXL U137 ( .A(n312), .Y(n313) );
  NAND2XL U138 ( .A(n352), .B(n351), .Y(n358) );
  AOI31XL U139 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI22XL U140 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  NOR3XL U141 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI211XL U142 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  AOI22XL U143 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  NAND2XL U144 ( .A(n311), .B(n196), .Y(n40) );
  NOR2XL U145 ( .A(n293), .B(n226), .Y(n39) );
  AOI22XL U146 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  NAND2XL U147 ( .A(n311), .B(n236), .Y(n346) );
  AOI22XL U148 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  INVXL U149 ( .A(n131), .Y(n351) );
  OAI22XL U150 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  NOR2XL U151 ( .A(n37), .B(n145), .Y(n99) );
  AOI22XL U152 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  AOI22XL U153 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  NOR2XL U154 ( .A(n181), .B(n269), .Y(n315) );
  AOI22XL U155 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  NOR2XL U156 ( .A(n268), .B(n354), .Y(n13) );
  AOI22XL U157 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  AND2X2 U158 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U159 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  AOI22XL U160 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AOI22XL U161 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  AOI22XL U162 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  OAI22XL U163 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  NAND2XL U164 ( .A(n350), .B(n245), .Y(n180) );
  NOR3XL U165 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  AOI2BB2XL U166 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U167 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  AOI22XL U168 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  AOI22XL U169 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  NAND2XL U170 ( .A(n107), .B(n348), .Y(n175) );
  AOI22XL U171 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  AOI22XL U172 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  NOR2XL U173 ( .A(a[1]), .B(n329), .Y(n269) );
  AOI22XL U174 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NAND2XL U175 ( .A(n329), .B(n323), .Y(n245) );
  NAND2XL U176 ( .A(n306), .B(n267), .Y(n61) );
  AOI22XL U177 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  NOR2XL U178 ( .A(n187), .B(n186), .Y(n290) );
  NOR2XL U179 ( .A(n37), .B(a[1]), .Y(n195) );
  NOR2XL U180 ( .A(a[1]), .B(n249), .Y(n131) );
  NAND3XL U181 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  AOI22XL U182 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  AOI22XL U183 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  NAND2XL U184 ( .A(n311), .B(n303), .Y(n38) );
  NOR2XL U185 ( .A(n233), .B(n331), .Y(n108) );
  NAND3XL U186 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  INVXL U187 ( .A(n297), .Y(n284) );
  INVXL U188 ( .A(n197), .Y(n185) );
  NAND2XL U189 ( .A(a[1]), .B(n261), .Y(n303) );
  NAND2XL U190 ( .A(n328), .B(n311), .Y(n353) );
  NAND3XL U191 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  INVXL U192 ( .A(n332), .Y(n234) );
  AOI22XL U193 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U194 ( .A(a[1]), .B(n198), .Y(n160) );
  AOI22XL U195 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  INVXL U196 ( .A(n274), .Y(n251) );
  NAND2XL U197 ( .A(n264), .B(n275), .Y(n252) );
  NOR2XL U198 ( .A(n264), .B(n273), .Y(n330) );
  NAND2XL U199 ( .A(a[3]), .B(a[1]), .Y(n20) );
  INVX2 U200 ( .A(a[7]), .Y(n264) );
  NOR2XL U201 ( .A(a[3]), .B(a[1]), .Y(n225) );
  NAND2XL U202 ( .A(a[4]), .B(a[1]), .Y(n274) );
  CLKINVX3 U203 ( .A(n266), .Y(n329) );
  NAND2X2 U204 ( .A(a[4]), .B(n31), .Y(n266) );
  NAND2X2 U205 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U206 ( .A(a[5]), .Y(n275) );
  OAI21X1 U207 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U208 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U209 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NOR2X2 U210 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U211 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U212 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U213 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U214 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U215 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U216 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U217 ( .A(n233), .Y(n359) );
  NAND2X2 U218 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U219 ( .A(n349), .Y(n288) );
  NOR2X4 U220 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U221 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U222 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U223 ( .A(n347), .Y(n1) );
  CLKINVX3 U224 ( .A(a[2]), .Y(n273) );
  OAI21X1 U225 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U226 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U227 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U228 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U229 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U230 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  AOI31X4 U231 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  CLKINVX3 U232 ( .A(n309), .Y(n345) );
  NAND2X2 U233 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U234 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U235 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U236 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U237 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U238 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U239 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U240 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U241 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U242 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U243 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U244 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U245 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U246 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U247 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U248 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U249 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U250 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U251 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U252 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U253 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U254 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U255 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U256 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U257 ( .A(a[1]), .Y(n323) );
  NAND2X1 U258 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U259 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U260 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U261 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U262 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U263 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U264 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U265 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U266 ( .A(n242), .Y(n249) );
  OAI21XL U267 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U268 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U269 ( .A(n192), .Y(n205) );
  INVX1 U270 ( .A(n66), .Y(n111) );
  NOR2X1 U271 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U272 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U273 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U274 ( .A(a[6]), .B(a[0]), .Y(n360) );
  INVX1 U275 ( .A(a[6]), .Y(n16) );
  NOR2X1 U276 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U277 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U278 ( .A(n261), .Y(n307) );
  INVX1 U279 ( .A(n20), .Y(n326) );
  NAND2X1 U280 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U281 ( .A(n187), .Y(n196) );
  INVX1 U282 ( .A(n350), .Y(n335) );
  NAND2X1 U283 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U284 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U285 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U286 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U287 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U288 ( .A(n103), .Y(n37) );
  NOR2X1 U289 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U290 ( .A(n311), .Y(n268) );
  INVX1 U291 ( .A(n293), .Y(n209) );
  NOR2X1 U292 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U293 ( .A(n224), .Y(n235) );
  NAND2X1 U294 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U295 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U296 ( .A(n195), .Y(n142) );
  NAND2X1 U297 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U298 ( .A(n226), .Y(n253) );
  NAND2X1 U299 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U300 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U301 ( .A(n1), .Y(n301) );
  NAND2X1 U302 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U303 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U304 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U305 ( .A(n89), .Y(n340) );
  AOI211X1 U306 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U307 ( .A(n327), .Y(n248) );
  INVX1 U308 ( .A(n181), .Y(n109) );
  INVX1 U309 ( .A(n225), .Y(n302) );
  NAND2X1 U310 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U311 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U312 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U313 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U314 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U315 ( .A(n270), .Y(n107) );
  INVX1 U316 ( .A(n306), .Y(n145) );
  NAND4X1 U317 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U318 ( .A(n210), .Y(n236) );
  INVX1 U319 ( .A(n331), .Y(n78) );
  INVX1 U320 ( .A(n328), .Y(n314) );
  OAI21XL U321 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U322 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U323 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U324 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_10 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  AOI21XL U4 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  NAND2X1 U5 ( .A(n235), .B(n265), .Y(n338) );
  NAND2X1 U6 ( .A(n194), .B(n274), .Y(n344) );
  AOI211XL U7 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  AOI21XL U8 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  INVXL U9 ( .A(n116), .Y(n203) );
  INVXL U10 ( .A(n257), .Y(n289) );
  INVXL U11 ( .A(n150), .Y(n310) );
  NOR2XL U12 ( .A(n224), .B(n326), .Y(n257) );
  AOI22XL U13 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  NOR2XL U14 ( .A(n248), .B(n142), .Y(n357) );
  NAND2XL U15 ( .A(n109), .B(n78), .Y(n158) );
  NOR2XL U16 ( .A(n324), .B(n131), .Y(n262) );
  NOR2X1 U17 ( .A(a[1]), .B(n293), .Y(n318) );
  NOR2XL U18 ( .A(n181), .B(n95), .Y(n174) );
  NOR2X1 U19 ( .A(n268), .B(n354), .Y(n13) );
  NOR2X1 U20 ( .A(n293), .B(n323), .Y(n150) );
  NAND2XL U21 ( .A(a[1]), .B(n293), .Y(n82) );
  INVX2 U22 ( .A(n324), .Y(n265) );
  NOR2X1 U23 ( .A(a[1]), .B(n103), .Y(n331) );
  NOR2X4 U24 ( .A(n264), .B(n197), .Y(n350) );
  INVXL U25 ( .A(n352), .Y(n141) );
  NOR2XL U26 ( .A(a[1]), .B(n242), .Y(n186) );
  INVXL U27 ( .A(n267), .Y(n333) );
  NAND2X1 U28 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI211XL U29 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  AOI211XL U30 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  OR4X2 U31 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U32 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI31XL U33 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI31XL U34 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  OAI211XL U35 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U36 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI31XL U37 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI31XL U38 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI31XL U39 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI211XL U40 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U41 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  OAI211XL U42 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  OAI211XL U43 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI31XL U44 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI22XL U45 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  AOI31XL U46 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  AOI31XL U47 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI211XL U48 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI22XL U49 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  OAI22XL U50 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI22XL U51 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI211XL U52 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI31XL U53 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U54 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI211XL U55 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI211XL U56 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI211XL U57 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U58 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  AOI31XL U59 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  OAI211XL U60 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U61 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI2BB2XL U62 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  OAI211XL U63 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  NAND2XL U64 ( .A(n296), .B(n101), .Y(n94) );
  INVXL U65 ( .A(n101), .Y(n254) );
  AOI31XL U66 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  AOI22XL U67 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U68 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U69 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U70 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  NOR2XL U71 ( .A(n224), .B(n150), .Y(n116) );
  AOI31XL U72 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI22XL U73 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI22XL U74 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  AOI211XL U75 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI211XL U76 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  NOR2XL U77 ( .A(n150), .B(n331), .Y(n130) );
  AOI22XL U78 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  NAND2XL U79 ( .A(n235), .B(n274), .Y(n184) );
  AOI31XL U80 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI211XL U81 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  AOI221XL U82 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI31XL U83 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  OAI211XL U84 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  AOI211XL U85 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI211XL U86 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI211XL U87 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI22XL U88 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI22XL U89 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI22XL U90 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI211XL U91 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI2BB2XL U92 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI22XL U93 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI22XL U94 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI2BB2XL U95 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U96 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  OAI22XL U97 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI211XL U98 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI22XL U99 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  INVXL U100 ( .A(n152), .Y(n222) );
  AOI22XL U101 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI31XL U102 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI22XL U103 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  NAND2XL U104 ( .A(n265), .B(n348), .Y(n247) );
  AOI2BB2XL U105 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI211XL U106 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI22XL U107 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI22XL U108 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  AOI2BB2XL U109 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  INVXL U110 ( .A(n180), .Y(n183) );
  INVXL U111 ( .A(n82), .Y(n172) );
  AOI211XL U112 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  OAI2BB1XL U113 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  AOI22XL U114 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  NOR2XL U115 ( .A(n293), .B(n292), .Y(n294) );
  NAND2XL U116 ( .A(n103), .B(n253), .Y(n305) );
  AOI22XL U117 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  NAND2XL U118 ( .A(n352), .B(n351), .Y(n358) );
  OAI211XL U119 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U120 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI22XL U121 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI2BB2XL U122 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  AOI22XL U123 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  OAI22XL U124 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  INVXL U125 ( .A(n312), .Y(n313) );
  AOI22XL U126 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  NOR2XL U127 ( .A(n161), .B(n309), .Y(n162) );
  NAND2XL U128 ( .A(n109), .B(n242), .Y(n135) );
  AOI211XL U129 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI22XL U130 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  AOI32XL U131 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  AOI22XL U132 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  AOI22XL U133 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI22XL U134 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  OAI22XL U135 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  NAND3XL U136 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  NOR2XL U137 ( .A(n209), .B(n233), .Y(n256) );
  AOI2BB2XL U138 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U139 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  AOI22XL U140 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI22XL U141 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  AOI22XL U142 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  OAI22XL U143 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI22XL U144 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  AOI22XL U145 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  NOR2XL U146 ( .A(n293), .B(n226), .Y(n39) );
  NAND2XL U147 ( .A(n350), .B(n245), .Y(n180) );
  OAI22XL U148 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U149 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AOI22XL U150 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AND2X2 U151 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U152 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  NAND2XL U153 ( .A(n311), .B(n236), .Y(n346) );
  AOI22XL U154 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  NOR3XL U155 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  AOI22XL U156 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  NOR2XL U157 ( .A(n181), .B(n269), .Y(n315) );
  AOI211XL U158 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  NOR3XL U159 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  INVXL U160 ( .A(n131), .Y(n351) );
  AOI22XL U161 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  NAND2XL U162 ( .A(n311), .B(n196), .Y(n40) );
  NOR2XL U163 ( .A(n37), .B(n145), .Y(n99) );
  AOI22XL U164 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  AOI22XL U165 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  AOI31XL U166 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI22XL U167 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  AOI22XL U168 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  NOR2XL U169 ( .A(a[1]), .B(n249), .Y(n131) );
  AOI22XL U170 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NAND3XL U171 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  AOI22XL U172 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  AOI22XL U173 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  AOI22XL U174 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NOR2XL U175 ( .A(n233), .B(n331), .Y(n108) );
  NOR2XL U176 ( .A(n37), .B(a[1]), .Y(n195) );
  NOR2XL U177 ( .A(a[1]), .B(n329), .Y(n269) );
  NOR2XL U178 ( .A(n187), .B(n186), .Y(n290) );
  NAND2XL U179 ( .A(n306), .B(n267), .Y(n61) );
  NAND2XL U180 ( .A(n311), .B(n303), .Y(n38) );
  NAND3XL U181 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NAND2XL U182 ( .A(n107), .B(n348), .Y(n175) );
  AOI22XL U183 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  NAND2XL U184 ( .A(n329), .B(n323), .Y(n245) );
  NAND2XL U185 ( .A(n328), .B(n311), .Y(n353) );
  NAND2XL U186 ( .A(a[1]), .B(n261), .Y(n303) );
  NAND3XL U187 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  INVXL U188 ( .A(n197), .Y(n185) );
  INVXL U189 ( .A(n332), .Y(n234) );
  INVXL U190 ( .A(n297), .Y(n284) );
  NOR2XL U191 ( .A(a[1]), .B(n198), .Y(n160) );
  AOI22XL U192 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  AOI22XL U193 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  INVXL U194 ( .A(n274), .Y(n251) );
  NOR2XL U195 ( .A(n264), .B(n273), .Y(n330) );
  NAND2XL U196 ( .A(n264), .B(n275), .Y(n252) );
  NOR2XL U197 ( .A(a[3]), .B(a[1]), .Y(n225) );
  NAND2XL U198 ( .A(a[3]), .B(a[1]), .Y(n20) );
  INVX2 U199 ( .A(a[7]), .Y(n264) );
  INVX1 U200 ( .A(a[6]), .Y(n16) );
  NAND2XL U201 ( .A(a[4]), .B(a[1]), .Y(n274) );
  CLKINVX3 U202 ( .A(n266), .Y(n329) );
  NAND2X2 U203 ( .A(a[4]), .B(n31), .Y(n266) );
  NAND2X2 U204 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U205 ( .A(a[5]), .Y(n275) );
  OAI21X1 U206 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U207 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U208 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NOR2X2 U209 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U210 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U211 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U212 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U213 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U214 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U215 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U216 ( .A(n233), .Y(n359) );
  NAND2X2 U217 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U218 ( .A(n349), .Y(n288) );
  NOR2X4 U219 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U220 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U221 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U222 ( .A(n347), .Y(n1) );
  CLKINVX3 U223 ( .A(a[2]), .Y(n273) );
  OAI21X1 U224 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U225 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U226 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U227 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U228 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U229 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  AOI31X4 U230 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  CLKINVX3 U231 ( .A(n309), .Y(n345) );
  NAND2X2 U232 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U233 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U234 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U235 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U236 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U237 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U238 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U239 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U240 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U241 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U242 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U243 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U244 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U245 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U246 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U247 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U248 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U249 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U250 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U251 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U252 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U253 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U254 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U255 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U256 ( .A(a[1]), .Y(n323) );
  NAND2X1 U257 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U258 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U259 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U260 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U261 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U262 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U263 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U264 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U265 ( .A(n242), .Y(n249) );
  OAI21XL U266 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U267 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U268 ( .A(n192), .Y(n205) );
  INVX1 U269 ( .A(n66), .Y(n111) );
  NOR2X1 U270 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U271 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U272 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U273 ( .A(a[6]), .B(a[0]), .Y(n360) );
  NOR2X1 U274 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U275 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U276 ( .A(n261), .Y(n307) );
  INVX1 U277 ( .A(n20), .Y(n326) );
  NAND2X1 U278 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U279 ( .A(n187), .Y(n196) );
  INVX1 U280 ( .A(n350), .Y(n335) );
  NAND2X1 U281 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U282 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U283 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U284 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U285 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U286 ( .A(n103), .Y(n37) );
  NOR2X1 U287 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U288 ( .A(n311), .Y(n268) );
  AOI22X1 U289 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  INVX1 U290 ( .A(n293), .Y(n209) );
  NOR2X1 U291 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U292 ( .A(n224), .Y(n235) );
  NAND2X1 U293 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U294 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U295 ( .A(n195), .Y(n142) );
  NAND2X1 U296 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U297 ( .A(n226), .Y(n253) );
  NAND2X1 U298 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U299 ( .A(n140), .B(n20), .Y(n151) );
  NAND2X1 U300 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U301 ( .A(n1), .Y(n301) );
  NAND2X1 U302 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U303 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U304 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U305 ( .A(n89), .Y(n340) );
  AOI211X1 U306 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U307 ( .A(n327), .Y(n248) );
  INVX1 U308 ( .A(n181), .Y(n109) );
  INVX1 U309 ( .A(n225), .Y(n302) );
  NAND2X1 U310 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U311 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U312 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U313 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U314 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U315 ( .A(n270), .Y(n107) );
  INVX1 U316 ( .A(n306), .Y(n145) );
  NAND4X1 U317 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U318 ( .A(n210), .Y(n236) );
  INVX1 U319 ( .A(n331), .Y(n78) );
  INVX1 U320 ( .A(n328), .Y(n314) );
  OAI21XL U321 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U322 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U323 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U324 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_11 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  AOI21XL U4 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  INVX1 U5 ( .A(n116), .Y(n203) );
  NAND2X1 U6 ( .A(n194), .B(n274), .Y(n344) );
  NAND2XL U7 ( .A(n140), .B(n20), .Y(n151) );
  INVX1 U8 ( .A(n324), .Y(n265) );
  AOI211XL U9 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  AOI2BB2XL U10 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI21XL U11 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  INVXL U12 ( .A(n257), .Y(n289) );
  NAND2XL U13 ( .A(n235), .B(n265), .Y(n338) );
  NOR2XL U14 ( .A(n224), .B(n326), .Y(n257) );
  INVXL U15 ( .A(n150), .Y(n310) );
  AOI22XL U16 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NOR2XL U17 ( .A(n248), .B(n142), .Y(n357) );
  NAND2XL U18 ( .A(n109), .B(n78), .Y(n158) );
  NOR2X1 U19 ( .A(a[1]), .B(n293), .Y(n318) );
  NOR2X1 U20 ( .A(n293), .B(n323), .Y(n150) );
  NOR2XL U21 ( .A(n181), .B(n95), .Y(n174) );
  NOR2XL U22 ( .A(n324), .B(n131), .Y(n262) );
  NAND2XL U23 ( .A(a[1]), .B(n293), .Y(n82) );
  INVXL U24 ( .A(n352), .Y(n141) );
  NOR2X4 U25 ( .A(n264), .B(n197), .Y(n350) );
  NOR2X1 U26 ( .A(a[1]), .B(n103), .Y(n331) );
  INVXL U27 ( .A(n267), .Y(n333) );
  NOR2XL U28 ( .A(a[1]), .B(n242), .Y(n186) );
  NAND2X1 U29 ( .A(a[1]), .B(n31), .Y(n352) );
  OR4X2 U30 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U31 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U32 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI211XL U33 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  AOI31XL U34 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI31XL U35 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI211XL U36 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U37 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U38 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI31XL U39 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  OAI211XL U40 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U41 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI31XL U42 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI211XL U43 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI22XL U44 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  AOI31XL U45 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U46 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI211XL U47 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI211XL U48 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U49 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI31XL U50 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI22XL U51 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI22XL U52 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  OAI211XL U53 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI31XL U54 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  OAI22XL U55 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI31XL U56 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  OAI211XL U57 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI211XL U58 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI211XL U59 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  OAI211XL U60 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U61 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI22XL U62 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U63 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U64 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  AOI31XL U65 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  INVXL U66 ( .A(n101), .Y(n254) );
  AOI31XL U67 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  NAND2XL U68 ( .A(n296), .B(n101), .Y(n94) );
  AOI211XL U69 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  OAI211XL U70 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  AOI221XL U71 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI211XL U72 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  NOR2XL U73 ( .A(n150), .B(n331), .Y(n130) );
  OAI211XL U74 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  AOI22XL U75 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  NAND2XL U76 ( .A(n235), .B(n274), .Y(n184) );
  AOI31XL U77 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  NOR2XL U78 ( .A(n224), .B(n150), .Y(n116) );
  AOI31XL U79 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  AOI22XL U80 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI22XL U81 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  AOI211XL U82 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI211XL U83 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI31XL U84 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI22XL U85 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI22XL U86 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI22XL U87 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI2BB2XL U88 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI211XL U89 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI22XL U90 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI211XL U91 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI22XL U92 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI22XL U93 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI2BB2XL U94 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U95 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI22XL U96 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI22XL U97 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI2BB2XL U98 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI211XL U99 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI211XL U100 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI31XL U101 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI211XL U102 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  INVXL U103 ( .A(n152), .Y(n222) );
  NAND2XL U104 ( .A(n265), .B(n348), .Y(n247) );
  AOI211XL U105 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI22XL U106 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  OAI22XL U107 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  NOR2XL U108 ( .A(n161), .B(n309), .Y(n162) );
  NAND2XL U109 ( .A(n109), .B(n242), .Y(n135) );
  AOI22XL U110 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  AOI211XL U111 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  INVXL U112 ( .A(n312), .Y(n313) );
  AOI22XL U113 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI22XL U114 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  AOI22XL U115 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  NAND3XL U116 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  NAND2XL U117 ( .A(n352), .B(n351), .Y(n358) );
  OAI22XL U118 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  AOI22XL U119 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  AOI22XL U120 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  AOI22XL U121 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  OAI22XL U122 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI2BB2XL U123 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U124 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  NOR2XL U125 ( .A(n293), .B(n292), .Y(n294) );
  AOI22XL U126 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  NAND2XL U127 ( .A(n103), .B(n253), .Y(n305) );
  AOI22XL U128 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  AOI2BB2XL U129 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  AOI22XL U130 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI22XL U131 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  OAI211XL U132 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  OAI2BB1XL U133 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  NOR2XL U134 ( .A(n209), .B(n233), .Y(n256) );
  AOI32XL U135 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  INVXL U136 ( .A(n180), .Y(n183) );
  INVXL U137 ( .A(n82), .Y(n172) );
  AOI211XL U138 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  OAI22XL U139 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI22XL U140 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  AOI22XL U141 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  NOR2XL U142 ( .A(n37), .B(n145), .Y(n99) );
  AOI31XL U143 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI22XL U144 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  AOI22XL U145 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  AOI211XL U146 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  AOI22XL U147 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  NOR2XL U148 ( .A(n268), .B(n354), .Y(n13) );
  AOI22XL U149 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  AOI22XL U150 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  NAND2XL U151 ( .A(n311), .B(n196), .Y(n40) );
  NOR2XL U152 ( .A(n293), .B(n226), .Y(n39) );
  NOR2XL U153 ( .A(n181), .B(n269), .Y(n315) );
  AOI22XL U154 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AOI22XL U155 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  NOR3XL U156 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  NOR3XL U157 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI22XL U158 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  NAND2XL U159 ( .A(n311), .B(n236), .Y(n346) );
  AOI22XL U160 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  AOI2BB2XL U161 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U162 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  NAND2XL U163 ( .A(n350), .B(n245), .Y(n180) );
  AOI22XL U164 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  OAI22XL U165 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U166 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AND2X2 U167 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U168 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  INVXL U169 ( .A(n131), .Y(n351) );
  AOI22XL U170 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  AOI22XL U171 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NAND2XL U172 ( .A(n306), .B(n267), .Y(n61) );
  NAND3XL U173 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  AOI22XL U174 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  NAND2XL U175 ( .A(n329), .B(n323), .Y(n245) );
  NOR2XL U176 ( .A(n37), .B(a[1]), .Y(n195) );
  AOI22XL U177 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  NAND2XL U178 ( .A(n311), .B(n303), .Y(n38) );
  NAND2XL U179 ( .A(n107), .B(n348), .Y(n175) );
  NOR2XL U180 ( .A(n187), .B(n186), .Y(n290) );
  NOR2XL U181 ( .A(n233), .B(n331), .Y(n108) );
  NAND3XL U182 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  NOR2XL U183 ( .A(a[1]), .B(n249), .Y(n131) );
  NOR2XL U184 ( .A(a[1]), .B(n329), .Y(n269) );
  AOI22XL U185 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  AOI22XL U186 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  INVXL U187 ( .A(n332), .Y(n234) );
  NAND2XL U188 ( .A(a[1]), .B(n261), .Y(n303) );
  NAND2XL U189 ( .A(n328), .B(n311), .Y(n353) );
  INVXL U190 ( .A(n197), .Y(n185) );
  INVXL U191 ( .A(n297), .Y(n284) );
  NAND3XL U192 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  AOI22XL U193 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  AOI22XL U194 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U195 ( .A(a[1]), .B(n198), .Y(n160) );
  INVXL U196 ( .A(n274), .Y(n251) );
  NOR2XL U197 ( .A(n264), .B(n273), .Y(n330) );
  NAND2XL U198 ( .A(n264), .B(n275), .Y(n252) );
  NOR2XL U199 ( .A(a[3]), .B(a[1]), .Y(n225) );
  NAND2XL U200 ( .A(a[4]), .B(a[1]), .Y(n274) );
  INVX2 U201 ( .A(a[7]), .Y(n264) );
  NAND2XL U202 ( .A(a[3]), .B(a[1]), .Y(n20) );
  CLKINVX3 U203 ( .A(n266), .Y(n329) );
  NAND2X2 U204 ( .A(a[4]), .B(n31), .Y(n266) );
  NAND2X2 U205 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U206 ( .A(a[5]), .Y(n275) );
  OAI21X1 U207 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U208 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U209 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NOR2X2 U210 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U211 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U212 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U213 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U214 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U215 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U216 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U217 ( .A(n233), .Y(n359) );
  NAND2X2 U218 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U219 ( .A(n349), .Y(n288) );
  NOR2X4 U220 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U221 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U222 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U223 ( .A(n347), .Y(n1) );
  CLKINVX3 U224 ( .A(a[2]), .Y(n273) );
  OAI21X1 U225 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U226 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U227 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U228 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U229 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U230 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  AOI31X4 U231 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  CLKINVX3 U232 ( .A(n309), .Y(n345) );
  NAND2X2 U233 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U234 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U235 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U236 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U237 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U238 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U239 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U240 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U241 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U242 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U243 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U244 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U245 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U246 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U247 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U248 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U249 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U250 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U251 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U252 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U253 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U254 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U255 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U256 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U257 ( .A(a[1]), .Y(n323) );
  NAND2X1 U258 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U259 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U260 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U261 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U262 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U263 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U264 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U265 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U266 ( .A(n242), .Y(n249) );
  OAI21XL U267 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U268 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U269 ( .A(n192), .Y(n205) );
  INVX1 U270 ( .A(n66), .Y(n111) );
  NOR2X1 U271 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U272 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U273 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U274 ( .A(a[6]), .B(a[0]), .Y(n360) );
  INVX1 U275 ( .A(a[6]), .Y(n16) );
  NOR2X1 U276 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U277 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U278 ( .A(n261), .Y(n307) );
  INVX1 U279 ( .A(n20), .Y(n326) );
  NAND2X1 U280 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U281 ( .A(n187), .Y(n196) );
  INVX1 U282 ( .A(n350), .Y(n335) );
  NAND2X1 U283 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U284 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U285 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U286 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U287 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U288 ( .A(n103), .Y(n37) );
  NOR2X1 U289 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U290 ( .A(n311), .Y(n268) );
  INVX1 U291 ( .A(n293), .Y(n209) );
  NOR2X1 U292 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U293 ( .A(n224), .Y(n235) );
  NAND2X1 U294 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U295 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U296 ( .A(n195), .Y(n142) );
  NAND2X1 U297 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U298 ( .A(n226), .Y(n253) );
  NAND2X1 U299 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U300 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U301 ( .A(n1), .Y(n301) );
  NAND2X1 U302 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U303 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U304 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U305 ( .A(n89), .Y(n340) );
  AOI211X1 U306 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U307 ( .A(n327), .Y(n248) );
  INVX1 U308 ( .A(n181), .Y(n109) );
  INVX1 U309 ( .A(n225), .Y(n302) );
  NAND2X1 U310 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U311 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U312 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U313 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U314 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U315 ( .A(n270), .Y(n107) );
  INVX1 U316 ( .A(n306), .Y(n145) );
  NAND4X1 U317 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U318 ( .A(n210), .Y(n236) );
  INVX1 U319 ( .A(n331), .Y(n78) );
  INVX1 U320 ( .A(n328), .Y(n314) );
  OAI21XL U321 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U322 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U323 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U324 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_12 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  AOI211XL U4 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  INVX1 U5 ( .A(n116), .Y(n203) );
  NAND2XL U6 ( .A(n140), .B(n20), .Y(n151) );
  NAND2X1 U7 ( .A(n194), .B(n274), .Y(n344) );
  INVX1 U8 ( .A(n324), .Y(n265) );
  AOI21XL U9 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  INVXL U10 ( .A(n257), .Y(n289) );
  NAND2XL U11 ( .A(n235), .B(n265), .Y(n338) );
  OAI211XL U12 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  NOR2XL U13 ( .A(n224), .B(n326), .Y(n257) );
  AOI22XL U14 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NOR2XL U15 ( .A(n248), .B(n142), .Y(n357) );
  NAND2XL U16 ( .A(n109), .B(n78), .Y(n158) );
  NAND2XL U17 ( .A(a[1]), .B(n293), .Y(n82) );
  NOR2X1 U18 ( .A(a[1]), .B(n293), .Y(n318) );
  NOR2X1 U19 ( .A(n293), .B(n323), .Y(n150) );
  NOR2XL U20 ( .A(n324), .B(n131), .Y(n262) );
  NOR2X1 U21 ( .A(a[1]), .B(n103), .Y(n331) );
  NOR2X4 U22 ( .A(n264), .B(n197), .Y(n350) );
  INVXL U23 ( .A(n352), .Y(n141) );
  NOR2XL U24 ( .A(a[1]), .B(n242), .Y(n186) );
  NAND2X1 U25 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI211XL U26 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI31XL U27 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI211XL U28 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI211XL U29 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  OR4X2 U30 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI31XL U31 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U32 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  OAI211XL U33 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U34 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI31XL U35 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI211XL U36 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U37 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U38 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI211XL U39 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI211XL U40 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI31XL U41 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  AOI211XL U42 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI31XL U43 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  OAI211XL U44 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI22XL U45 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI22XL U46 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  OAI22XL U47 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI22XL U48 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  AOI31XL U49 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI211XL U50 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI31XL U51 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI21X1 U52 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  OAI211XL U53 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI211XL U54 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U55 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  INVXL U56 ( .A(n101), .Y(n254) );
  OAI211XL U57 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI22XL U58 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U59 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI211XL U60 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  AOI2BB2XL U61 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI211XL U62 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  NAND2XL U63 ( .A(n296), .B(n101), .Y(n94) );
  AOI31XL U64 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  AOI211XL U65 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U66 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI31XL U67 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  AOI22XL U68 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI31XL U69 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  NAND2XL U70 ( .A(n235), .B(n274), .Y(n184) );
  AOI211XL U71 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  AOI221XL U72 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI211XL U73 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI31XL U74 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI22XL U75 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  AOI22XL U76 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  OAI211XL U77 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  INVXL U78 ( .A(n150), .Y(n310) );
  NOR2XL U79 ( .A(n150), .B(n331), .Y(n130) );
  AOI211XL U80 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI31XL U81 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  NOR2XL U82 ( .A(n224), .B(n150), .Y(n116) );
  AOI22XL U83 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI22XL U84 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  NAND2XL U85 ( .A(n265), .B(n348), .Y(n247) );
  AOI22XL U86 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI22XL U87 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI22XL U88 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI211XL U89 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI2BB2XL U90 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI22XL U91 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI22XL U92 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  INVXL U93 ( .A(n152), .Y(n222) );
  AOI211XL U94 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI2BB2XL U95 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI211XL U96 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI22XL U97 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI2BB2XL U98 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U99 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI211XL U100 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI31XL U101 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI211XL U102 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  OAI22XL U103 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI211XL U104 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI22XL U105 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI22XL U106 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  AOI22XL U107 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  NAND2XL U108 ( .A(n109), .B(n242), .Y(n135) );
  AOI22XL U109 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  NOR2XL U110 ( .A(n161), .B(n309), .Y(n162) );
  OAI22XL U111 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI2BB2XL U112 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U113 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI22XL U114 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  AOI211XL U115 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI22XL U116 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI22XL U117 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  NAND3XL U118 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  OAI22XL U119 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  NAND2XL U120 ( .A(n352), .B(n351), .Y(n358) );
  NOR2XL U121 ( .A(n293), .B(n292), .Y(n294) );
  NAND2XL U122 ( .A(n103), .B(n253), .Y(n305) );
  AOI22XL U123 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  INVXL U124 ( .A(n312), .Y(n313) );
  OAI211XL U125 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U126 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI2BB2XL U127 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  NOR2XL U128 ( .A(n209), .B(n233), .Y(n256) );
  AOI22XL U129 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  AOI22XL U130 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  AOI211XL U131 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  INVXL U132 ( .A(n180), .Y(n183) );
  AOI32XL U133 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  INVXL U134 ( .A(n82), .Y(n172) );
  AOI22XL U135 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  OAI2BB1XL U136 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  AOI22XL U137 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  NOR2XL U138 ( .A(n293), .B(n226), .Y(n39) );
  AOI22XL U139 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  NAND2XL U140 ( .A(n311), .B(n196), .Y(n40) );
  NOR2XL U141 ( .A(n37), .B(n145), .Y(n99) );
  AOI22XL U142 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  AOI22XL U143 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  OAI22XL U144 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI2BB2XL U145 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  NOR2XL U146 ( .A(n181), .B(n269), .Y(n315) );
  AOI22XL U147 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  AOI31XL U148 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI22XL U149 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  NOR2XL U150 ( .A(n268), .B(n354), .Y(n13) );
  AOI211XL U151 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  AOI22XL U152 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  AOI22XL U153 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  AOI22XL U154 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI22XL U155 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  INVXL U156 ( .A(n131), .Y(n351) );
  AOI22XL U157 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  NOR3XL U158 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI22XL U159 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  NAND2XL U160 ( .A(n350), .B(n245), .Y(n180) );
  AOI22XL U161 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  NOR3XL U162 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  NAND2XL U163 ( .A(n311), .B(n236), .Y(n346) );
  OAI22XL U164 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U165 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  AOI22XL U166 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AND2X2 U167 ( .A(n303), .B(n78), .Y(n221) );
  NAND2XL U168 ( .A(n306), .B(n267), .Y(n61) );
  AOI22XL U169 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NAND3XL U170 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  AOI22XL U171 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  AOI22XL U172 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  NAND2XL U173 ( .A(n311), .B(n303), .Y(n38) );
  AOI22XL U174 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  AOI22XL U175 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NOR2XL U176 ( .A(a[1]), .B(n249), .Y(n131) );
  NOR2XL U177 ( .A(a[1]), .B(n329), .Y(n269) );
  NAND3XL U178 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NAND2XL U179 ( .A(n329), .B(n323), .Y(n245) );
  NOR2XL U180 ( .A(n233), .B(n331), .Y(n108) );
  AOI22XL U181 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  NOR2XL U182 ( .A(n37), .B(a[1]), .Y(n195) );
  NOR2XL U183 ( .A(n187), .B(n186), .Y(n290) );
  NAND2XL U184 ( .A(n107), .B(n348), .Y(n175) );
  INVXL U185 ( .A(n197), .Y(n185) );
  NAND2XL U186 ( .A(n328), .B(n311), .Y(n353) );
  NAND2XL U187 ( .A(a[1]), .B(n261), .Y(n303) );
  INVXL U188 ( .A(n297), .Y(n284) );
  INVXL U189 ( .A(n332), .Y(n234) );
  NAND3XL U190 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  INVXL U191 ( .A(n267), .Y(n333) );
  INVXL U192 ( .A(n274), .Y(n251) );
  AOI22XL U193 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U194 ( .A(n264), .B(n273), .Y(n330) );
  NOR2XL U195 ( .A(a[1]), .B(n198), .Y(n160) );
  AOI22XL U196 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  NAND2XL U197 ( .A(n264), .B(n275), .Y(n252) );
  NAND2XL U198 ( .A(a[3]), .B(a[1]), .Y(n20) );
  INVX2 U199 ( .A(a[7]), .Y(n264) );
  NAND2XL U200 ( .A(a[4]), .B(a[1]), .Y(n274) );
  NOR2XL U201 ( .A(a[3]), .B(a[1]), .Y(n225) );
  CLKINVX3 U202 ( .A(n266), .Y(n329) );
  NAND2X2 U203 ( .A(a[4]), .B(n31), .Y(n266) );
  OAI21X1 U204 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U205 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U206 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U207 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U208 ( .A(a[5]), .Y(n275) );
  NOR2X2 U209 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U210 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U211 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U212 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U213 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U214 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U215 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U216 ( .A(n233), .Y(n359) );
  NAND2X2 U217 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U218 ( .A(n349), .Y(n288) );
  NOR2X4 U219 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U220 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U221 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U222 ( .A(n347), .Y(n1) );
  CLKINVX3 U223 ( .A(a[2]), .Y(n273) );
  OAI21X1 U224 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U225 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U226 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U227 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U228 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U229 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31X4 U230 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  CLKINVX3 U231 ( .A(n309), .Y(n345) );
  NAND2X2 U232 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U233 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U234 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U235 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U236 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U237 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U238 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U239 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U240 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U241 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U242 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U243 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U244 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U245 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U246 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U247 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U248 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U249 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U250 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U251 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U252 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U253 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U254 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U255 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U256 ( .A(a[1]), .Y(n323) );
  NAND2X1 U257 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U258 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U259 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U260 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U261 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U262 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U263 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U264 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U265 ( .A(n242), .Y(n249) );
  OAI21XL U266 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U267 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U268 ( .A(n192), .Y(n205) );
  INVX1 U269 ( .A(n66), .Y(n111) );
  NOR2X1 U270 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U271 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U272 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U273 ( .A(a[6]), .B(a[0]), .Y(n360) );
  INVX1 U274 ( .A(a[6]), .Y(n16) );
  NOR2X1 U275 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U276 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U277 ( .A(n261), .Y(n307) );
  INVX1 U278 ( .A(n20), .Y(n326) );
  NAND2X1 U279 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U280 ( .A(n187), .Y(n196) );
  INVX1 U281 ( .A(n350), .Y(n335) );
  NAND2X1 U282 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U283 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U284 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U285 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U286 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U287 ( .A(n103), .Y(n37) );
  NOR2X1 U288 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U289 ( .A(n311), .Y(n268) );
  INVX1 U290 ( .A(n293), .Y(n209) );
  NOR2X1 U291 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U292 ( .A(n224), .Y(n235) );
  NAND2X1 U293 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U294 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U295 ( .A(n195), .Y(n142) );
  NAND2X1 U296 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U297 ( .A(n226), .Y(n253) );
  NAND2X1 U298 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U299 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U300 ( .A(n1), .Y(n301) );
  NAND2X1 U301 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U302 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U303 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U304 ( .A(n89), .Y(n340) );
  AOI211X1 U305 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U306 ( .A(n327), .Y(n248) );
  INVX1 U307 ( .A(n181), .Y(n109) );
  INVX1 U308 ( .A(n225), .Y(n302) );
  NAND2X1 U309 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U310 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U311 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U312 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U313 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U314 ( .A(n270), .Y(n107) );
  INVX1 U315 ( .A(n306), .Y(n145) );
  NAND4X1 U316 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U317 ( .A(n210), .Y(n236) );
  INVX1 U318 ( .A(n331), .Y(n78) );
  INVX1 U319 ( .A(n328), .Y(n314) );
  OAI21XL U320 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U321 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U322 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U323 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  NOR2X1 U324 ( .A(n181), .B(n95), .Y(n174) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_13 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  AOI211XL U4 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  INVX1 U5 ( .A(n116), .Y(n203) );
  NAND2X1 U6 ( .A(n194), .B(n274), .Y(n344) );
  NAND2X1 U7 ( .A(n140), .B(n20), .Y(n151) );
  INVX1 U8 ( .A(n324), .Y(n265) );
  AOI21XL U9 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  OAI211XL U10 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  INVXL U11 ( .A(n257), .Y(n289) );
  NAND2XL U12 ( .A(n235), .B(n265), .Y(n338) );
  NOR2XL U13 ( .A(n224), .B(n326), .Y(n257) );
  NAND2XL U14 ( .A(n109), .B(n78), .Y(n158) );
  AOI22XL U15 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NOR2XL U16 ( .A(n248), .B(n142), .Y(n357) );
  NOR2X1 U17 ( .A(n293), .B(n323), .Y(n150) );
  NOR2X1 U18 ( .A(a[1]), .B(n293), .Y(n318) );
  NAND2XL U19 ( .A(a[1]), .B(n293), .Y(n82) );
  NOR2XL U20 ( .A(n324), .B(n131), .Y(n262) );
  INVXL U21 ( .A(n352), .Y(n141) );
  INVXL U22 ( .A(n267), .Y(n333) );
  NOR2X1 U23 ( .A(a[1]), .B(n103), .Y(n331) );
  NOR2XL U24 ( .A(a[1]), .B(n242), .Y(n186) );
  NOR2X4 U25 ( .A(n264), .B(n197), .Y(n350) );
  NAND2X1 U26 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI211XL U27 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI211XL U28 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  OR4X2 U29 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI31XL U30 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI211XL U31 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U32 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U33 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI31XL U34 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U35 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U36 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI31XL U37 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  OAI211XL U38 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U39 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  OAI211XL U40 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI211XL U41 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI22XL U42 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  OAI211XL U43 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  OAI22XL U44 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI211XL U45 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U46 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI21X1 U47 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  AOI211XL U48 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI22XL U49 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI22XL U50 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI211XL U51 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI31XL U52 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI31XL U53 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI31XL U54 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI31XL U55 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  AOI211XL U56 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI211XL U57 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  NAND2XL U58 ( .A(n296), .B(n101), .Y(n94) );
  AOI211XL U59 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  AOI31XL U60 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  INVXL U61 ( .A(n101), .Y(n254) );
  AOI31XL U62 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  OAI211XL U63 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI2BB2XL U64 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI211XL U65 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  AOI211XL U66 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U67 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI22XL U68 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  OAI211XL U69 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  AOI22XL U70 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  AOI31XL U71 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI22XL U72 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI211XL U73 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI22XL U74 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  INVXL U75 ( .A(n150), .Y(n310) );
  AOI211XL U76 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  NAND2XL U77 ( .A(n235), .B(n274), .Y(n184) );
  AOI211XL U78 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  NOR2XL U79 ( .A(n224), .B(n150), .Y(n116) );
  AOI31XL U80 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI31XL U81 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  NOR2XL U82 ( .A(n150), .B(n331), .Y(n130) );
  AOI221XL U83 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI22XL U84 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  INVXL U85 ( .A(n152), .Y(n222) );
  AOI22XL U86 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI2BB2XL U87 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI211XL U88 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI22XL U89 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI2BB2XL U90 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI22XL U91 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  NAND2XL U92 ( .A(n265), .B(n348), .Y(n247) );
  AOI2BB2XL U93 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI211XL U94 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI211XL U95 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI211XL U96 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI211XL U97 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI31XL U98 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI22XL U99 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI22XL U100 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI22XL U101 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI22XL U102 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI211XL U103 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  OAI22XL U104 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI22XL U105 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI22XL U106 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI22XL U107 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  NAND2XL U108 ( .A(n109), .B(n242), .Y(n135) );
  AOI22XL U109 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  AOI22XL U110 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  AOI22XL U111 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI211XL U112 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI2BB2XL U113 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U114 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI22XL U115 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  AOI22XL U116 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  OAI22XL U117 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  NAND3XL U118 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  AOI22XL U119 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  OAI22XL U120 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI22XL U121 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  AOI22XL U122 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  OAI2BB1XL U123 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  INVXL U124 ( .A(n312), .Y(n313) );
  NAND2XL U125 ( .A(n103), .B(n253), .Y(n305) );
  NOR2XL U126 ( .A(n293), .B(n292), .Y(n294) );
  OAI211XL U127 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U128 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  NOR2XL U129 ( .A(n209), .B(n233), .Y(n256) );
  AOI2BB2XL U130 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  INVXL U131 ( .A(n82), .Y(n172) );
  AOI32XL U132 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  NOR2XL U133 ( .A(n161), .B(n309), .Y(n162) );
  INVXL U134 ( .A(n180), .Y(n183) );
  AOI211XL U135 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  NAND2XL U136 ( .A(n352), .B(n351), .Y(n358) );
  AOI22XL U137 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  AOI22XL U138 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  NOR2XL U139 ( .A(n293), .B(n226), .Y(n39) );
  AOI22XL U140 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  NAND2XL U141 ( .A(n311), .B(n196), .Y(n40) );
  AOI22XL U142 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AOI22XL U143 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  INVXL U144 ( .A(n131), .Y(n351) );
  AOI22XL U145 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AOI22XL U146 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  OAI22XL U147 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U148 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  NOR2XL U149 ( .A(n268), .B(n354), .Y(n13) );
  NAND2XL U150 ( .A(n311), .B(n236), .Y(n346) );
  AOI22XL U151 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  NAND2XL U152 ( .A(n350), .B(n245), .Y(n180) );
  AND2X2 U153 ( .A(n303), .B(n78), .Y(n221) );
  NOR3XL U154 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  NOR2XL U155 ( .A(n37), .B(n145), .Y(n99) );
  AOI22XL U156 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  AOI22XL U157 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI22XL U158 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  OAI22XL U159 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  NOR3XL U160 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  AOI22XL U161 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  AOI22XL U162 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  AOI22XL U163 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  AOI211XL U164 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  NOR2XL U165 ( .A(n181), .B(n269), .Y(n315) );
  AOI31XL U166 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI2BB2XL U167 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U168 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  NAND2XL U169 ( .A(n329), .B(n323), .Y(n245) );
  AOI22XL U170 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NAND2XL U171 ( .A(n306), .B(n267), .Y(n61) );
  NAND2XL U172 ( .A(n311), .B(n303), .Y(n38) );
  NOR2XL U173 ( .A(n187), .B(n186), .Y(n290) );
  NAND2XL U174 ( .A(n107), .B(n348), .Y(n175) );
  NOR2XL U175 ( .A(n233), .B(n331), .Y(n108) );
  NAND3XL U176 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  AOI22XL U177 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  AOI22XL U178 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  AOI22XL U179 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  NAND3XL U180 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NOR2XL U181 ( .A(n37), .B(a[1]), .Y(n195) );
  AOI22XL U182 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  NOR2XL U183 ( .A(a[1]), .B(n329), .Y(n269) );
  AOI22XL U184 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  NOR2XL U185 ( .A(a[1]), .B(n249), .Y(n131) );
  INVXL U186 ( .A(n197), .Y(n185) );
  NAND3XL U187 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  NAND2XL U188 ( .A(a[1]), .B(n261), .Y(n303) );
  NAND2XL U189 ( .A(n328), .B(n311), .Y(n353) );
  INVXL U190 ( .A(n297), .Y(n284) );
  INVXL U191 ( .A(n332), .Y(n234) );
  NOR2XL U192 ( .A(n264), .B(n273), .Y(n330) );
  NAND2XL U193 ( .A(n264), .B(n275), .Y(n252) );
  INVXL U194 ( .A(n274), .Y(n251) );
  AOI22XL U195 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  NOR2XL U196 ( .A(a[1]), .B(n198), .Y(n160) );
  AOI22XL U197 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U198 ( .A(a[3]), .B(a[1]), .Y(n225) );
  INVX2 U199 ( .A(a[7]), .Y(n264) );
  NAND2XL U200 ( .A(a[3]), .B(a[1]), .Y(n20) );
  NAND2XL U201 ( .A(a[4]), .B(a[1]), .Y(n274) );
  CLKINVX3 U202 ( .A(n266), .Y(n329) );
  NAND2X2 U203 ( .A(a[4]), .B(n31), .Y(n266) );
  OAI21X1 U204 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U205 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U206 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U207 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U208 ( .A(a[5]), .Y(n275) );
  NOR2X2 U209 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U210 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U211 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U212 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U213 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U214 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U215 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U216 ( .A(n233), .Y(n359) );
  NAND2X2 U217 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U218 ( .A(n349), .Y(n288) );
  NOR2X4 U219 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U220 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U221 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U222 ( .A(n347), .Y(n1) );
  CLKINVX3 U223 ( .A(a[2]), .Y(n273) );
  OAI21X1 U224 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U225 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U226 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U227 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U228 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U229 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31X4 U230 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  CLKINVX3 U231 ( .A(n309), .Y(n345) );
  NAND2X2 U232 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U233 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U234 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U235 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U236 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U237 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U238 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U239 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U240 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U241 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U242 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U243 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U244 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U245 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U246 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U247 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U248 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U249 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U250 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U251 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U252 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U253 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U254 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U255 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U256 ( .A(a[1]), .Y(n323) );
  NAND2X1 U257 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U258 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U259 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U260 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U261 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U262 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U263 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U264 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U265 ( .A(n242), .Y(n249) );
  OAI21XL U266 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U267 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U268 ( .A(n192), .Y(n205) );
  INVX1 U269 ( .A(n66), .Y(n111) );
  NOR2X1 U270 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U271 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U272 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U273 ( .A(a[6]), .B(a[0]), .Y(n360) );
  INVX1 U274 ( .A(a[6]), .Y(n16) );
  NOR2X1 U275 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U276 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U277 ( .A(n261), .Y(n307) );
  INVX1 U278 ( .A(n20), .Y(n326) );
  NAND2X1 U279 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U280 ( .A(n187), .Y(n196) );
  INVX1 U281 ( .A(n350), .Y(n335) );
  NAND2X1 U282 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U283 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U284 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U285 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U286 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U287 ( .A(n103), .Y(n37) );
  NOR2X1 U288 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U289 ( .A(n311), .Y(n268) );
  INVX1 U290 ( .A(n293), .Y(n209) );
  NOR2X1 U291 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U292 ( .A(n224), .Y(n235) );
  NAND2X1 U293 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U294 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U295 ( .A(n195), .Y(n142) );
  NAND2X1 U296 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U297 ( .A(n226), .Y(n253) );
  NAND2X1 U298 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U299 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U300 ( .A(n1), .Y(n301) );
  NAND2X1 U301 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U302 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U303 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U304 ( .A(n89), .Y(n340) );
  AOI211X1 U305 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U306 ( .A(n327), .Y(n248) );
  INVX1 U307 ( .A(n181), .Y(n109) );
  INVX1 U308 ( .A(n225), .Y(n302) );
  NAND2X1 U309 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U310 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U311 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U312 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U313 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U314 ( .A(n270), .Y(n107) );
  INVX1 U315 ( .A(n306), .Y(n145) );
  NAND4X1 U316 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U317 ( .A(n210), .Y(n236) );
  INVX1 U318 ( .A(n331), .Y(n78) );
  INVX1 U319 ( .A(n328), .Y(n314) );
  OAI21XL U320 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U321 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U322 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U323 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  NOR2X1 U324 ( .A(n181), .B(n95), .Y(n174) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_14 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  AOI211XL U4 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  INVX1 U5 ( .A(n116), .Y(n203) );
  NAND2X1 U6 ( .A(n194), .B(n274), .Y(n344) );
  NAND2XL U7 ( .A(n140), .B(n20), .Y(n151) );
  INVX1 U8 ( .A(n324), .Y(n265) );
  AOI21XL U9 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  NAND2XL U10 ( .A(n235), .B(n265), .Y(n338) );
  OAI211XL U11 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  INVXL U12 ( .A(n257), .Y(n289) );
  NOR2XL U13 ( .A(n224), .B(n326), .Y(n257) );
  NAND2XL U14 ( .A(n109), .B(n78), .Y(n158) );
  NOR2XL U15 ( .A(n248), .B(n142), .Y(n357) );
  AOI22XL U16 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NOR2XL U17 ( .A(n324), .B(n131), .Y(n262) );
  NAND2XL U18 ( .A(a[1]), .B(n293), .Y(n82) );
  NOR2X1 U19 ( .A(a[1]), .B(n293), .Y(n318) );
  NOR2X1 U20 ( .A(n293), .B(n323), .Y(n150) );
  NOR2X4 U21 ( .A(n264), .B(n197), .Y(n350) );
  NOR2XL U22 ( .A(a[1]), .B(n242), .Y(n186) );
  NOR2X1 U23 ( .A(a[1]), .B(n103), .Y(n331) );
  INVXL U24 ( .A(n267), .Y(n333) );
  INVXL U25 ( .A(n352), .Y(n141) );
  NAND2X1 U26 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI31XL U27 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI211XL U28 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  AOI211XL U29 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI211XL U30 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  OR4X2 U31 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI31XL U32 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI211XL U33 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U34 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U35 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI31XL U36 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  OAI211XL U37 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U38 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U39 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  OAI22XL U40 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  OAI211XL U41 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI22XL U42 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  AOI211XL U43 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U44 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  OAI211XL U45 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI31XL U46 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U47 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI31XL U48 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  AOI211XL U49 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI31XL U50 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI31XL U51 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI22XL U52 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI211XL U53 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI211XL U54 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI22XL U55 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI21X1 U56 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  NAND2XL U57 ( .A(n296), .B(n101), .Y(n94) );
  AOI31XL U58 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  AOI22XL U59 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U60 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  AOI211XL U61 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  OAI211XL U62 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U63 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U64 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  AOI2BB2XL U65 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI31XL U66 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  INVXL U67 ( .A(n101), .Y(n254) );
  AOI211XL U68 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI31XL U69 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI31XL U70 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI211XL U71 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI22XL U72 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  OAI211XL U73 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  AOI22XL U74 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  INVXL U75 ( .A(n150), .Y(n310) );
  NOR2XL U76 ( .A(n150), .B(n331), .Y(n130) );
  NAND2XL U77 ( .A(n235), .B(n274), .Y(n184) );
  AOI211XL U78 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  AOI22XL U79 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  AOI211XL U80 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  NOR2XL U81 ( .A(n224), .B(n150), .Y(n116) );
  AOI31XL U82 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  AOI221XL U83 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI2BB2XL U84 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI31XL U85 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI2BB2XL U86 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI211XL U87 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI211XL U88 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  OAI22XL U89 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  INVXL U90 ( .A(n152), .Y(n222) );
  AOI22XL U91 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI211XL U92 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  NAND2XL U93 ( .A(n265), .B(n348), .Y(n247) );
  AOI22XL U94 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI22XL U95 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI211XL U96 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI22XL U97 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI22XL U98 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI22XL U99 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI2BB2XL U100 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U101 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI22XL U102 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI211XL U103 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI211XL U104 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI22XL U105 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI22XL U106 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  NAND2XL U107 ( .A(n109), .B(n242), .Y(n135) );
  OAI211XL U108 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U109 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  NOR2XL U110 ( .A(n209), .B(n233), .Y(n256) );
  NAND2XL U111 ( .A(n103), .B(n253), .Y(n305) );
  AOI22XL U112 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI2BB2XL U113 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  NOR2XL U114 ( .A(n293), .B(n292), .Y(n294) );
  AOI22XL U115 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  NAND2XL U116 ( .A(n352), .B(n351), .Y(n358) );
  OAI22XL U117 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI22XL U118 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  AOI22XL U119 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  AOI2BB2XL U120 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U121 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  INVXL U122 ( .A(n82), .Y(n172) );
  AOI22XL U123 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI22XL U124 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  NOR2XL U125 ( .A(n161), .B(n309), .Y(n162) );
  AOI22XL U126 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  AOI32XL U127 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  AOI211XL U128 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  AOI22XL U129 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  INVXL U130 ( .A(n180), .Y(n183) );
  AOI211XL U131 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  INVXL U132 ( .A(n312), .Y(n313) );
  AOI22XL U133 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  OAI22XL U134 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  AOI22XL U135 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  NAND3XL U136 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  OAI2BB1XL U137 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  AOI22XL U138 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  AOI22XL U139 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  NAND2XL U140 ( .A(n350), .B(n245), .Y(n180) );
  OAI22XL U141 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U142 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AOI22XL U143 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  NOR2XL U144 ( .A(n268), .B(n354), .Y(n13) );
  AND2X2 U145 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U146 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  AOI22XL U147 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  AOI22XL U148 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  AOI22XL U149 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  NOR3XL U150 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  AOI31XL U151 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI22XL U152 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  NOR2XL U153 ( .A(n37), .B(n145), .Y(n99) );
  AOI22XL U154 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  AOI211XL U155 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  OAI22XL U156 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI22XL U157 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  AOI22XL U158 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  AOI22XL U159 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  AOI22XL U160 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  NAND2XL U161 ( .A(n311), .B(n196), .Y(n40) );
  NOR2XL U162 ( .A(n293), .B(n226), .Y(n39) );
  AOI2BB2XL U163 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  NOR2XL U164 ( .A(n181), .B(n269), .Y(n315) );
  NAND2XL U165 ( .A(n311), .B(n236), .Y(n346) );
  AOI22XL U166 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  INVXL U167 ( .A(n131), .Y(n351) );
  NOR3XL U168 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI22XL U169 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NAND3XL U170 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NAND3XL U171 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  NOR2XL U172 ( .A(n37), .B(a[1]), .Y(n195) );
  NAND2XL U173 ( .A(n306), .B(n267), .Y(n61) );
  AOI22XL U174 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NOR2XL U175 ( .A(a[1]), .B(n249), .Y(n131) );
  NAND2XL U176 ( .A(n329), .B(n323), .Y(n245) );
  AOI22XL U177 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  NAND2XL U178 ( .A(n311), .B(n303), .Y(n38) );
  NOR2XL U179 ( .A(a[1]), .B(n329), .Y(n269) );
  AOI22XL U180 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  NOR2XL U181 ( .A(n233), .B(n331), .Y(n108) );
  NOR2XL U182 ( .A(n187), .B(n186), .Y(n290) );
  AOI22XL U183 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  AOI22XL U184 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  NAND2XL U185 ( .A(n107), .B(n348), .Y(n175) );
  NAND3XL U186 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  INVXL U187 ( .A(n197), .Y(n185) );
  NAND2XL U188 ( .A(n328), .B(n311), .Y(n353) );
  NAND2XL U189 ( .A(a[1]), .B(n261), .Y(n303) );
  INVXL U190 ( .A(n332), .Y(n234) );
  INVXL U191 ( .A(n297), .Y(n284) );
  NOR2XL U192 ( .A(n264), .B(n273), .Y(n330) );
  NAND2XL U193 ( .A(n264), .B(n275), .Y(n252) );
  INVXL U194 ( .A(n274), .Y(n251) );
  AOI22XL U195 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  NOR2XL U196 ( .A(a[1]), .B(n198), .Y(n160) );
  AOI22XL U197 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U198 ( .A(a[3]), .B(a[1]), .Y(n225) );
  INVX2 U199 ( .A(a[7]), .Y(n264) );
  NAND2XL U200 ( .A(a[4]), .B(a[1]), .Y(n274) );
  NAND2XL U201 ( .A(a[3]), .B(a[1]), .Y(n20) );
  CLKINVX3 U202 ( .A(n266), .Y(n329) );
  NAND2X2 U203 ( .A(a[4]), .B(n31), .Y(n266) );
  OAI21X1 U204 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U205 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U206 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U207 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U208 ( .A(a[5]), .Y(n275) );
  NOR2X2 U209 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U210 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U211 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U212 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U213 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U214 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U215 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U216 ( .A(n233), .Y(n359) );
  NAND2X2 U217 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U218 ( .A(n349), .Y(n288) );
  NOR2X4 U219 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U220 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U221 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U222 ( .A(n347), .Y(n1) );
  CLKINVX3 U223 ( .A(a[2]), .Y(n273) );
  OAI21X1 U224 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U225 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U226 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U227 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U228 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U229 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31X4 U230 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  CLKINVX3 U231 ( .A(n309), .Y(n345) );
  NAND2X2 U232 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U233 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U234 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U235 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U236 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U237 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U238 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U239 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U240 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U241 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U242 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U243 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U244 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U245 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U246 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U247 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U248 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U249 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U250 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U251 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U252 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U253 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U254 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U255 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U256 ( .A(a[1]), .Y(n323) );
  NAND2X1 U257 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U258 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U259 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U260 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U261 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U262 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U263 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U264 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U265 ( .A(n242), .Y(n249) );
  OAI21XL U266 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U267 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U268 ( .A(n192), .Y(n205) );
  INVX1 U269 ( .A(n66), .Y(n111) );
  NOR2X1 U270 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U271 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U272 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U273 ( .A(a[6]), .B(a[0]), .Y(n360) );
  INVX1 U274 ( .A(a[6]), .Y(n16) );
  NOR2X1 U275 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U276 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U277 ( .A(n261), .Y(n307) );
  INVX1 U278 ( .A(n20), .Y(n326) );
  NAND2X1 U279 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U280 ( .A(n187), .Y(n196) );
  INVX1 U281 ( .A(n350), .Y(n335) );
  NAND2X1 U282 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U283 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U284 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U285 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U286 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U287 ( .A(n103), .Y(n37) );
  NOR2X1 U288 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U289 ( .A(n311), .Y(n268) );
  INVX1 U290 ( .A(n293), .Y(n209) );
  NOR2X1 U291 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U292 ( .A(n224), .Y(n235) );
  NAND2X1 U293 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U294 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U295 ( .A(n195), .Y(n142) );
  NAND2X1 U296 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U297 ( .A(n226), .Y(n253) );
  NAND2X1 U298 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U299 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U300 ( .A(n1), .Y(n301) );
  NAND2X1 U301 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U302 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U303 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U304 ( .A(n89), .Y(n340) );
  AOI211X1 U305 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U306 ( .A(n327), .Y(n248) );
  INVX1 U307 ( .A(n181), .Y(n109) );
  INVX1 U308 ( .A(n225), .Y(n302) );
  NAND2X1 U309 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U310 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U311 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U312 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U313 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U314 ( .A(n270), .Y(n107) );
  INVX1 U315 ( .A(n306), .Y(n145) );
  NAND4X1 U316 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U317 ( .A(n210), .Y(n236) );
  INVX1 U318 ( .A(n331), .Y(n78) );
  INVX1 U319 ( .A(n328), .Y(n314) );
  OAI21XL U320 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U321 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U322 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U323 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  NOR2X1 U324 ( .A(n181), .B(n95), .Y(n174) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_15 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  NAND2X1 U4 ( .A(n194), .B(n274), .Y(n344) );
  INVX1 U5 ( .A(n324), .Y(n265) );
  AOI21XL U6 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  AOI211XL U7 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  INVXL U8 ( .A(n257), .Y(n289) );
  OAI211XL U9 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  NAND2XL U10 ( .A(n235), .B(n265), .Y(n338) );
  INVXL U11 ( .A(n116), .Y(n203) );
  NOR2XL U12 ( .A(n224), .B(n326), .Y(n257) );
  AOI22XL U13 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NAND2XL U14 ( .A(n109), .B(n78), .Y(n158) );
  NOR2XL U15 ( .A(n248), .B(n142), .Y(n357) );
  NOR2X1 U16 ( .A(a[1]), .B(n293), .Y(n318) );
  NOR2X1 U17 ( .A(n293), .B(n323), .Y(n150) );
  NAND2XL U18 ( .A(a[1]), .B(n293), .Y(n82) );
  NOR2XL U19 ( .A(n324), .B(n131), .Y(n262) );
  NOR2X4 U20 ( .A(n264), .B(n197), .Y(n350) );
  NOR2X1 U21 ( .A(a[1]), .B(n103), .Y(n331) );
  INVXL U22 ( .A(n352), .Y(n141) );
  NOR2XL U23 ( .A(a[1]), .B(n242), .Y(n186) );
  INVXL U24 ( .A(n267), .Y(n333) );
  NAND2X1 U25 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI211XL U26 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U27 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI211XL U28 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  OR4X2 U29 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI31XL U30 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI211XL U31 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U32 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI31XL U33 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI31XL U34 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U35 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  OAI211XL U36 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U37 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI31XL U38 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  OAI211XL U39 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI22XL U40 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  OAI22XL U41 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI211XL U42 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI31XL U43 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI31XL U44 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI211XL U45 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI211XL U46 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U47 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI31XL U48 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  AOI21X1 U49 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  OAI211XL U50 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI31XL U51 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U52 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI22XL U53 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI211XL U54 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI22XL U55 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  AOI211XL U56 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  INVXL U57 ( .A(n101), .Y(n254) );
  NAND2XL U58 ( .A(n296), .B(n101), .Y(n94) );
  AOI31XL U59 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  AOI31XL U60 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  AOI2BB2XL U61 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI211XL U62 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  AOI22XL U63 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U64 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U65 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  OAI211XL U66 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U67 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI31XL U68 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI22XL U69 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  NAND2XL U70 ( .A(n235), .B(n274), .Y(n184) );
  AOI221XL U71 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI22XL U72 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  NOR2XL U73 ( .A(n150), .B(n331), .Y(n130) );
  AOI211XL U74 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI211XL U75 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI31XL U76 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  AOI31XL U77 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI211XL U78 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  OAI211XL U79 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  INVXL U80 ( .A(n150), .Y(n310) );
  AOI22XL U81 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  NOR2XL U82 ( .A(n224), .B(n150), .Y(n116) );
  AOI22XL U83 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI22XL U84 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI22XL U85 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI22XL U86 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI2BB2XL U87 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U88 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI31XL U89 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI211XL U90 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI22XL U91 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI2BB2XL U92 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI22XL U93 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  NAND2XL U94 ( .A(n265), .B(n348), .Y(n247) );
  AOI211XL U95 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI211XL U96 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI211XL U97 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI211XL U98 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  INVXL U99 ( .A(n152), .Y(n222) );
  OAI22XL U100 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI2BB2XL U101 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI22XL U102 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI22XL U103 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI211XL U104 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI22XL U105 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  OAI211XL U106 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U107 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  NAND2XL U108 ( .A(n103), .B(n253), .Y(n305) );
  AOI22XL U109 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  NAND2XL U110 ( .A(n352), .B(n351), .Y(n358) );
  AOI22XL U111 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  INVXL U112 ( .A(n312), .Y(n313) );
  NOR2XL U113 ( .A(n293), .B(n292), .Y(n294) );
  NOR2XL U114 ( .A(n209), .B(n233), .Y(n256) );
  AOI22XL U115 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  NAND3XL U116 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  AOI22XL U117 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  AOI22XL U118 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI2BB2XL U119 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  OAI22XL U120 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  INVXL U121 ( .A(n82), .Y(n172) );
  AOI2BB2XL U122 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U123 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI22XL U124 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  NOR2XL U125 ( .A(n161), .B(n309), .Y(n162) );
  AOI22XL U126 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  AOI22XL U127 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  AOI211XL U128 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  OAI2BB1XL U129 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  AOI22XL U130 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  NAND2XL U131 ( .A(n109), .B(n242), .Y(n135) );
  AOI22XL U132 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  AOI32XL U133 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  OAI22XL U134 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  INVXL U135 ( .A(n180), .Y(n183) );
  AOI211XL U136 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  AOI31XL U137 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI22XL U138 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  NOR2XL U139 ( .A(n37), .B(n145), .Y(n99) );
  NOR3XL U140 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI22XL U141 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  AOI2BB2XL U142 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  INVXL U143 ( .A(n131), .Y(n351) );
  AOI211XL U144 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  NOR2XL U145 ( .A(n181), .B(n269), .Y(n315) );
  AOI22XL U146 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  AND2X2 U147 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U148 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  OAI22XL U149 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI22XL U150 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  AOI22XL U151 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  AOI22XL U152 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  NAND2XL U153 ( .A(n350), .B(n245), .Y(n180) );
  AOI22XL U154 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  NOR3XL U155 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  AOI22XL U156 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  AOI22XL U157 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  AOI22XL U158 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  NAND2XL U159 ( .A(n311), .B(n236), .Y(n346) );
  AOI22XL U160 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  NAND2XL U161 ( .A(n311), .B(n196), .Y(n40) );
  NOR2XL U162 ( .A(n293), .B(n226), .Y(n39) );
  AOI22XL U163 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  OAI22XL U164 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U165 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  NOR2XL U166 ( .A(n268), .B(n354), .Y(n13) );
  AOI22XL U167 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AOI22XL U168 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  NAND2XL U169 ( .A(n329), .B(n323), .Y(n245) );
  NOR2XL U170 ( .A(n187), .B(n186), .Y(n290) );
  AOI22XL U171 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  NOR2XL U172 ( .A(n233), .B(n331), .Y(n108) );
  NAND3XL U173 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  AOI22XL U174 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  AOI22XL U175 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  AOI22XL U176 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NAND2XL U177 ( .A(n306), .B(n267), .Y(n61) );
  AOI22XL U178 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  NAND2XL U179 ( .A(n311), .B(n303), .Y(n38) );
  NAND3XL U180 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NOR2XL U181 ( .A(a[1]), .B(n249), .Y(n131) );
  NOR2XL U182 ( .A(n37), .B(a[1]), .Y(n195) );
  NAND2XL U183 ( .A(n107), .B(n348), .Y(n175) );
  NOR2XL U184 ( .A(a[1]), .B(n329), .Y(n269) );
  NAND3XL U185 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  INVXL U186 ( .A(n332), .Y(n234) );
  INVXL U187 ( .A(n197), .Y(n185) );
  INVXL U188 ( .A(n297), .Y(n284) );
  NAND2XL U189 ( .A(n328), .B(n311), .Y(n353) );
  NAND2XL U190 ( .A(a[1]), .B(n261), .Y(n303) );
  NOR2XL U191 ( .A(a[1]), .B(n198), .Y(n160) );
  AOI22XL U192 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  INVXL U193 ( .A(n274), .Y(n251) );
  NOR2XL U194 ( .A(n264), .B(n273), .Y(n330) );
  NAND2XL U195 ( .A(n264), .B(n275), .Y(n252) );
  AOI22XL U196 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  INVX2 U197 ( .A(a[7]), .Y(n264) );
  NOR2XL U198 ( .A(a[3]), .B(a[1]), .Y(n225) );
  NAND2XL U199 ( .A(a[4]), .B(a[1]), .Y(n274) );
  INVX1 U200 ( .A(a[6]), .Y(n16) );
  NAND2XL U201 ( .A(a[3]), .B(a[1]), .Y(n20) );
  CLKINVX3 U202 ( .A(n266), .Y(n329) );
  NAND2X2 U203 ( .A(a[4]), .B(n31), .Y(n266) );
  OAI21X1 U204 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U205 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U206 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U207 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U208 ( .A(a[5]), .Y(n275) );
  NOR2X2 U209 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U210 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U211 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U212 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U213 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U214 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U215 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U216 ( .A(n233), .Y(n359) );
  NAND2X2 U217 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U218 ( .A(n349), .Y(n288) );
  NOR2X4 U219 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U220 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U221 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U222 ( .A(n347), .Y(n1) );
  CLKINVX3 U223 ( .A(a[2]), .Y(n273) );
  OAI21X1 U224 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U225 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U226 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U227 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U228 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U229 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31X4 U230 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  CLKINVX3 U231 ( .A(n309), .Y(n345) );
  NAND2X2 U232 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U233 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U234 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U235 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U236 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U237 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U238 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U239 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U240 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U241 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U242 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U243 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U244 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U245 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U246 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U247 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U248 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U249 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U250 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U251 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U252 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U253 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U254 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U255 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U256 ( .A(a[1]), .Y(n323) );
  NAND2X1 U257 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U258 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U259 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U260 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U261 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U262 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U263 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U264 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U265 ( .A(n242), .Y(n249) );
  OAI21XL U266 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U267 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U268 ( .A(n192), .Y(n205) );
  INVX1 U269 ( .A(n66), .Y(n111) );
  NOR2X1 U270 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U271 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U272 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U273 ( .A(a[6]), .B(a[0]), .Y(n360) );
  NOR2X1 U274 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U275 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U276 ( .A(n261), .Y(n307) );
  INVX1 U277 ( .A(n20), .Y(n326) );
  NAND2X1 U278 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U279 ( .A(n187), .Y(n196) );
  INVX1 U280 ( .A(n350), .Y(n335) );
  NAND2X1 U281 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U282 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U283 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U284 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U285 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U286 ( .A(n103), .Y(n37) );
  NOR2X1 U287 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U288 ( .A(n311), .Y(n268) );
  INVX1 U289 ( .A(n293), .Y(n209) );
  NOR2X1 U290 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U291 ( .A(n224), .Y(n235) );
  NAND2X1 U292 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U293 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U294 ( .A(n195), .Y(n142) );
  NAND2X1 U295 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U296 ( .A(n226), .Y(n253) );
  NAND2X1 U297 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U298 ( .A(n140), .B(n20), .Y(n151) );
  NAND2X1 U299 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U300 ( .A(n1), .Y(n301) );
  NAND2X1 U301 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U302 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U303 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U304 ( .A(n89), .Y(n340) );
  AOI211X1 U305 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U306 ( .A(n327), .Y(n248) );
  INVX1 U307 ( .A(n181), .Y(n109) );
  INVX1 U308 ( .A(n225), .Y(n302) );
  NAND2X1 U309 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U310 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U311 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U312 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U313 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U314 ( .A(n270), .Y(n107) );
  INVX1 U315 ( .A(n306), .Y(n145) );
  NAND4X1 U316 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U317 ( .A(n210), .Y(n236) );
  INVX1 U318 ( .A(n331), .Y(n78) );
  INVX1 U319 ( .A(n328), .Y(n314) );
  OAI21XL U320 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U321 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U322 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U323 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  NOR2X1 U324 ( .A(n181), .B(n95), .Y(n174) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U334 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U335 ( .A(n125), .Y(n319) );
  NAND2X1 U336 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U337 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U338 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U339 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U340 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U341 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U342 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U343 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U344 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U345 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U346 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U347 ( .A(n117), .Y(n188) );
  OAI21XL U348 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U349 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U350 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_16 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  AOI21XL U4 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  AOI211XL U5 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  INVX1 U6 ( .A(n116), .Y(n203) );
  NAND2X1 U7 ( .A(n140), .B(n20), .Y(n151) );
  INVX1 U8 ( .A(n324), .Y(n265) );
  AOI2BB2XL U9 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI21XL U10 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  NAND2XL U11 ( .A(n235), .B(n265), .Y(n338) );
  INVXL U12 ( .A(n257), .Y(n289) );
  NOR2XL U13 ( .A(n224), .B(n326), .Y(n257) );
  NAND2XL U14 ( .A(n109), .B(n78), .Y(n158) );
  AOI22XL U15 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NOR2XL U16 ( .A(n324), .B(n131), .Y(n262) );
  NAND2XL U17 ( .A(n194), .B(n274), .Y(n344) );
  NOR2X1 U18 ( .A(a[1]), .B(n293), .Y(n318) );
  NOR2X1 U19 ( .A(n293), .B(n323), .Y(n150) );
  NOR2XL U20 ( .A(n181), .B(n95), .Y(n174) );
  NAND2XL U21 ( .A(a[1]), .B(n293), .Y(n82) );
  NOR2XL U22 ( .A(a[1]), .B(n242), .Y(n186) );
  INVXL U23 ( .A(n352), .Y(n141) );
  NOR2X4 U24 ( .A(n264), .B(n197), .Y(n350) );
  NOR2X1 U25 ( .A(a[1]), .B(n103), .Y(n331) );
  INVXL U26 ( .A(n267), .Y(n333) );
  NAND2X1 U27 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI211XL U28 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U29 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI211XL U30 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  OR4X2 U31 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI31XL U32 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI31XL U33 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U34 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI31XL U35 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  AOI31XL U36 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI31XL U37 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  OAI211XL U38 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI211XL U39 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U40 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI22XL U41 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI31XL U42 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI31XL U43 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI22XL U44 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  OAI211XL U45 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI22XL U46 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  OAI22XL U47 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  OAI211XL U48 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI211XL U49 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI211XL U50 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI211XL U51 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI31XL U52 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  AOI211XL U53 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI211XL U54 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI31XL U55 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U56 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  INVXL U57 ( .A(n101), .Y(n254) );
  NAND2XL U58 ( .A(n296), .B(n101), .Y(n94) );
  AOI31XL U59 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  OAI211XL U60 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  OAI211XL U61 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U62 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI22XL U63 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U64 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U65 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U66 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  AOI211XL U67 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  AOI31XL U68 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  INVXL U69 ( .A(n150), .Y(n310) );
  AOI211XL U70 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  AOI31XL U71 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI221XL U72 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI211XL U73 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI22XL U74 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  NOR2XL U75 ( .A(n224), .B(n150), .Y(n116) );
  AOI22XL U76 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  AOI31XL U77 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  NAND2XL U78 ( .A(n235), .B(n274), .Y(n184) );
  NOR2XL U79 ( .A(n150), .B(n331), .Y(n130) );
  AOI211XL U80 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI31XL U81 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI22XL U82 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  OAI211XL U83 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  AOI211XL U84 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI22XL U85 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI2BB2XL U86 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  NAND2XL U87 ( .A(n265), .B(n348), .Y(n247) );
  AOI2BB2XL U88 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U89 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI22XL U90 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  INVXL U91 ( .A(n152), .Y(n222) );
  AOI22XL U92 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI22XL U93 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI211XL U94 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI22XL U95 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI22XL U96 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  OAI22XL U97 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI211XL U98 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI22XL U99 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI22XL U100 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI2BB2XL U101 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI211XL U102 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI211XL U103 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI31XL U104 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI22XL U105 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI211XL U106 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  AOI211XL U107 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  INVXL U108 ( .A(n180), .Y(n183) );
  OAI2BB1XL U109 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  OAI22XL U110 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI22XL U111 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  INVXL U112 ( .A(n82), .Y(n172) );
  AOI22XL U113 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  INVXL U114 ( .A(n312), .Y(n313) );
  OAI211XL U115 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U116 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  NAND2XL U117 ( .A(n352), .B(n351), .Y(n358) );
  NOR2XL U118 ( .A(n293), .B(n292), .Y(n294) );
  AOI2BB2XL U119 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  AOI22XL U120 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI22XL U121 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  AOI22XL U122 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  NOR2XL U123 ( .A(n161), .B(n309), .Y(n162) );
  NAND2XL U124 ( .A(n103), .B(n253), .Y(n305) );
  AOI22XL U125 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  AOI22XL U126 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI22XL U127 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI22XL U128 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  OAI22XL U129 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  AOI22XL U130 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  NOR2XL U131 ( .A(n209), .B(n233), .Y(n256) );
  NAND3XL U132 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  AOI32XL U133 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  NAND2XL U134 ( .A(n109), .B(n242), .Y(n135) );
  AOI211XL U135 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI2BB2XL U136 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U137 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  NOR2XL U138 ( .A(n37), .B(n145), .Y(n99) );
  AND2X2 U139 ( .A(n303), .B(n78), .Y(n221) );
  INVXL U140 ( .A(n131), .Y(n351) );
  NOR2XL U141 ( .A(n293), .B(n226), .Y(n39) );
  AOI31XL U142 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  NOR3XL U143 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI211XL U144 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  AOI22XL U145 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  AOI22XL U146 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  NOR2XL U147 ( .A(n181), .B(n269), .Y(n315) );
  AOI22XL U148 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  NOR2XL U149 ( .A(n268), .B(n354), .Y(n13) );
  AOI22XL U150 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  AOI22XL U151 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI2BB2XL U152 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U153 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  NAND2XL U154 ( .A(n311), .B(n196), .Y(n40) );
  AOI22XL U155 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  AOI22XL U156 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  NAND2XL U157 ( .A(n350), .B(n245), .Y(n180) );
  OAI22XL U158 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U159 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AOI22XL U160 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AOI22XL U161 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  AOI22XL U162 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  OAI22XL U163 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI22XL U164 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  NOR3XL U165 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  AOI22XL U166 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  NAND2XL U167 ( .A(n311), .B(n236), .Y(n346) );
  AOI22XL U168 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  NAND2XL U169 ( .A(n107), .B(n348), .Y(n175) );
  AOI22XL U170 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  AOI22XL U171 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  NOR2XL U172 ( .A(a[1]), .B(n329), .Y(n269) );
  NAND2XL U173 ( .A(n329), .B(n323), .Y(n245) );
  NOR2XL U174 ( .A(n187), .B(n186), .Y(n290) );
  NAND3XL U175 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  NAND3XL U176 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NOR2XL U177 ( .A(n233), .B(n331), .Y(n108) );
  NOR2XL U178 ( .A(n37), .B(a[1]), .Y(n195) );
  NOR2XL U179 ( .A(a[1]), .B(n249), .Y(n131) );
  NAND2XL U180 ( .A(n311), .B(n303), .Y(n38) );
  AOI22XL U181 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  AOI22XL U182 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  AOI22XL U183 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  AOI22XL U184 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  NAND2XL U185 ( .A(n306), .B(n267), .Y(n61) );
  INVXL U186 ( .A(n197), .Y(n185) );
  INVXL U187 ( .A(n332), .Y(n234) );
  NAND3XL U188 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  NAND2XL U189 ( .A(n328), .B(n311), .Y(n353) );
  INVXL U190 ( .A(n297), .Y(n284) );
  NAND2XL U191 ( .A(a[1]), .B(n261), .Y(n303) );
  AOI22XL U192 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  NOR2XL U193 ( .A(a[1]), .B(n198), .Y(n160) );
  NAND2XL U194 ( .A(n264), .B(n275), .Y(n252) );
  AOI22XL U195 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U196 ( .A(n264), .B(n273), .Y(n330) );
  INVXL U197 ( .A(n274), .Y(n251) );
  NAND2XL U198 ( .A(a[3]), .B(a[1]), .Y(n20) );
  NAND2XL U199 ( .A(a[4]), .B(a[1]), .Y(n274) );
  INVX2 U200 ( .A(a[7]), .Y(n264) );
  NOR2XL U201 ( .A(a[3]), .B(a[1]), .Y(n225) );
  CLKINVX3 U202 ( .A(n266), .Y(n329) );
  NAND2X2 U203 ( .A(a[4]), .B(n31), .Y(n266) );
  OAI21X1 U204 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U205 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U206 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U207 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U208 ( .A(a[5]), .Y(n275) );
  NOR2X2 U209 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U210 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U211 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U212 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U213 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U214 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U215 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U216 ( .A(n233), .Y(n359) );
  NAND2X2 U217 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U218 ( .A(n349), .Y(n288) );
  NOR2X4 U219 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U220 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U221 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U222 ( .A(n347), .Y(n1) );
  CLKINVX3 U223 ( .A(a[2]), .Y(n273) );
  OAI21X1 U224 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U225 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U226 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U227 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U228 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U229 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31X4 U230 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  CLKINVX3 U231 ( .A(n309), .Y(n345) );
  NAND2X2 U232 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U233 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U234 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U235 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U236 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U237 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U238 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U239 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U240 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U241 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U242 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U243 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U244 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U245 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U246 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U247 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U248 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U249 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U250 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U251 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U252 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U253 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U254 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U255 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U256 ( .A(a[1]), .Y(n323) );
  NAND2X1 U257 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U258 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U259 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U260 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U261 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U262 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U263 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U264 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U265 ( .A(n242), .Y(n249) );
  OAI21XL U266 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U267 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U268 ( .A(n192), .Y(n205) );
  INVX1 U269 ( .A(n66), .Y(n111) );
  NOR2X1 U270 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U271 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U272 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U273 ( .A(a[6]), .B(a[0]), .Y(n360) );
  INVX1 U274 ( .A(a[6]), .Y(n16) );
  NOR2X1 U275 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U276 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U277 ( .A(n261), .Y(n307) );
  INVX1 U278 ( .A(n20), .Y(n326) );
  NAND2X1 U279 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U280 ( .A(n187), .Y(n196) );
  INVX1 U281 ( .A(n350), .Y(n335) );
  NAND2X1 U282 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U283 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U284 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U285 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U286 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U287 ( .A(n103), .Y(n37) );
  NOR2X1 U288 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U289 ( .A(n311), .Y(n268) );
  INVX1 U290 ( .A(n293), .Y(n209) );
  NOR2X1 U291 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U292 ( .A(n224), .Y(n235) );
  NAND2X1 U293 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U294 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U295 ( .A(n195), .Y(n142) );
  NAND2X1 U296 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U297 ( .A(n226), .Y(n253) );
  NAND2X1 U298 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U299 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U300 ( .A(n1), .Y(n301) );
  NAND2X1 U301 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U302 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U303 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U304 ( .A(n89), .Y(n340) );
  AOI211X1 U305 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U306 ( .A(n327), .Y(n248) );
  INVX1 U307 ( .A(n181), .Y(n109) );
  INVX1 U308 ( .A(n225), .Y(n302) );
  NAND2X1 U309 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U310 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U311 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U312 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U313 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U314 ( .A(n270), .Y(n107) );
  INVX1 U315 ( .A(n306), .Y(n145) );
  NAND4X1 U316 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U317 ( .A(n210), .Y(n236) );
  INVX1 U318 ( .A(n331), .Y(n78) );
  INVX1 U319 ( .A(n328), .Y(n314) );
  OAI21XL U320 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U321 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U322 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U323 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U324 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U325 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U326 ( .A(n186), .Y(n194) );
  NAND2X1 U327 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U328 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U329 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U330 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U331 ( .A(n72), .Y(n204) );
  OAI21XL U332 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U333 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U334 ( .A(n125), .Y(n319) );
  NAND2X1 U335 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U336 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U337 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U338 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U339 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U340 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U341 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U342 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U343 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U344 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U345 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U346 ( .A(n117), .Y(n188) );
  OAI21XL U347 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U348 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U349 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  NOR2X1 U350 ( .A(n248), .B(n142), .Y(n357) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_17 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  AOI211XL U4 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  AOI21XL U5 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  INVX1 U6 ( .A(n116), .Y(n203) );
  NAND2XL U7 ( .A(n235), .B(n265), .Y(n338) );
  NAND2XL U8 ( .A(n345), .B(n209), .Y(n93) );
  NAND2X1 U9 ( .A(n194), .B(n274), .Y(n344) );
  INVX1 U10 ( .A(n324), .Y(n265) );
  AOI31XL U11 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  AOI21XL U12 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  AOI2BB2XL U13 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  INVXL U14 ( .A(n257), .Y(n289) );
  NOR2XL U15 ( .A(n224), .B(n326), .Y(n257) );
  AOI22XL U16 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NAND2XL U17 ( .A(n109), .B(n78), .Y(n158) );
  NOR2XL U18 ( .A(n181), .B(n95), .Y(n174) );
  NOR2X1 U19 ( .A(n293), .B(n323), .Y(n150) );
  NOR2X1 U20 ( .A(a[1]), .B(n293), .Y(n318) );
  NAND2XL U21 ( .A(n140), .B(n20), .Y(n151) );
  NAND2XL U22 ( .A(a[1]), .B(n293), .Y(n82) );
  NOR2XL U23 ( .A(n324), .B(n131), .Y(n262) );
  INVXL U24 ( .A(n352), .Y(n141) );
  NOR2X4 U25 ( .A(n264), .B(n197), .Y(n350) );
  NOR2XL U26 ( .A(a[1]), .B(n242), .Y(n186) );
  INVXL U27 ( .A(n267), .Y(n333) );
  NOR2X1 U28 ( .A(a[1]), .B(n103), .Y(n331) );
  NAND2X1 U29 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI211XL U30 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI211XL U31 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  AOI31XL U32 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  OR4X2 U33 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U34 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U35 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  OAI211XL U36 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U37 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI31XL U38 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U39 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI31XL U40 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U41 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI31XL U42 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  OAI22XL U43 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI31XL U44 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI211XL U45 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI211XL U46 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  OAI211XL U47 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI211XL U48 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U49 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI211XL U50 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI22XL U51 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI22XL U52 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI31XL U53 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  AOI211XL U54 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI31XL U55 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  OAI211XL U56 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI22XL U57 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  NAND2XL U58 ( .A(n296), .B(n101), .Y(n94) );
  AOI22XL U59 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI211XL U60 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  OAI211XL U61 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  INVXL U62 ( .A(n101), .Y(n254) );
  AOI31XL U63 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  AOI31XL U64 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  AOI211XL U65 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  OAI211XL U66 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI211XL U67 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U68 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U69 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  AOI211XL U70 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  AOI31XL U71 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  AOI22XL U72 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  OAI211XL U73 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  AOI211XL U74 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI221XL U75 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI22XL U76 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI211XL U77 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  NAND2XL U78 ( .A(n235), .B(n274), .Y(n184) );
  AOI31XL U79 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  AOI22XL U80 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  NOR2XL U81 ( .A(n150), .B(n331), .Y(n130) );
  AOI31XL U82 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  INVXL U83 ( .A(n150), .Y(n310) );
  NOR2XL U84 ( .A(n224), .B(n150), .Y(n116) );
  NAND2XL U85 ( .A(n265), .B(n348), .Y(n247) );
  AOI22XL U86 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  AOI22XL U87 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI22XL U88 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  INVXL U89 ( .A(n152), .Y(n222) );
  AOI211XL U90 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI22XL U91 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI22XL U92 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI2BB2XL U93 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI22XL U94 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI22XL U95 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI211XL U96 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI211XL U97 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI31XL U98 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI2BB2XL U99 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  AOI22XL U100 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI211XL U101 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI22XL U102 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  AOI211XL U103 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI22XL U104 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI211XL U105 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  OAI22XL U106 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI2BB2XL U107 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  OAI22XL U108 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI211XL U109 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  AOI22XL U110 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  AOI22XL U111 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  AOI22XL U112 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  AOI2BB2XL U113 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U114 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  AOI22XL U115 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  OAI22XL U116 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  NAND3XL U117 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  OAI2BB1XL U118 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  NOR2XL U119 ( .A(n209), .B(n233), .Y(n256) );
  INVXL U120 ( .A(n312), .Y(n313) );
  AOI2BB2XL U121 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  AOI22XL U122 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  NOR2XL U123 ( .A(n293), .B(n292), .Y(n294) );
  OAI211XL U124 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  NOR2XL U125 ( .A(n161), .B(n309), .Y(n162) );
  NAND2XL U126 ( .A(n352), .B(n351), .Y(n358) );
  AOI22XL U127 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  NAND2XL U128 ( .A(n103), .B(n253), .Y(n305) );
  NAND2XL U129 ( .A(n109), .B(n242), .Y(n135) );
  AOI22XL U130 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  AOI22XL U131 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  AOI22XL U132 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  AOI32XL U133 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  INVXL U134 ( .A(n180), .Y(n183) );
  AOI211XL U135 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  AOI22XL U136 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  AOI22XL U137 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  INVXL U138 ( .A(n82), .Y(n172) );
  AOI22XL U139 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  AOI22XL U140 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  NAND2XL U141 ( .A(n311), .B(n236), .Y(n346) );
  INVXL U142 ( .A(n131), .Y(n351) );
  AOI22XL U143 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  AOI22XL U144 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  AOI22XL U145 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  AOI22XL U146 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  NOR2XL U147 ( .A(n293), .B(n226), .Y(n39) );
  AOI2BB2XL U148 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U149 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  NOR2XL U150 ( .A(n181), .B(n269), .Y(n315) );
  NOR2XL U151 ( .A(n268), .B(n354), .Y(n13) );
  NOR3XL U152 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  AOI22XL U153 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  AOI22XL U154 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AND2X2 U155 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U156 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  AOI22XL U157 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  OAI22XL U158 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  NAND2XL U159 ( .A(n350), .B(n245), .Y(n180) );
  AOI22XL U160 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  AOI22XL U161 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  NOR2XL U162 ( .A(n37), .B(n145), .Y(n99) );
  NAND2XL U163 ( .A(n311), .B(n196), .Y(n40) );
  AOI22XL U164 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  NOR3XL U165 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  AOI211XL U166 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  AOI31XL U167 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  OAI22XL U168 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  AOI22XL U169 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  AOI22XL U170 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  NAND2XL U171 ( .A(n329), .B(n323), .Y(n245) );
  NAND2XL U172 ( .A(n107), .B(n348), .Y(n175) );
  AOI22XL U173 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  AOI22XL U174 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NAND2XL U175 ( .A(n306), .B(n267), .Y(n61) );
  NOR2XL U176 ( .A(n233), .B(n331), .Y(n108) );
  AOI22XL U177 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  AOI22XL U178 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  NAND3XL U179 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NOR2XL U180 ( .A(n37), .B(a[1]), .Y(n195) );
  NOR2XL U181 ( .A(n187), .B(n186), .Y(n290) );
  NAND3XL U182 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  AOI22XL U183 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  NAND2XL U184 ( .A(n311), .B(n303), .Y(n38) );
  NOR2XL U185 ( .A(a[1]), .B(n329), .Y(n269) );
  NOR2XL U186 ( .A(a[1]), .B(n249), .Y(n131) );
  NAND3XL U187 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  NAND2XL U188 ( .A(n328), .B(n311), .Y(n353) );
  INVXL U189 ( .A(n332), .Y(n234) );
  NAND2XL U190 ( .A(a[1]), .B(n261), .Y(n303) );
  INVXL U191 ( .A(n197), .Y(n185) );
  INVXL U192 ( .A(n297), .Y(n284) );
  INVXL U193 ( .A(n274), .Y(n251) );
  AOI22XL U194 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  AOI22XL U195 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U196 ( .A(n264), .B(n273), .Y(n330) );
  NOR2XL U197 ( .A(a[1]), .B(n198), .Y(n160) );
  NAND2XL U198 ( .A(n264), .B(n275), .Y(n252) );
  NAND2XL U199 ( .A(a[4]), .B(a[1]), .Y(n274) );
  NAND2XL U200 ( .A(a[3]), .B(a[1]), .Y(n20) );
  INVX2 U201 ( .A(a[7]), .Y(n264) );
  NOR2XL U202 ( .A(a[3]), .B(a[1]), .Y(n225) );
  CLKINVX3 U203 ( .A(n266), .Y(n329) );
  NAND2X2 U204 ( .A(a[4]), .B(n31), .Y(n266) );
  OAI21X1 U205 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U206 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U207 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U208 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U209 ( .A(a[5]), .Y(n275) );
  NOR2X2 U210 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U211 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U212 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U213 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U214 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U215 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U216 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U217 ( .A(n233), .Y(n359) );
  NAND2X2 U218 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U219 ( .A(n349), .Y(n288) );
  NOR2X4 U220 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U221 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U222 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U223 ( .A(n347), .Y(n1) );
  CLKINVX3 U224 ( .A(a[2]), .Y(n273) );
  OAI21X1 U225 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U226 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U227 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U228 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U229 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U230 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31X4 U231 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  CLKINVX3 U232 ( .A(n309), .Y(n345) );
  NAND2X2 U233 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U234 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U235 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U236 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U237 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U238 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U239 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U240 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U241 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U242 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U243 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U244 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U245 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U246 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U247 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U248 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U249 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U250 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U251 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U252 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U253 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U254 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U255 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U256 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U257 ( .A(a[1]), .Y(n323) );
  NAND2X1 U258 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U259 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U260 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U261 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U262 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U263 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U264 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U265 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U266 ( .A(n242), .Y(n249) );
  OAI21XL U267 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U268 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U269 ( .A(n192), .Y(n205) );
  INVX1 U270 ( .A(n66), .Y(n111) );
  NOR2X1 U271 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U272 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U273 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U274 ( .A(a[6]), .B(a[0]), .Y(n360) );
  INVX1 U275 ( .A(a[6]), .Y(n16) );
  NOR2X1 U276 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U277 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U278 ( .A(n261), .Y(n307) );
  INVX1 U279 ( .A(n20), .Y(n326) );
  NAND2X1 U280 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U281 ( .A(n187), .Y(n196) );
  INVX1 U282 ( .A(n350), .Y(n335) );
  NAND2X1 U283 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U284 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U285 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U286 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U287 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U288 ( .A(n103), .Y(n37) );
  NOR2X1 U289 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U290 ( .A(n311), .Y(n268) );
  INVX1 U291 ( .A(n293), .Y(n209) );
  NOR2X1 U292 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U293 ( .A(n224), .Y(n235) );
  NAND2X1 U294 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U295 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U296 ( .A(n195), .Y(n142) );
  NAND2X1 U297 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U298 ( .A(n226), .Y(n253) );
  NAND2X1 U299 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U300 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U301 ( .A(n1), .Y(n301) );
  NAND2X1 U302 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U303 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U304 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U305 ( .A(n89), .Y(n340) );
  AOI211X1 U306 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U307 ( .A(n327), .Y(n248) );
  INVX1 U308 ( .A(n181), .Y(n109) );
  INVX1 U309 ( .A(n225), .Y(n302) );
  NAND2X1 U310 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U311 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U312 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U313 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U314 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U315 ( .A(n270), .Y(n107) );
  INVX1 U316 ( .A(n306), .Y(n145) );
  NAND4X1 U317 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U318 ( .A(n210), .Y(n236) );
  INVX1 U319 ( .A(n331), .Y(n78) );
  INVX1 U320 ( .A(n328), .Y(n314) );
  OAI21XL U321 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U322 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U323 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U324 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U325 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U326 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U327 ( .A(n186), .Y(n194) );
  NAND2X1 U328 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U329 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U330 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U331 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U332 ( .A(n72), .Y(n204) );
  OAI21XL U333 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  INVX1 U334 ( .A(n125), .Y(n319) );
  NAND2X1 U335 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U336 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U337 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U338 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U339 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U340 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U341 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U342 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U343 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U344 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U345 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U346 ( .A(n117), .Y(n188) );
  OAI21XL U347 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U348 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U349 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  NOR2X1 U350 ( .A(n248), .B(n142), .Y(n357) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule


module aes_sbox_18 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367;

  INVX1 U1 ( .A(n296), .Y(n354) );
  INVX1 U2 ( .A(a[3]), .Y(n31) );
  NOR2BX1 U3 ( .AN(n348), .B(n309), .Y(n246) );
  AOI21XL U4 ( .A0(n359), .A1(n223), .B0(n65), .Y(n91) );
  AOI211XL U5 ( .A0(n185), .A1(n184), .B0(n183), .C0(n182), .Y(n191) );
  INVX1 U6 ( .A(n116), .Y(n203) );
  NAND2X1 U7 ( .A(n194), .B(n274), .Y(n344) );
  INVX1 U8 ( .A(n324), .Y(n265) );
  AOI2BB2XL U9 ( .B0(n359), .B1(n289), .A0N(n288), .A1N(n287), .Y(n300) );
  AOI21XL U10 ( .A0(n339), .A1(n338), .B0(n337), .Y(n341) );
  NAND2XL U11 ( .A(n235), .B(n265), .Y(n338) );
  INVXL U12 ( .A(n257), .Y(n289) );
  NOR2XL U13 ( .A(n224), .B(n326), .Y(n257) );
  AOI22XL U14 ( .A0(n161), .A1(n327), .B0(n13), .B1(n265), .Y(n18) );
  NAND2XL U15 ( .A(n109), .B(n78), .Y(n158) );
  NOR2XL U16 ( .A(n324), .B(n131), .Y(n262) );
  NOR2X1 U17 ( .A(a[1]), .B(n293), .Y(n318) );
  NOR2X1 U18 ( .A(n293), .B(n323), .Y(n150) );
  NAND2XL U19 ( .A(a[1]), .B(n293), .Y(n82) );
  NAND2XL U20 ( .A(n140), .B(n20), .Y(n151) );
  NOR2XL U21 ( .A(n181), .B(n95), .Y(n174) );
  NOR2X4 U22 ( .A(n264), .B(n197), .Y(n350) );
  NOR2XL U23 ( .A(a[1]), .B(n242), .Y(n186) );
  NOR2X1 U24 ( .A(a[1]), .B(n103), .Y(n331) );
  INVXL U25 ( .A(n267), .Y(n333) );
  INVXL U26 ( .A(n352), .Y(n141) );
  NAND2X1 U27 ( .A(a[1]), .B(n31), .Y(n352) );
  AOI31XL U28 ( .A0(n260), .A1(n259), .A2(n258), .B0(n340), .Y(n282) );
  AOI211XL U29 ( .A0(n89), .A1(n88), .B0(n87), .C0(n86), .Y(n90) );
  AOI211XL U30 ( .A0(n125), .A1(n58), .B0(n57), .C0(n56), .Y(n59) );
  OR4X2 U31 ( .A(n367), .B(n366), .C(n365), .D(n364), .Y(d[0]) );
  AOI211XL U32 ( .A0(n125), .A1(n124), .B0(n123), .C0(n122), .Y(n126) );
  AOI211XL U33 ( .A0(n328), .A1(n257), .B0(n256), .C0(n255), .Y(n258) );
  AOI31XL U34 ( .A0(n322), .A1(n321), .A2(n320), .B0(n319), .Y(n366) );
  OAI211XL U35 ( .A0(n288), .A1(n265), .B0(n137), .C0(n136), .Y(n138) );
  AOI31XL U36 ( .A0(n55), .A1(n54), .A2(n53), .B0(n340), .Y(n56) );
  AOI31XL U37 ( .A0(n85), .A1(n84), .A2(n83), .B0(n297), .Y(n86) );
  AOI31XL U38 ( .A0(n25), .A1(n24), .A2(n23), .B0(n340), .Y(n26) );
  AOI31XL U39 ( .A0(n121), .A1(n120), .A2(n119), .B0(n340), .Y(n122) );
  AOI31XL U40 ( .A0(n19), .A1(n18), .A2(n17), .B0(n297), .Y(n27) );
  AOI22XL U41 ( .A0(n327), .A1(n203), .B0(n188), .B1(n118), .Y(n119) );
  AOI211XL U42 ( .A0(n327), .A1(n135), .B0(n134), .C0(n133), .Y(n136) );
  AOI31XL U43 ( .A0(n157), .A1(n156), .A2(n155), .B0(n319), .Y(n168) );
  AOI31XL U44 ( .A0(n166), .A1(n165), .A2(n164), .B0(n340), .Y(n167) );
  OAI211XL U45 ( .A0(n193), .A1(n192), .B0(n191), .C0(n190), .Y(n218) );
  AOI211XL U46 ( .A0(n257), .A1(n359), .B0(n15), .C0(n14), .Y(n17) );
  AOI211XL U47 ( .A0(n246), .A1(n236), .B0(n174), .C0(n52), .Y(n53) );
  AOI211XL U48 ( .A0(n328), .A1(n158), .B0(n81), .C0(n80), .Y(n84) );
  AOI22XL U49 ( .A0(n254), .A1(n296), .B0(n265), .B1(n102), .Y(n105) );
  AOI31XL U50 ( .A0(n300), .A1(n299), .A2(n298), .B0(n297), .Y(n367) );
  OAI211XL U51 ( .A0(n245), .A1(n354), .B0(n244), .C0(n243), .Y(n283) );
  AOI31XL U52 ( .A0(n343), .A1(n342), .A2(n341), .B0(n340), .Y(n365) );
  AOI22XL U53 ( .A0(n327), .A1(n223), .B0(n1), .B1(n222), .Y(n230) );
  OAI22XL U54 ( .A0(n254), .A1(n288), .B0(n253), .B1(n252), .Y(n255) );
  AOI211XL U55 ( .A0(n349), .A1(n203), .B0(n202), .C0(n201), .Y(n207) );
  AOI211XL U56 ( .A0(n318), .A1(n349), .B0(n317), .C0(n316), .Y(n320) );
  AOI211XL U57 ( .A0(a[7]), .A1(n338), .B0(n92), .C0(n111), .Y(n15) );
  INVXL U58 ( .A(n101), .Y(n254) );
  AOI211XL U59 ( .A0(a[2]), .A1(n130), .B0(n315), .C0(n129), .Y(n134) );
  AOI211XL U60 ( .A0(n350), .A1(n338), .B0(n357), .C0(n144), .Y(n147) );
  AOI211XL U61 ( .A0(n327), .A1(n289), .B0(n163), .C0(n162), .Y(n164) );
  OAI211XL U62 ( .A0(n336), .A1(n233), .B0(n177), .C0(n176), .Y(n178) );
  AOI31XL U63 ( .A0(n242), .A1(n253), .A2(n241), .B0(n240), .Y(n244) );
  OAI211XL U64 ( .A0(n70), .A1(n117), .B0(n69), .C0(n68), .Y(n88) );
  AOI211XL U65 ( .A0(n325), .A1(n184), .B0(n48), .C0(n163), .Y(n49) );
  NAND2XL U66 ( .A(n296), .B(n101), .Y(n94) );
  AOI31XL U67 ( .A0(n114), .A1(n113), .A2(n243), .B0(n360), .Y(n123) );
  AOI22XL U68 ( .A0(n1), .A1(n130), .B0(n359), .B1(n263), .Y(n9) );
  AOI31XL U69 ( .A0(n77), .A1(n76), .A2(n93), .B0(n319), .Y(n87) );
  OAI211XL U70 ( .A0(n249), .A1(n335), .B0(n64), .C0(n63), .Y(n65) );
  INVXL U71 ( .A(n150), .Y(n310) );
  AOI22XL U72 ( .A0(n66), .A1(n150), .B0(n350), .B1(n263), .Y(n69) );
  AOI22XL U73 ( .A0(n296), .A1(n150), .B0(n350), .B1(n262), .Y(n4) );
  AOI211XL U74 ( .A0(n1), .A1(n82), .B0(n47), .C0(n46), .Y(n50) );
  AOI31XL U75 ( .A0(n363), .A1(n362), .A2(n361), .B0(n360), .Y(n364) );
  AOI22XL U76 ( .A0(n1), .A1(n188), .B0(n359), .B1(n150), .Y(n157) );
  NAND2XL U77 ( .A(n235), .B(n274), .Y(n184) );
  NOR2XL U78 ( .A(n224), .B(n150), .Y(n116) );
  NOR2XL U79 ( .A(n150), .B(n331), .Y(n130) );
  AOI31XL U80 ( .A0(n215), .A1(n214), .A2(n213), .B0(n319), .Y(n216) );
  AOI211XL U81 ( .A0(n296), .A1(n175), .B0(n174), .C0(n173), .Y(n177) );
  AOI211XL U82 ( .A0(n350), .A1(n247), .B0(n246), .C0(n312), .Y(n260) );
  AOI221XL U83 ( .A0(n345), .A1(n329), .B0(n1), .B1(n266), .C0(n112), .Y(n113)
         );
  AOI22XL U84 ( .A0(n349), .A1(n305), .B0(n350), .B1(n38), .Y(n25) );
  NAND2XL U85 ( .A(n265), .B(n348), .Y(n247) );
  AOI2BB2XL U86 ( .B0(n350), .B1(n100), .A0N(n192), .A1N(n99), .Y(n106) );
  AOI211XL U87 ( .A0(n345), .A1(n265), .B0(n139), .C0(n115), .Y(n121) );
  AOI22XL U88 ( .A0(n188), .A1(n273), .B0(n233), .B1(n314), .Y(n189) );
  AOI22XL U89 ( .A0(n349), .A1(n210), .B0(n328), .B1(n265), .Y(n54) );
  AOI2BB2XL U90 ( .B0(n350), .B1(n82), .A0N(n233), .A1N(n100), .Y(n51) );
  AOI22XL U91 ( .A0(n349), .A1(n287), .B0(n345), .B1(n266), .Y(n153) );
  AOI211XL U92 ( .A0(n296), .A1(n287), .B0(n75), .C0(n74), .Y(n76) );
  AOI22XL U93 ( .A0(n350), .A1(n158), .B0(n328), .B1(n175), .Y(n166) );
  AOI22XL U94 ( .A0(n329), .A1(n1), .B0(n296), .B1(n135), .Y(n64) );
  OAI22XL U95 ( .A0(n355), .A1(n353), .B0(n172), .B1(n180), .Y(n173) );
  AOI211XL U96 ( .A0(n328), .A1(n194), .B0(n67), .C0(n139), .Y(n68) );
  INVXL U97 ( .A(n152), .Y(n222) );
  AOI22XL U98 ( .A0(n349), .A1(n100), .B0(n325), .B1(n172), .Y(n34) );
  AOI22XL U99 ( .A0(n349), .A1(n291), .B0(n256), .B1(n265), .Y(n79) );
  AOI22XL U100 ( .A0(n224), .A1(n328), .B0(n296), .B1(n99), .Y(n43) );
  AOI211XL U101 ( .A0(n328), .A1(n263), .B0(n212), .C0(n211), .Y(n214) );
  AOI22XL U102 ( .A0(n1), .A1(n40), .B0(n345), .B1(n287), .Y(n41) );
  AOI211XL U103 ( .A0(n359), .A1(n358), .B0(n357), .C0(n356), .Y(n361) );
  AOI211XL U104 ( .A0(n296), .A1(n351), .B0(n295), .C0(n294), .Y(n298) );
  AOI31XL U105 ( .A0(n327), .A1(n352), .A2(n351), .B0(n308), .Y(n321) );
  AOI2BB2XL U106 ( .B0(n327), .B1(n291), .A0N(n314), .A1N(n290), .Y(n299) );
  NOR2XL U107 ( .A(n209), .B(n233), .Y(n256) );
  NAND3XL U108 ( .A(n1), .B(n140), .C(n82), .Y(n83) );
  AOI22XL U109 ( .A0(n327), .A1(n117), .B0(n328), .B1(n151), .Y(n24) );
  AOI2BB2XL U110 ( .B0(n261), .B1(n359), .A0N(n288), .A1N(n262), .Y(n280) );
  AOI22XL U111 ( .A0(n185), .A1(n318), .B0(n327), .B1(n262), .Y(n110) );
  NAND2XL U112 ( .A(n109), .B(n242), .Y(n135) );
  OAI22XL U113 ( .A0(n161), .A1(n301), .B0(n92), .B1(n233), .Y(n98) );
  OAI22XL U114 ( .A0(n31), .A1(n248), .B0(n197), .B1(n151), .Y(n36) );
  AOI22XL U115 ( .A0(n1), .A1(n226), .B0(n350), .B1(n221), .Y(n199) );
  AOI22XL U116 ( .A0(n327), .A1(n92), .B0(n345), .B1(n323), .Y(n45) );
  INVXL U117 ( .A(n82), .Y(n172) );
  AOI211XL U118 ( .A0(n327), .A1(n268), .B0(n62), .C0(n295), .Y(n63) );
  NOR2XL U119 ( .A(n293), .B(n292), .Y(n294) );
  AOI22XL U120 ( .A0(n195), .A1(n332), .B0(n328), .B1(n344), .Y(n208) );
  AOI32XL U121 ( .A0(n109), .A1(a[7]), .A2(n266), .B0(n159), .B1(n264), .Y(
        n193) );
  INVXL U122 ( .A(n312), .Y(n313) );
  NAND2XL U123 ( .A(n103), .B(n253), .Y(n305) );
  INVXL U124 ( .A(n180), .Y(n183) );
  AOI211XL U125 ( .A0(n288), .A1(n301), .B0(n181), .C0(n261), .Y(n182) );
  AOI22XL U126 ( .A0(n1), .A1(n263), .B0(n328), .B1(n262), .Y(n279) );
  AOI22XL U127 ( .A0(n349), .A1(n20), .B0(n345), .B1(n318), .Y(n5) );
  AOI22XL U128 ( .A0(n296), .A1(n142), .B0(n350), .B1(n159), .Y(n85) );
  AOI2BB2XL U129 ( .B0(n350), .B1(n336), .A0N(n288), .A1N(n175), .Y(n44) );
  AOI22XL U130 ( .A0(n268), .A1(n350), .B0(n327), .B1(n151), .Y(n156) );
  OAI2BB1XL U131 ( .A0N(n210), .A1N(n325), .B0(n243), .Y(n211) );
  OAI211XL U132 ( .A0(n274), .A1(n273), .B0(n272), .C0(n271), .Y(n276) );
  AOI22XL U133 ( .A0(n327), .A1(n39), .B0(n359), .B1(n38), .Y(n42) );
  NAND2XL U134 ( .A(n352), .B(n351), .Y(n358) );
  AOI22XL U135 ( .A0(n92), .A1(n349), .B0(n350), .B1(n303), .Y(n77) );
  NOR2XL U136 ( .A(n161), .B(n309), .Y(n162) );
  AOI22XL U137 ( .A0(n1), .A1(n346), .B0(n345), .B1(n344), .Y(n363) );
  AOI22XL U138 ( .A0(n186), .A1(n359), .B0(n328), .B1(n103), .Y(n33) );
  AOI22XL U139 ( .A0(a[4]), .A1(n296), .B0(n345), .B1(n306), .Y(n21) );
  NOR2XL U140 ( .A(n268), .B(n354), .Y(n13) );
  AOI22XL U141 ( .A0(n349), .A1(n293), .B0(n296), .B1(n326), .Y(n11) );
  AOI22XL U142 ( .A0(n226), .A1(n205), .B0(n359), .B1(n311), .Y(n6) );
  AOI22XL U143 ( .A0(a[3]), .A1(n345), .B0(n327), .B1(n198), .Y(n200) );
  OAI22XL U144 ( .A0(n326), .A1(n233), .B0(n197), .B1(n196), .Y(n202) );
  NAND2XL U145 ( .A(n350), .B(n245), .Y(n180) );
  NAND2XL U146 ( .A(n311), .B(n236), .Y(n346) );
  AOI2BB2XL U147 ( .B0(n359), .B1(n160), .A0N(n301), .A1N(n159), .Y(n165) );
  AOI22XL U148 ( .A0(a[3]), .A1(n350), .B0(n349), .B1(n348), .Y(n362) );
  AOI22XL U149 ( .A0(n268), .A1(n359), .B0(n339), .B1(n331), .Y(n143) );
  AOI22XL U150 ( .A0(a[1]), .A1(n296), .B0(n1), .B1(n140), .Y(n149) );
  AOI22XL U151 ( .A0(n296), .A1(n128), .B0(n359), .B1(n306), .Y(n137) );
  INVXL U152 ( .A(n131), .Y(n351) );
  NOR3XL U153 ( .A(n181), .B(n261), .C(n309), .Y(n295) );
  NOR3XL U154 ( .A(n324), .B(n249), .C(n248), .Y(n250) );
  NOR2XL U155 ( .A(n181), .B(n269), .Y(n315) );
  AOI22XL U156 ( .A0(n327), .A1(n290), .B0(n333), .B1(n350), .Y(n237) );
  AOI22XL U157 ( .A0(n349), .A1(n226), .B0(n249), .B1(n328), .Y(n229) );
  AND2X2 U158 ( .A(n303), .B(n78), .Y(n221) );
  AOI22XL U159 ( .A0(a[1]), .A1(n350), .B0(n349), .B1(n333), .Y(n215) );
  AOI31XL U160 ( .A0(n354), .A1(n233), .A2(n176), .B0(n329), .Y(n67) );
  AOI211XL U161 ( .A0(a[7]), .A1(n61), .B0(n187), .C0(n111), .Y(n62) );
  NAND2XL U162 ( .A(n311), .B(n196), .Y(n40) );
  NOR2XL U163 ( .A(n293), .B(n226), .Y(n39) );
  AOI22XL U164 ( .A0(n226), .A1(n350), .B0(n339), .B1(n355), .Y(n120) );
  OAI22XL U165 ( .A0(n354), .A1(n194), .B0(n306), .B1(n314), .Y(n115) );
  AOI22XL U166 ( .A0(n350), .A1(n352), .B0(n108), .B1(n107), .Y(n114) );
  NOR2XL U167 ( .A(n37), .B(n145), .Y(n99) );
  AOI22XL U168 ( .A0(n181), .A1(n350), .B0(n328), .B1(n269), .Y(n96) );
  NOR2XL U169 ( .A(a[1]), .B(n249), .Y(n131) );
  NAND2XL U170 ( .A(n311), .B(n303), .Y(n38) );
  NOR2XL U171 ( .A(n233), .B(n331), .Y(n108) );
  AOI22XL U172 ( .A0(n325), .A1(n324), .B0(n1), .B1(n323), .Y(n343) );
  NAND3XL U173 ( .A(n1), .B(a[3]), .C(n204), .Y(n73) );
  NAND2XL U174 ( .A(n107), .B(n348), .Y(n175) );
  NOR2XL U175 ( .A(n37), .B(a[1]), .Y(n195) );
  AOI22XL U176 ( .A0(n141), .A1(n332), .B0(n251), .B1(n330), .Y(n148) );
  NOR2XL U177 ( .A(a[1]), .B(n329), .Y(n269) );
  AOI22XL U178 ( .A0(n187), .A1(n205), .B0(n328), .B1(n307), .Y(n12) );
  NAND2XL U179 ( .A(n329), .B(n323), .Y(n245) );
  AOI22XL U180 ( .A0(n268), .A1(n325), .B0(n330), .B1(n267), .Y(n272) );
  AOI22XL U181 ( .A0(n333), .A1(n332), .B0(n331), .B1(n330), .Y(n334) );
  NOR2XL U182 ( .A(n187), .B(n186), .Y(n290) );
  NAND3XL U183 ( .A(n205), .B(n242), .C(n204), .Y(n206) );
  NAND2XL U184 ( .A(n306), .B(n267), .Y(n61) );
  AOI22XL U185 ( .A0(n329), .A1(n328), .B0(n327), .B1(n326), .Y(n342) );
  NAND2XL U186 ( .A(n328), .B(n311), .Y(n353) );
  NAND2XL U187 ( .A(a[1]), .B(n261), .Y(n303) );
  INVXL U188 ( .A(n197), .Y(n185) );
  NAND3XL U189 ( .A(n332), .B(n72), .C(n242), .Y(n71) );
  INVXL U190 ( .A(n297), .Y(n284) );
  INVXL U191 ( .A(n332), .Y(n234) );
  AOI22XL U192 ( .A0(a[2]), .A1(a[4]), .B0(a[3]), .B1(n273), .Y(n132) );
  NOR2XL U193 ( .A(a[1]), .B(n198), .Y(n160) );
  AOI22XL U194 ( .A0(a[1]), .A1(a[7]), .B0(n264), .B1(n323), .Y(n72) );
  INVXL U195 ( .A(n274), .Y(n251) );
  NAND2XL U196 ( .A(n264), .B(n275), .Y(n252) );
  NOR2XL U197 ( .A(n264), .B(n273), .Y(n330) );
  INVX2 U198 ( .A(a[7]), .Y(n264) );
  NAND2XL U199 ( .A(a[4]), .B(a[1]), .Y(n274) );
  NAND2XL U200 ( .A(a[3]), .B(a[1]), .Y(n20) );
  NOR2XL U201 ( .A(a[3]), .B(a[1]), .Y(n225) );
  CLKINVX3 U202 ( .A(n266), .Y(n329) );
  NAND2X2 U203 ( .A(a[4]), .B(n31), .Y(n266) );
  OAI21X1 U204 ( .A0(n60), .A1(n297), .B0(n59), .Y(d[6]) );
  OAI21X1 U205 ( .A0(n286), .A1(n319), .B0(n285), .Y(d[1]) );
  OAI21X1 U206 ( .A0(n127), .A1(n297), .B0(n126), .Y(d[4]) );
  NAND2X2 U207 ( .A(n275), .B(n273), .Y(n197) );
  CLKINVX3 U208 ( .A(a[5]), .Y(n275) );
  NOR2X2 U209 ( .A(n31), .B(n198), .Y(n261) );
  NOR2X2 U210 ( .A(n37), .B(n323), .Y(n181) );
  NOR2X2 U211 ( .A(n273), .B(a[7]), .Y(n325) );
  NOR2X2 U212 ( .A(n249), .B(n329), .Y(n293) );
  NOR2X2 U213 ( .A(n329), .B(n323), .Y(n226) );
  NAND2X2 U214 ( .A(n198), .B(n323), .Y(n311) );
  CLKINVX3 U215 ( .A(a[4]), .Y(n198) );
  CLKINVX3 U216 ( .A(n233), .Y(n359) );
  NAND2X2 U217 ( .A(a[5]), .B(n325), .Y(n233) );
  CLKINVX3 U218 ( .A(n349), .Y(n288) );
  NOR2X4 U219 ( .A(a[7]), .B(n111), .Y(n349) );
  NOR2X4 U220 ( .A(n264), .B(n192), .Y(n327) );
  NOR2X4 U221 ( .A(a[2]), .B(n129), .Y(n328) );
  BUFX3 U222 ( .A(n347), .Y(n1) );
  CLKINVX3 U223 ( .A(a[2]), .Y(n273) );
  OAI21X1 U224 ( .A0(n220), .A1(n340), .B0(n219), .Y(d[2]) );
  NOR2X4 U225 ( .A(a[7]), .B(n197), .Y(n296) );
  OAI21X1 U226 ( .A0(n171), .A1(n360), .B0(n170), .Y(d[3]) );
  OAI21X1 U227 ( .A0(n91), .A1(n360), .B0(n90), .Y(d[5]) );
  OAI21X1 U228 ( .A0(n30), .A1(n360), .B0(n29), .Y(d[7]) );
  AOI31X4 U229 ( .A0(n208), .A1(n207), .A2(n206), .B0(n360), .Y(n217) );
  AOI31X4 U230 ( .A0(n280), .A1(n279), .A2(n278), .B0(n360), .Y(n281) );
  CLKINVX3 U231 ( .A(n309), .Y(n345) );
  NAND2X2 U232 ( .A(n275), .B(n325), .Y(n309) );
  NAND2X2 U233 ( .A(a[1]), .B(n242), .Y(n306) );
  NAND2X2 U234 ( .A(a[3]), .B(n198), .Y(n242) );
  AOI21XL U235 ( .A0(n50), .A1(n49), .B0(n360), .Y(n57) );
  AOI21XL U236 ( .A0(n236), .A1(n78), .B0(n314), .Y(n47) );
  AOI21XL U237 ( .A0(n266), .A1(n265), .B0(n264), .Y(n277) );
  AOI21XL U238 ( .A0(n251), .A1(n1), .B0(n250), .Y(n259) );
  AOI21XL U239 ( .A0(n345), .A1(n346), .B0(n238), .Y(n239) );
  AOI21XL U240 ( .A0(n209), .A1(n306), .B0(n248), .Y(n212) );
  AOI21XL U241 ( .A0(n267), .A1(n352), .B0(n309), .Y(n179) );
  AOI21XL U242 ( .A0(n311), .A1(n310), .B0(n309), .Y(n317) );
  AOI21XL U243 ( .A0(n307), .A1(n306), .B0(n335), .Y(n308) );
  AOI21XL U244 ( .A0(n359), .A1(n305), .B0(n304), .Y(n322) );
  AOI21XL U245 ( .A0(n303), .A1(n302), .B0(n301), .Y(n304) );
  AOI21XL U246 ( .A0(n350), .A1(n306), .B0(n1), .Y(n292) );
  AOI21XL U247 ( .A0(n236), .A1(n245), .B0(n248), .Y(n81) );
  AOI21XL U248 ( .A0(n205), .A1(n318), .B0(n345), .Y(n70) );
  AOI21XL U249 ( .A0(n328), .A1(n222), .B0(n154), .Y(n155) );
  AOI21XL U250 ( .A0(n132), .A1(n351), .B0(n309), .Y(n133) );
  AOI21XL U251 ( .A0(n359), .A1(n287), .B0(n22), .Y(n23) );
  AOI21XL U252 ( .A0(n142), .A1(n352), .B0(n335), .Y(n14) );
  AOI21XL U253 ( .A0(n327), .A1(n247), .B0(n48), .Y(n10) );
  AOI21XL U254 ( .A0(n311), .A1(n196), .B0(n335), .Y(n48) );
  NOR2X1 U255 ( .A(n273), .B(n129), .Y(n347) );
  CLKINVX3 U256 ( .A(a[1]), .Y(n323) );
  NAND2X1 U257 ( .A(a[7]), .B(a[5]), .Y(n129) );
  NOR2X1 U258 ( .A(n323), .B(n242), .Y(n210) );
  NAND2X1 U259 ( .A(a[2]), .B(n275), .Y(n192) );
  NAND2X1 U260 ( .A(n327), .B(n266), .Y(n95) );
  NOR2X1 U261 ( .A(a[4]), .B(n323), .Y(n270) );
  OAI21XL U262 ( .A0(n270), .A1(n225), .B0(n1), .Y(n3) );
  NOR2X1 U263 ( .A(a[2]), .B(n275), .Y(n66) );
  NOR2X1 U264 ( .A(a[7]), .B(a[2]), .Y(n339) );
  INVX1 U265 ( .A(n242), .Y(n249) );
  OAI21XL U266 ( .A0(n66), .A1(n339), .B0(n131), .Y(n2) );
  NAND3X1 U267 ( .A(n95), .B(n3), .C(n2), .Y(n8) );
  INVX1 U268 ( .A(n192), .Y(n205) );
  INVX1 U269 ( .A(n66), .Y(n111) );
  NOR2X1 U270 ( .A(n261), .B(n323), .Y(n324) );
  NAND3X1 U271 ( .A(n6), .B(n5), .C(n4), .Y(n7) );
  AOI211X1 U272 ( .A0(n328), .A1(n210), .B0(n8), .C0(n7), .Y(n30) );
  NAND2X1 U273 ( .A(a[6]), .B(a[0]), .Y(n360) );
  INVX1 U274 ( .A(a[6]), .Y(n16) );
  NOR2X1 U275 ( .A(a[0]), .B(n16), .Y(n125) );
  NOR2X1 U276 ( .A(n323), .B(n266), .Y(n187) );
  INVX1 U277 ( .A(n261), .Y(n307) );
  INVX1 U278 ( .A(n20), .Y(n326) );
  NAND2X1 U279 ( .A(n261), .B(n323), .Y(n348) );
  INVX1 U280 ( .A(n187), .Y(n196) );
  INVX1 U281 ( .A(n350), .Y(n335) );
  NAND2X1 U282 ( .A(n31), .B(n198), .Y(n103) );
  NAND2X1 U283 ( .A(n20), .B(n245), .Y(n263) );
  NAND4X1 U284 ( .A(n12), .B(n11), .C(n10), .D(n9), .Y(n28) );
  NAND2X1 U285 ( .A(a[3]), .B(n323), .Y(n267) );
  AOI22X1 U286 ( .A0(n1), .A1(n39), .B0(n345), .B1(n61), .Y(n19) );
  INVX1 U287 ( .A(n103), .Y(n37) );
  NOR2X1 U288 ( .A(n195), .B(n270), .Y(n161) );
  INVX1 U289 ( .A(n311), .Y(n268) );
  INVX1 U290 ( .A(n293), .Y(n209) );
  NOR2X1 U291 ( .A(a[1]), .B(n209), .Y(n224) );
  INVX1 U292 ( .A(n224), .Y(n235) );
  NAND2X1 U293 ( .A(n323), .B(n307), .Y(n140) );
  NOR2BX1 U294 ( .AN(n140), .B(n181), .Y(n92) );
  INVX1 U295 ( .A(n195), .Y(n142) );
  NAND2X1 U296 ( .A(a[0]), .B(n16), .Y(n297) );
  INVX1 U297 ( .A(n226), .Y(n253) );
  NAND2X1 U298 ( .A(n196), .B(n348), .Y(n117) );
  NAND2X1 U299 ( .A(n307), .B(n82), .Y(n287) );
  INVX1 U300 ( .A(n1), .Y(n301) );
  NAND2X1 U301 ( .A(n235), .B(n352), .Y(n101) );
  OAI21XL U302 ( .A0(n301), .A1(n101), .B0(n21), .Y(n22) );
  NOR2X1 U303 ( .A(a[6]), .B(a[0]), .Y(n89) );
  INVX1 U304 ( .A(n89), .Y(n340) );
  AOI211X1 U305 ( .A0(n125), .A1(n28), .B0(n27), .C0(n26), .Y(n29) );
  INVX1 U306 ( .A(n327), .Y(n248) );
  INVX1 U307 ( .A(n181), .Y(n109) );
  INVX1 U308 ( .A(n225), .Y(n302) );
  NAND2X1 U309 ( .A(n109), .B(n302), .Y(n100) );
  OAI21XL U310 ( .A0(n270), .A1(n160), .B0(n1), .Y(n32) );
  NAND4BXL U311 ( .AN(n246), .B(n34), .C(n33), .D(n32), .Y(n35) );
  AOI211X1 U312 ( .A0(n296), .A1(n101), .B0(n36), .C0(n35), .Y(n60) );
  NOR2X1 U313 ( .A(n141), .B(n331), .Y(n336) );
  INVX1 U314 ( .A(n270), .Y(n107) );
  INVX1 U315 ( .A(n306), .Y(n145) );
  NAND4X1 U316 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n58) );
  INVX1 U317 ( .A(n210), .Y(n236) );
  INVX1 U318 ( .A(n331), .Y(n78) );
  INVX1 U319 ( .A(n328), .Y(n314) );
  OAI21XL U320 ( .A0(a[4]), .A1(n288), .B0(n45), .Y(n46) );
  NAND2X1 U321 ( .A(n311), .B(n253), .Y(n291) );
  NOR2X1 U322 ( .A(n354), .B(n291), .Y(n163) );
  OAI21XL U323 ( .A0(n324), .A1(n225), .B0(n296), .Y(n55) );
  OAI21XL U324 ( .A0(n116), .A1(n301), .B0(n51), .Y(n52) );
  NAND2X1 U325 ( .A(n267), .B(n310), .Y(n223) );
  INVX1 U326 ( .A(n186), .Y(n194) );
  NAND2X1 U327 ( .A(n1), .B(n311), .Y(n176) );
  NOR2X1 U328 ( .A(n288), .B(n311), .Y(n139) );
  NOR2X1 U329 ( .A(n275), .B(n273), .Y(n332) );
  OAI21XL U330 ( .A0(n352), .A1(n248), .B0(n71), .Y(n75) );
  INVX1 U331 ( .A(n72), .Y(n204) );
  OAI21XL U332 ( .A0(n221), .A1(n314), .B0(n73), .Y(n74) );
  NAND2X1 U333 ( .A(n345), .B(n209), .Y(n93) );
  INVX1 U334 ( .A(n125), .Y(n319) );
  NAND2X1 U335 ( .A(n107), .B(n267), .Y(n159) );
  OAI21XL U336 ( .A0(n116), .A1(n309), .B0(n79), .Y(n80) );
  NOR2X1 U337 ( .A(n145), .B(n318), .Y(n152) );
  NAND4X1 U338 ( .A(n96), .B(n95), .C(n94), .D(n93), .Y(n97) );
  AOI211X1 U339 ( .A0(n349), .A1(n152), .B0(n98), .C0(n97), .Y(n127) );
  OAI21XL U340 ( .A0(n249), .A1(n288), .B0(n176), .Y(n102) );
  NOR2X1 U341 ( .A(n103), .B(n323), .Y(n355) );
  OAI21XL U342 ( .A0(n186), .A1(n355), .B0(n328), .Y(n104) );
  NAND4BXL U343 ( .AN(n108), .B(n106), .C(n105), .D(n104), .Y(n124) );
  OAI21XL U344 ( .A0(n111), .A1(n193), .B0(n110), .Y(n112) );
  NAND2X1 U345 ( .A(n296), .B(n226), .Y(n243) );
  INVX1 U346 ( .A(n117), .Y(n188) );
  OAI21XL U347 ( .A0(n194), .A1(n234), .B0(n233), .Y(n118) );
  OAI21XL U348 ( .A0(a[1]), .A1(n132), .B0(n306), .Y(n128) );
  AOI211X1 U349 ( .A0(n188), .A1(n350), .B0(n139), .C0(n138), .Y(n171) );
  NOR2X1 U350 ( .A(n248), .B(n142), .Y(n357) );
  OAI21XL U351 ( .A0(n309), .A1(n302), .B0(n143), .Y(n144) );
  OAI21XL U352 ( .A0(n329), .A1(n145), .B0(n328), .Y(n146) );
  NAND4X1 U353 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n169) );
  OAI21XL U354 ( .A0(n209), .A1(n252), .B0(n153), .Y(n154) );
  AOI211X1 U355 ( .A0(n284), .A1(n169), .B0(n168), .C0(n167), .Y(n170) );
  AOI211X1 U356 ( .A0(n349), .A1(n306), .B0(n179), .C0(n178), .Y(n220) );
  OAI21XL U357 ( .A0(n290), .A1(n273), .B0(n189), .Y(n190) );
  OAI21XL U358 ( .A0(n200), .A1(n204), .B0(n199), .Y(n201) );
  OAI21XL U359 ( .A0(n318), .A1(n355), .B0(n1), .Y(n213) );
  AOI211X1 U360 ( .A0(n284), .A1(n218), .B0(n217), .C0(n216), .Y(n219) );
  NOR2X1 U361 ( .A(n221), .B(n335), .Y(n232) );
  OAI21XL U362 ( .A0(n224), .A1(n270), .B0(n345), .Y(n228) );
  OAI21XL U363 ( .A0(n226), .A1(n225), .B0(n359), .Y(n227) );
  NAND4X1 U364 ( .A(n230), .B(n229), .C(n228), .D(n227), .Y(n231) );
  AOI211X1 U365 ( .A0(n336), .A1(n296), .B0(n232), .C0(n231), .Y(n286) );
  OAI21XL U366 ( .A0(n235), .A1(n234), .B0(n233), .Y(n241) );
  OAI21XL U367 ( .A0(n329), .A1(n314), .B0(n237), .Y(n238) );
  OAI21XL U368 ( .A0(n288), .A1(n346), .B0(n239), .Y(n240) );
  NOR2X1 U369 ( .A(n354), .B(n302), .Y(n312) );
  OAI21XL U370 ( .A0(n270), .A1(n269), .B0(n339), .Y(n271) );
  OAI21XL U371 ( .A0(n277), .A1(n276), .B0(n275), .Y(n278) );
  AOI211X1 U372 ( .A0(n284), .A1(n283), .B0(n282), .C0(n281), .Y(n285) );
  OAI21XL U373 ( .A0(n315), .A1(n314), .B0(n313), .Y(n316) );
  OAI21XL U374 ( .A0(n336), .A1(n335), .B0(n334), .Y(n337) );
  OAI21XL U375 ( .A0(n355), .A1(n354), .B0(n353), .Y(n356) );
endmodule

//wddl nand
module WDDLNAND2X (A,B,clkinv,Y);
  input A, B,clkinv;
  output Y;
  wire Ainv, Binv, Apre, Bpre, Ainvpre, Binvpre, y, y_bar, y_buf, y_barinv;
  AND2XL U1 ( .A(A), .B(clkinv), .Y(Apre));
  AND2XL U2 ( .A(B), .B(clkinv), .Y(Bpre));
  INVXL U3 ( .A(A), .Y(Ainv) );
  INVXL U4 ( .A(B), .Y(Binv) );
  AND2XL U5 ( .A(Ainv), .B(clkinv), .Y(Ainvpre));
  AND2XL U6 ( .A(Binv), .B(clkinv), .Y(Binvpre));
  AND2XL U7 ( .A(Apre), .B(Bpre), .Y(y_bar));
  OR2XL U8 ( .A(Ainvpre), .B(Binvpre), .Y(y));
  BUFXL U9 ( .A(y), .Y(y_buf) );
  INVXL U10 ( .A(y_bar), .Y(y_barinv));
  OR2XL U11 ( .A(y_buf), .B(y_barinv), .Y(Y));
  
  
endmodule

//wddl nor
module WDDLNOR2X (A,B,clkinv,Y);
  input A, B,clkinv;
  output Y;
  wire Ainv, Binv, Apre, Bpre, Ainvpre, Binvpre, y, y_bar, y_buf, y_barinv;
  AND2XL U1 ( .A(A), .B(clkinv), .Y(Apre));
  AND2XL U2 ( .A(B), .B(clkinv), .Y(Bpre));
  INVXL U3 ( .A(A), .Y(Ainv) );
  INVXL U4 ( .A(B), .Y(Binv) );
  AND2XL U5 ( .A(Ainv), .B(clkinv), .Y(Ainvpre));
  AND2XL U6 ( .A(Binv), .B(clkinv), .Y(Binvpre));
  OR2XL U7 ( .A(Apre), .B(Bpre), .Y(y_bar));
  AND2XL U8 ( .A(Ainvpre), .B(Binvpre), .Y(y));
  BUFXL U9 ( .A(y), .Y(y_buf) );
  INVXL U10 ( .A(y_bar), .Y(y_barinv));
  OR2XL U11 ( .A(y_buf), .B(y_barinv), .Y(Y));
  
  
endmodule

//wddl inv 
module WDDLINV (A,clkinv,Y);
  input A, clkinv;
  output Y;
  wire Ainv, y_bar, y, y_barinv, y_buf;
  AND2XL U1 ( .A(A), .B(clkinv), .Y(y_bar));
  INVXL U2 ( .A(A), .Y(Ainv) );
  AND2XL U3 ( .A(Ainv), .B(clkinv), .Y(y));
  BUFXL U4 ( .A(y), .Y(y_buf) );
  INVXL U5 ( .A(y_bar), .Y(y_barinv));
  OR2XL U6 ( .A(y_buf), .B(y_barinv), .Y(Y));

endmodule


//wddl: mux
module MUX2X(S, A, B, Y);
  input S, A, B;
  output Y;
  wire z1, z2, Sinv;
  AND2XL U1 ( .A(A), .B(S), .Y(z1));
  INVXL U2 ( .A(S), .Y(Sinv) );
  AND2XL U3 ( .A(B), .B(Sinv), .Y(z2));
  OR2XL U4 ( .A(z1), .B(z2), .Y(Y));
endmodule

//m master slave DFF
module WDDLDFFMS ( D,CK,Q );
  input D, CK;
  output Q; 
  wire z;
  DFFHQX1 reg_1 ( .D(D), .CK(CK), .Q(z));
  DFFHQX1 reg_2 ( .D(z), .CK(CK), .Q(Q));
  
endmodule

// WDDL register with DFF
/*
module WDDLDFFHQX2 ( D, Dinv, CLK, PRECLK, Q );
  input D, Dinv, CLK, PRECLK;
  output Q;
  wire q, qinv,z, zinv, clkinv,preclkinv, qpre, qinvpre, qbuf, qbarinv;
  //wire dinv, clkinv, qpre, qinvpre, qbuf, qbarinv;
  //reg q, qinv;
//  INVX1 U1 ( .A(D), .Y(Dinv));
  DFFHQX1 reg_11 ( .D(D), .CK(CLK), .Q(z));
  DFFHQX1 reg_12 ( .D(z), .CK(CLK), .Q(q));
  DFFHQX1 reg_21 ( .D(Dinv), .CK(CLK), .Q(zinv));
  DFFHQX1 reg_22 ( .D(zinv), .CK(CLK), .Q(qinv));
  CLKINVX1 U2 ( .A(PRECLK), .Y(preclkinv));
//  AND2X1 U3 ( .A(q), .B(preclkinv), .Y(qpre));
//  AND2X1 U4 ( .A(qinv), .B(preclkinv), .Y(qinvpre));
  BUFX1 U5 ( .A(q), .Y(qbuf));
  INVX1 U6 ( .A(qinv), .Y(qbarinv));
  OR2X1 U7 ( .A(qbuf), .B(qbarinv), .Y(Q));
endmodule */

//module WDDLDFFHQX2 ( D, Dinv, CLK, PRECLK, Q );
//  input D, Dinv, CLK, PRECLK;
//  output Q;
//  wire q, qinv,z, zinv, qpre, qinvpre, qbuf, qbarinv;
// // assign qpre = PRECLK?q:z;
//  //assign qinvpre = PRECLK?qinv:zinv;
//  //wire dinv, clkinv, qpre, qinvpre, qbuf, qbarinv;
//  //reg q, qinv;
////  INVX1 U1 ( .A(D), .Y(Dinv));
//  DFFHQX1 reg_11 ( .D(D), .CK(CLK), .Q(z));
//  DFFHQX1 reg_12 ( .D(z), .CK(CLK), .Q(q));
//  DFFHQX1 reg_21 ( .D(Dinv), .CK(CLK), .Q(zinv));
//  DFFHQX1 reg_22 ( .D(zinv), .CK(CLK), .Q(qinv));
////  CLKINVX1 U2 ( .A(PRECLK), .Y(preclkinv));
//  MUX2X m1 (.S(PRECLK), .A(z), .B(q), .Y(qpre));
//  MUX2X m2 (.S(PRECLK), .A(zinv), .B(qinv), .Y(qinvpre));
////  AND2X1 U3 ( .A(q), .B(preclkinv), .Y(qpre));
////  AND2X1 U4 ( .A(qinv), .B(preclkinv), .Y(qinvpre));
//  BUFX1 U5 ( .A(qpre), .Y(qbuf));
//  INVX1 U6 ( .A(qinvpre), .Y(qbarinv));
//  OR2X1 U7 ( .A(qbuf), .B(qbarinv), .Y(Q));
//endmodule

module WDDLDFFHQX2 ( D, Dinv, CLK, PRECLK, Q );
  input D, Dinv, CLK, PRECLK;
  output Q;
  wire q, qinv,z, zinv, qpre, qinvpre, qbuf, qbarinv, preclkinv, qmux, qinvmux;
 // assign qpre = PRECLK?q:z;
  //assign qinvpre = PRECLK?qinv:zinv;
  //wire dinv, clkinv, qpre, qinvpre, qbuf, qbarinv;
  //reg q, qinv;
//  INVX1 U1 ( .A(D), .Y(Dinv));
  DFFHQX1 reg_11 ( .D(D), .CK(CLK), .Q(z));
  DFFHQX1 reg_12 ( .D(z), .CK(CLK), .Q(q));
  DFFHQX1 reg_21 ( .D(Dinv), .CK(CLK), .Q(zinv));
  DFFHQX1 reg_22 ( .D(zinv), .CK(CLK), .Q(qinv));
  CLKINVX1 U2 ( .A(PRECLK), .Y(preclkinv));
//  MUX2X m1 (.S(PRECLK), .A(z), .B(q), .Y(qmux));
//  MUX2X m2 (.S(PRECLK), .A(zinv), .B(qinv), .Y(qinvmux));
  AND2X1 U3 ( .A(q), .B(preclkinv), .Y(qpre));
  AND2X1 U4 ( .A(qinv), .B(preclkinv), .Y(qinvpre));
  BUFX1 U5 ( .A(qpre), .Y(qbuf));
  INVX1 U6 ( .A(qinvpre), .Y(qbarinv));
  OR2X1 U7 ( .A(qbuf), .B(qbarinv), .Y(Q));
endmodule

// wddl precharge signal, half the clock signal

module precharge(clk,rst, preclk);
  input clk, rst;
  output preclk;
  wire q_bar;

 // DFFHQX1 reg_1 ( .D(d), .CK(clk), .Q(q));
  DFFRX4 reg_1 (.D(q_bar), .CK(clk), .Q(preclk), .QN(q_bar), .RN(rst));
  //CLKINVX1 U2 ( .A(q), .Y(d));
endmodule


module WDDLNANDCOMP ( A, B , C, clkinv, Y, Y_bar);
  input A, B, C, clkinv;
  output Y, Y_bar;
  wire Ainv, Binv, Apre, Bpre, Ainvpre, Binvpre, z, z_bar, Cpre, Cinvpre, Cinv;
  AND2X1 U1 ( .A(A), .B(clkinv), .Y(Apre));
  AND2X1 U2 ( .A(B), .B(clkinv), .Y(Bpre));
  AND2X1 U3 ( .A(C), .B(clkinv), .Y(Cpre));
  INVX1 U4 ( .A(A), .Y(Ainv) );
  INVX1 U5 ( .A(B), .Y(Binv) );
  INVX1 U6 ( .A(C), .Y(Cinv) );
  AND2X1 U7 ( .A(Ainv), .B(clkinv), .Y(Ainvpre));
  AND2X1 U8 ( .A(Binv), .B(clkinv), .Y(Binvpre));
  AND2X1 U9 ( .A(Cinv), .B(clkinv), .Y(Cinvpre));
  AND2X1 U10 ( .A(Apre), .B(Bpre), .Y(z_bar));
  OR2X1 U11 ( .A(Ainvpre), .B(Binvpre), .Y(z));
  AND2X1 U12 ( .A(z), .B(Cpre), .Y(Y_bar));
  OR2X1 U13 ( .A(z_bar), .B(Cinvpre), .Y(Y));
endmodule


//module aes_cipher_top ( clk, rst, ld, done, key, text_in, text_out );
//module aes_cipher_top ( clk, rst, ld, done, key, text_in, text_out );
module aes_cipher_top ( divclk,clk, rst, ld, done, key, text_in, text_out, m_in0_U179, m_in1_U179, m_out_U179, precharge_lmdpl);
  input [127:0] key;
  input [127:0] text_in;
  output [127:0] text_out;
  input divclk;
  // lmdpl inputs:
  input  m_in0_U179, m_in1_U179, m_out_U179, precharge_lmdpl;
  //input divclk, rst, ld;
  input clk, rst, ld;
  output done;
  wire   dcnt_2_, N21, N32, N33, N34, N35, N36, N37, N38, N39, N48, N49, N50,
         N51, N52, N53, N54, N55, N64, N65, N66, N67, N68, N69, N70, N71, N80,
         N81, N82, N83, N84, N85, N86, N87, N96, N97, N98, N99, N100, N101,
         N102, N103, N112, N113, N114, N115, N116, N117, N118, N119, N128,
         N129, N130, N131, N132, N133, N134, N135, N144, N145, N146, N147,
         N148, N149, N150, N151, N160, N161, N162, N163, N164, N165, N166,
         N167, N176, N177, N178, N179, N180, N181, N182, N183, N192, N193,
         N194, N195, N196, N197, N198, N199, N208, N209, N210, N211, N212,
         N213, N214, N215, N224, N225, N226, N227, N228, N229, N230, N231,
         N240, N241, N242, N243, N244, N245, N246, N247, N256, N257, N258,
         N259, N260, N261, N262, N263, N272, N273, N274, N275, N276, N277,
         N278, N279, N376, N377, N378, N379, N380, N381, N382, N383, N384,
         N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395,
         N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406,
         N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417,
         N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428,
         N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439,
         N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450,
         N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461,
         N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472,
         N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483,
         N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494,
         N495, N496, N497, N498, N499, N500, N501, N502, N503, n2, n3, n4,
         n137, n139, n398, n399, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n472, n473, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n508, n509, n510, n511, n512, n513, n514, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n581, n582, n583, n584, n585, n586, n587, n588, n589, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n607,
         n608, n609, n610, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n652, n653, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n746,
         n747, n748, n749, n750, n751, n752, n753, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, preclk, N49inv, clk_originv, clk_bar;
  wire   [127:0] text_in_r;
  wire   [31:0] w3;
  wire   [7:0] sa33;
  wire   [7:0] sa33_next;
  wire   [7:0] sa23;
  wire   [7:0] sa23_next;
  wire   [7:0] sa13;
  wire   [7:1] sa13_next;
  wire   [7:0] sa03;
  wire   [7:0] sa03_next;
  wire   [31:0] w2;
  wire   [7:0] sa32;
  wire   [7:1] sa32_next;
  wire   [7:0] sa22;
  wire   [7:1] sa22_next;
  wire   [7:0] sa12;
  wire   [7:1] sa12_next;
  wire   [7:0] sa02;
  wire   [7:1] sa02_next;
  wire   [31:0] w1;
  wire   [7:0] sa31;
  wire   [7:1] sa31_next;
  wire   [7:0] sa21;
  wire   [7:1] sa21_next;
  wire   [7:0] sa11;
  wire   [7:1] sa11_next;
  wire   [7:0] sa01;
  wire   [7:1] sa01_next;
  wire   [31:0] w0;
  wire   [7:0] sa30;
  wire   [7:0] sa30_next;
  wire   [7:0] sa20;
  wire   [7:0] sa20_next;
  wire   [7:0] sa10;
  wire   [7:0] sa10_next;
  wire   [7:0] sa00;
  wire   [7:0] sa00_next;
  wire   [7:0] sa00_sr;
  wire   [7:0] sa01_sr;
  wire   [7:0] sa02_sr;
  wire   [7:0] sa03_sr;
  wire   [7:0] sa10_sr;
  wire   [7:0] sa11_sr;
  wire   [7:0] sa12_sr;
  wire   [7:0] sa13_sr;
  wire   [7:0] sa20_sr;
  wire   [7:0] sa21_sr;
  wire   [7:0] sa22_sr;
  wire   [7:0] sa23_sr;
  wire   [7:0] sa30_sr;
  wire   [7:0] sa31_sr;
  wire   [7:0] sa32_sr;
  wire   [7:0] sa33_sr;

  aes_key_expand_128 u0 ( .clk(divclk), .kld(ld), .key(key), .wo_0(w0), .wo_1(w1), 
        .wo_2(w2), .wo_3(w3) );
 // aes_key_expand_128 u0 ( .clk(preclk), .kld(ld), .key(key), .wo_0(w0), .wo_1(w1), 
       // .wo_2(w2), .wo_3(w3) );
  aes_sbox_19 us00 ( .a(sa00), .d(sa00_sr) );
  aes_sbox_18 us01 ( .a(sa01), .d(sa01_sr) );
  aes_sbox_17 us02 ( .a(sa02), .d(sa02_sr) );
  aes_sbox_16 us03 ( .a(sa03), .d(sa03_sr) );
  aes_sbox_15 us10 ( .a(sa10), .d(sa13_sr) );
  aes_sbox_14 us11 ( .a(sa11), .d(sa10_sr) );
  aes_sbox_13 us12 ( .a(sa12), .d(sa11_sr) );
  aes_sbox_12 us13 ( .a(sa13), .d(sa12_sr) );
  aes_sbox_11 us20 ( .a(sa20), .d(sa22_sr) );
  aes_sbox_10 us21 ( .a(sa21), .d(sa23_sr) );
  aes_sbox_9 us22 ( .a(sa22), .d(sa20_sr) );
  //aes_sbox_8 us23 ( .a(sa23), .d(sa21_sr) );
  //wddl
  //aes_sbox_8 us23 ( .a(sa23), .d(sa21_sr), .preclkbar(clk_bar));
  aes_sbox_8 us23 ( .a(sa23), .d(sa21_sr), .clk(clk), .rst(rst), .preclkbar(clk_bar), .m_in0_U179(m_in0_U179), .m_in1_U179(m_in1_U179), .m_out_U179(m_out_U179), .precharge_lmdpl(precharge_lmdpl));
  aes_sbox_7 us30 ( .a(sa30), .d(sa31_sr) );
  aes_sbox_6 us31 ( .a(sa31), .d(sa32_sr) );
  aes_sbox_5 us32 ( .a(sa32), .d(sa33_sr) );
  aes_sbox_4 us33 ( .a(sa33), .d(sa30_sr) );
 //wddl: generate precharge clock
 // assign clkinput = rst ? divclk : 1'b0;
 // CLKINVX3 Uinv (.A(clk), .Y(clk_originv));
 // precharge pre(.clk(clk), .preclk(divclk),.rst(rst));
  DFFTRX1 dcnt_reg_0_ ( .D(n139), .RN(n137), .CK(divclk), .Q(n959) );
  DFFHQX1 done_reg ( .D(N21), .CK(divclk), .Q(done) );
WDDLDFFMS text_out_reg_127_ ( .D(N376), .CK(clk), .Q(text_out[127]) );
WDDLDFFMS text_out_reg_126_ ( .D(N377), .CK(clk), .Q(text_out[126]) );
WDDLDFFMS text_out_reg_125_ ( .D(N378), .CK(clk), .Q(text_out[125]) );
WDDLDFFMS text_out_reg_124_ ( .D(N379), .CK(clk), .Q(text_out[124]) );
WDDLDFFMS text_out_reg_123_ ( .D(N380), .CK(clk), .Q(text_out[123]) );
WDDLDFFMS text_out_reg_122_ ( .D(N381), .CK(clk), .Q(text_out[122]) );
WDDLDFFMS text_out_reg_121_ ( .D(N382), .CK(clk), .Q(text_out[121]) );
WDDLDFFMS text_out_reg_120_ ( .D(N383), .CK(clk), .Q(text_out[120]) );
WDDLDFFMS text_out_reg_95_ ( .D(N384), .CK(clk), .Q(text_out[95]) );
WDDLDFFMS text_out_reg_94_ ( .D(N385), .CK(clk), .Q(text_out[94]) );
WDDLDFFMS text_out_reg_93_ ( .D(N386), .CK(clk), .Q(text_out[93]) );
WDDLDFFMS text_out_reg_92_ ( .D(N387), .CK(clk), .Q(text_out[92]) );
WDDLDFFMS text_out_reg_91_ ( .D(N388), .CK(clk), .Q(text_out[91]) );
WDDLDFFMS text_out_reg_90_ ( .D(N389), .CK(clk), .Q(text_out[90]) );
WDDLDFFMS text_out_reg_89_ ( .D(N390), .CK(clk), .Q(text_out[89]) );
WDDLDFFMS text_out_reg_88_ ( .D(N391), .CK(clk), .Q(text_out[88]) );
WDDLDFFMS text_out_reg_63_ ( .D(N392), .CK(clk), .Q(text_out[63]) );
WDDLDFFMS text_out_reg_62_ ( .D(N393), .CK(clk), .Q(text_out[62]) );
WDDLDFFMS text_out_reg_61_ ( .D(N394), .CK(clk), .Q(text_out[61]) );
WDDLDFFMS text_out_reg_60_ ( .D(N395), .CK(clk), .Q(text_out[60]) );
WDDLDFFMS text_out_reg_59_ ( .D(N396), .CK(clk), .Q(text_out[59]) );
WDDLDFFMS text_out_reg_58_ ( .D(N397), .CK(clk), .Q(text_out[58]) );
WDDLDFFMS text_out_reg_57_ ( .D(N398), .CK(clk), .Q(text_out[57]) );
WDDLDFFMS text_out_reg_56_ ( .D(N399), .CK(clk), .Q(text_out[56]) );
WDDLDFFMS text_out_reg_31_ ( .D(N400), .CK(clk), .Q(text_out[31]) );
WDDLDFFMS text_out_reg_30_ ( .D(N401), .CK(clk), .Q(text_out[30]) );
WDDLDFFMS text_out_reg_29_ ( .D(N402), .CK(clk), .Q(text_out[29]) );
WDDLDFFMS text_out_reg_28_ ( .D(N403), .CK(clk), .Q(text_out[28]) );
WDDLDFFMS text_out_reg_27_ ( .D(N404), .CK(clk), .Q(text_out[27]) );
WDDLDFFMS text_out_reg_26_ ( .D(N405), .CK(clk), .Q(text_out[26]) );
WDDLDFFMS text_out_reg_25_ ( .D(N406), .CK(clk), .Q(text_out[25]) );
WDDLDFFMS text_out_reg_24_ ( .D(N407), .CK(clk), .Q(text_out[24]) );
WDDLDFFMS text_out_reg_119_ ( .D(N408), .CK(clk), .Q(text_out[119]) );
WDDLDFFMS text_out_reg_118_ ( .D(N409), .CK(clk), .Q(text_out[118]) );
WDDLDFFMS text_out_reg_117_ ( .D(N410), .CK(clk), .Q(text_out[117]) );
WDDLDFFMS text_out_reg_116_ ( .D(N411), .CK(clk), .Q(text_out[116]) );
WDDLDFFMS text_out_reg_115_ ( .D(N412), .CK(clk), .Q(text_out[115]) );
WDDLDFFMS text_out_reg_114_ ( .D(N413), .CK(clk), .Q(text_out[114]) );
WDDLDFFMS text_out_reg_113_ ( .D(N414), .CK(clk), .Q(text_out[113]) );
WDDLDFFMS text_out_reg_112_ ( .D(N415), .CK(clk), .Q(text_out[112]) );
WDDLDFFMS text_out_reg_87_ ( .D(N416), .CK(clk), .Q(text_out[87]) );
WDDLDFFMS text_out_reg_86_ ( .D(N417), .CK(clk), .Q(text_out[86]) );
WDDLDFFMS text_out_reg_85_ ( .D(N418), .CK(clk), .Q(text_out[85]) );
WDDLDFFMS text_out_reg_84_ ( .D(N419), .CK(clk), .Q(text_out[84]) );
WDDLDFFMS text_out_reg_83_ ( .D(N420), .CK(clk), .Q(text_out[83]) );
WDDLDFFMS text_out_reg_82_ ( .D(N421), .CK(clk), .Q(text_out[82]) );
WDDLDFFMS text_out_reg_81_ ( .D(N422), .CK(clk), .Q(text_out[81]) );
WDDLDFFMS text_out_reg_80_ ( .D(N423), .CK(clk), .Q(text_out[80]) );
WDDLDFFMS text_out_reg_55_ ( .D(N424), .CK(clk), .Q(text_out[55]) );
WDDLDFFMS text_out_reg_54_ ( .D(N425), .CK(clk), .Q(text_out[54]) );
WDDLDFFMS text_out_reg_53_ ( .D(N426), .CK(clk), .Q(text_out[53]) );
WDDLDFFMS text_out_reg_52_ ( .D(N427), .CK(clk), .Q(text_out[52]) );
WDDLDFFMS text_out_reg_51_ ( .D(N428), .CK(clk), .Q(text_out[51]) );
WDDLDFFMS text_out_reg_50_ ( .D(N429), .CK(clk), .Q(text_out[50]) );
WDDLDFFMS text_out_reg_49_ ( .D(N430), .CK(clk), .Q(text_out[49]) );
WDDLDFFMS text_out_reg_48_ ( .D(N431), .CK(clk), .Q(text_out[48]) );
WDDLDFFMS text_out_reg_23_ ( .D(N432), .CK(clk), .Q(text_out[23]) );
WDDLDFFMS text_out_reg_22_ ( .D(N433), .CK(clk), .Q(text_out[22]) );
WDDLDFFMS text_out_reg_21_ ( .D(N434), .CK(clk), .Q(text_out[21]) );
WDDLDFFMS text_out_reg_20_ ( .D(N435), .CK(clk), .Q(text_out[20]) );
WDDLDFFMS text_out_reg_19_ ( .D(N436), .CK(clk), .Q(text_out[19]) );
WDDLDFFMS text_out_reg_18_ ( .D(N437), .CK(clk), .Q(text_out[18]) );
WDDLDFFMS text_out_reg_17_ ( .D(N438), .CK(clk), .Q(text_out[17]) );
WDDLDFFMS text_out_reg_16_ ( .D(N439), .CK(clk), .Q(text_out[16]) );
WDDLDFFMS text_out_reg_111_ ( .D(N440), .CK(clk), .Q(text_out[111]) );
WDDLDFFMS text_out_reg_110_ ( .D(N441), .CK(clk), .Q(text_out[110]) );
WDDLDFFMS text_out_reg_109_ ( .D(N442), .CK(clk), .Q(text_out[109]) );
WDDLDFFMS text_out_reg_108_ ( .D(N443), .CK(clk), .Q(text_out[108]) );
WDDLDFFMS text_out_reg_107_ ( .D(N444), .CK(clk), .Q(text_out[107]) );
WDDLDFFMS text_out_reg_106_ ( .D(N445), .CK(clk), .Q(text_out[106]) );
WDDLDFFMS text_out_reg_105_ ( .D(N446), .CK(clk), .Q(text_out[105]) );
WDDLDFFMS text_out_reg_104_ ( .D(N447), .CK(clk), .Q(text_out[104]) );
WDDLDFFMS text_out_reg_79_ ( .D(N448), .CK(clk), .Q(text_out[79]) );
WDDLDFFMS text_out_reg_78_ ( .D(N449), .CK(clk), .Q(text_out[78]) );
WDDLDFFMS text_out_reg_77_ ( .D(N450), .CK(clk), .Q(text_out[77]) );
WDDLDFFMS text_out_reg_76_ ( .D(N451), .CK(clk), .Q(text_out[76]) );
WDDLDFFMS text_out_reg_75_ ( .D(N452), .CK(clk), .Q(text_out[75]) );
WDDLDFFMS text_out_reg_74_ ( .D(N453), .CK(clk), .Q(text_out[74]) );
WDDLDFFMS text_out_reg_73_ ( .D(N454), .CK(clk), .Q(text_out[73]) );
WDDLDFFMS text_out_reg_72_ ( .D(N455), .CK(clk), .Q(text_out[72]) );
WDDLDFFMS text_out_reg_47_ ( .D(N456), .CK(clk), .Q(text_out[47]) );
WDDLDFFMS text_out_reg_46_ ( .D(N457), .CK(clk), .Q(text_out[46]) );
WDDLDFFMS text_out_reg_45_ ( .D(N458), .CK(clk), .Q(text_out[45]) );
WDDLDFFMS text_out_reg_44_ ( .D(N459), .CK(clk), .Q(text_out[44]) );
WDDLDFFMS text_out_reg_43_ ( .D(N460), .CK(clk), .Q(text_out[43]) );
WDDLDFFMS text_out_reg_42_ ( .D(N461), .CK(clk), .Q(text_out[42]) );
WDDLDFFMS text_out_reg_41_ ( .D(N462), .CK(clk), .Q(text_out[41]) );
WDDLDFFMS text_out_reg_40_ ( .D(N463), .CK(clk), .Q(text_out[40]) );
WDDLDFFMS text_out_reg_15_ ( .D(N464), .CK(clk), .Q(text_out[15]) );
WDDLDFFMS text_out_reg_14_ ( .D(N465), .CK(clk), .Q(text_out[14]) );
WDDLDFFMS text_out_reg_13_ ( .D(N466), .CK(clk), .Q(text_out[13]) );
WDDLDFFMS text_out_reg_12_ ( .D(N467), .CK(clk), .Q(text_out[12]) );
WDDLDFFMS text_out_reg_11_ ( .D(N468), .CK(clk), .Q(text_out[11]) );
WDDLDFFMS text_out_reg_10_ ( .D(N469), .CK(clk), .Q(text_out[10]) );
WDDLDFFMS text_out_reg_9_ ( .D(N470), .CK(clk), .Q(text_out[9]) );
WDDLDFFMS text_out_reg_8_ ( .D(N471), .CK(clk), .Q(text_out[8]) );
WDDLDFFMS text_out_reg_103_ ( .D(N472), .CK(clk), .Q(text_out[103]) );
WDDLDFFMS text_out_reg_102_ ( .D(N473), .CK(clk), .Q(text_out[102]) );
WDDLDFFMS text_out_reg_101_ ( .D(N474), .CK(clk), .Q(text_out[101]) );
WDDLDFFMS text_out_reg_100_ ( .D(N475), .CK(clk), .Q(text_out[100]) );
WDDLDFFMS text_out_reg_99_ ( .D(N476), .CK(clk), .Q(text_out[99]) );
WDDLDFFMS text_out_reg_98_ ( .D(N477), .CK(clk), .Q(text_out[98]) );
WDDLDFFMS text_out_reg_97_ ( .D(N478), .CK(clk), .Q(text_out[97]) );
WDDLDFFMS text_out_reg_96_ ( .D(N479), .CK(clk), .Q(text_out[96]) );
WDDLDFFMS text_out_reg_71_ ( .D(N480), .CK(clk), .Q(text_out[71]) );
WDDLDFFMS text_out_reg_70_ ( .D(N481), .CK(clk), .Q(text_out[70]) );
WDDLDFFMS text_out_reg_69_ ( .D(N482), .CK(clk), .Q(text_out[69]) );
WDDLDFFMS text_out_reg_68_ ( .D(N483), .CK(clk), .Q(text_out[68]) );
WDDLDFFMS text_out_reg_67_ ( .D(N484), .CK(clk), .Q(text_out[67]) );
WDDLDFFMS text_out_reg_66_ ( .D(N485), .CK(clk), .Q(text_out[66]) );
WDDLDFFMS text_out_reg_65_ ( .D(N486), .CK(clk), .Q(text_out[65]) );
WDDLDFFMS text_out_reg_64_ ( .D(N487), .CK(clk), .Q(text_out[64]) );
WDDLDFFMS text_out_reg_39_ ( .D(N488), .CK(clk), .Q(text_out[39]) );
WDDLDFFMS text_out_reg_38_ ( .D(N489), .CK(clk), .Q(text_out[38]) );
WDDLDFFMS text_out_reg_37_ ( .D(N490), .CK(clk), .Q(text_out[37]) );
WDDLDFFMS text_out_reg_36_ ( .D(N491), .CK(clk), .Q(text_out[36]) );
WDDLDFFMS text_out_reg_35_ ( .D(N492), .CK(clk), .Q(text_out[35]) );
WDDLDFFMS text_out_reg_34_ ( .D(N493), .CK(clk), .Q(text_out[34]) );
WDDLDFFMS text_out_reg_33_ ( .D(N494), .CK(clk), .Q(text_out[33]) );
WDDLDFFMS text_out_reg_32_ ( .D(N495), .CK(clk), .Q(text_out[32]) );
WDDLDFFMS text_out_reg_7_ ( .D(N496), .CK(clk), .Q(text_out[7]) );
WDDLDFFMS text_out_reg_6_ ( .D(N497), .CK(clk), .Q(text_out[6]) );
WDDLDFFMS text_out_reg_5_ ( .D(N498), .CK(clk), .Q(text_out[5]) );
WDDLDFFMS text_out_reg_4_ ( .D(N499), .CK(clk), .Q(text_out[4]) );
WDDLDFFMS text_out_reg_3_ ( .D(N500), .CK(clk), .Q(text_out[3]) );
WDDLDFFMS text_out_reg_2_ ( .D(N501), .CK(clk), .Q(text_out[2]) );
WDDLDFFMS text_out_reg_1_ ( .D(N502), .CK(clk), .Q(text_out[1]) );
WDDLDFFMS text_out_reg_0_ ( .D(N503), .CK(clk), .Q(text_out[0]) );
  EDFFX1 text_in_r_reg_127_ ( .D(text_in[127]), .E(ld), .CK(divclk), .Q(
        text_in_r[127]) );
  EDFFX1 text_in_r_reg_126_ ( .D(text_in[126]), .E(ld), .CK(divclk), .Q(
        text_in_r[126]) );
  EDFFX1 text_in_r_reg_125_ ( .D(text_in[125]), .E(ld), .CK(divclk), .Q(
        text_in_r[125]) );
  EDFFX1 text_in_r_reg_124_ ( .D(text_in[124]), .E(ld), .CK(divclk), .Q(
        text_in_r[124]) );
  EDFFX1 text_in_r_reg_123_ ( .D(text_in[123]), .E(ld), .CK(divclk), .Q(
        text_in_r[123]) );
  EDFFX1 text_in_r_reg_122_ ( .D(text_in[122]), .E(ld), .CK(divclk), .Q(
        text_in_r[122]) );
  EDFFX1 text_in_r_reg_121_ ( .D(text_in[121]), .E(ld), .CK(divclk), .Q(
        text_in_r[121]) );
  EDFFX1 text_in_r_reg_120_ ( .D(text_in[120]), .E(ld), .CK(divclk), .Q(
        text_in_r[120]) );
  EDFFX1 text_in_r_reg_119_ ( .D(text_in[119]), .E(ld), .CK(divclk), .Q(
        text_in_r[119]) );
  EDFFX1 text_in_r_reg_118_ ( .D(text_in[118]), .E(ld), .CK(divclk), .Q(
        text_in_r[118]) );
  EDFFX1 text_in_r_reg_117_ ( .D(text_in[117]), .E(ld), .CK(divclk), .Q(
        text_in_r[117]) );
  EDFFX1 text_in_r_reg_116_ ( .D(text_in[116]), .E(ld), .CK(divclk), .Q(
        text_in_r[116]) );
  EDFFX1 text_in_r_reg_115_ ( .D(text_in[115]), .E(ld), .CK(divclk), .Q(
        text_in_r[115]) );
  EDFFX1 text_in_r_reg_114_ ( .D(text_in[114]), .E(ld), .CK(divclk), .Q(
        text_in_r[114]) );
  EDFFX1 text_in_r_reg_113_ ( .D(text_in[113]), .E(ld), .CK(divclk), .Q(
        text_in_r[113]) );
  EDFFX1 text_in_r_reg_112_ ( .D(text_in[112]), .E(ld), .CK(divclk), .Q(
        text_in_r[112]) );
  EDFFX1 text_in_r_reg_111_ ( .D(text_in[111]), .E(ld), .CK(divclk), .Q(
        text_in_r[111]) );
  EDFFX1 text_in_r_reg_110_ ( .D(text_in[110]), .E(ld), .CK(divclk), .Q(
        text_in_r[110]) );
  EDFFX1 text_in_r_reg_109_ ( .D(text_in[109]), .E(ld), .CK(divclk), .Q(
        text_in_r[109]) );
  EDFFX1 text_in_r_reg_108_ ( .D(text_in[108]), .E(ld), .CK(divclk), .Q(
        text_in_r[108]) );
  EDFFX1 text_in_r_reg_107_ ( .D(text_in[107]), .E(ld), .CK(divclk), .Q(
        text_in_r[107]) );
  EDFFX1 text_in_r_reg_106_ ( .D(text_in[106]), .E(ld), .CK(divclk), .Q(
        text_in_r[106]) );
  EDFFX1 text_in_r_reg_105_ ( .D(text_in[105]), .E(ld), .CK(divclk), .Q(
        text_in_r[105]) );
  EDFFX1 text_in_r_reg_104_ ( .D(text_in[104]), .E(ld), .CK(divclk), .Q(
        text_in_r[104]) );
  EDFFX1 text_in_r_reg_103_ ( .D(text_in[103]), .E(ld), .CK(divclk), .Q(
        text_in_r[103]) );
  EDFFX1 text_in_r_reg_102_ ( .D(text_in[102]), .E(ld), .CK(divclk), .Q(
        text_in_r[102]) );
  EDFFX1 text_in_r_reg_101_ ( .D(text_in[101]), .E(ld), .CK(divclk), .Q(
        text_in_r[101]) );
  EDFFX1 text_in_r_reg_100_ ( .D(text_in[100]), .E(ld), .CK(divclk), .Q(
        text_in_r[100]) );
  EDFFX1 text_in_r_reg_99_ ( .D(text_in[99]), .E(ld), .CK(divclk), .Q(
        text_in_r[99]) );
  EDFFX1 text_in_r_reg_98_ ( .D(text_in[98]), .E(ld), .CK(divclk), .Q(
        text_in_r[98]) );
  EDFFX1 text_in_r_reg_97_ ( .D(text_in[97]), .E(ld), .CK(divclk), .Q(
        text_in_r[97]) );
  EDFFX1 text_in_r_reg_96_ ( .D(text_in[96]), .E(ld), .CK(divclk), .Q(
        text_in_r[96]) );
  EDFFX1 text_in_r_reg_95_ ( .D(text_in[95]), .E(ld), .CK(divclk), .Q(
        text_in_r[95]) );
  EDFFX1 text_in_r_reg_94_ ( .D(text_in[94]), .E(ld), .CK(divclk), .Q(
        text_in_r[94]) );
  EDFFX1 text_in_r_reg_93_ ( .D(text_in[93]), .E(ld), .CK(divclk), .Q(
        text_in_r[93]) );
  EDFFX1 text_in_r_reg_92_ ( .D(text_in[92]), .E(ld), .CK(divclk), .Q(
        text_in_r[92]) );
  EDFFX1 text_in_r_reg_91_ ( .D(text_in[91]), .E(ld), .CK(divclk), .Q(
        text_in_r[91]) );
  EDFFX1 text_in_r_reg_90_ ( .D(text_in[90]), .E(ld), .CK(divclk), .Q(
        text_in_r[90]) );
  EDFFX1 text_in_r_reg_89_ ( .D(text_in[89]), .E(ld), .CK(divclk), .Q(
        text_in_r[89]) );
  EDFFX1 text_in_r_reg_88_ ( .D(text_in[88]), .E(ld), .CK(divclk), .Q(
        text_in_r[88]) );
  EDFFX1 text_in_r_reg_87_ ( .D(text_in[87]), .E(ld), .CK(divclk), .Q(
        text_in_r[87]) );
  EDFFX1 text_in_r_reg_86_ ( .D(text_in[86]), .E(ld), .CK(divclk), .Q(
        text_in_r[86]) );
  EDFFX1 text_in_r_reg_85_ ( .D(text_in[85]), .E(ld), .CK(divclk), .Q(
        text_in_r[85]) );
  EDFFX1 text_in_r_reg_84_ ( .D(text_in[84]), .E(ld), .CK(divclk), .Q(
        text_in_r[84]) );
  EDFFX1 text_in_r_reg_83_ ( .D(text_in[83]), .E(ld), .CK(divclk), .Q(
        text_in_r[83]) );
  EDFFX1 text_in_r_reg_82_ ( .D(text_in[82]), .E(ld), .CK(divclk), .Q(
        text_in_r[82]) );
  EDFFX1 text_in_r_reg_81_ ( .D(text_in[81]), .E(ld), .CK(divclk), .Q(
        text_in_r[81]) );
  EDFFX1 text_in_r_reg_80_ ( .D(text_in[80]), .E(ld), .CK(divclk), .Q(
        text_in_r[80]) );
  EDFFX1 text_in_r_reg_79_ ( .D(text_in[79]), .E(ld), .CK(divclk), .Q(
        text_in_r[79]) );
  EDFFX1 text_in_r_reg_78_ ( .D(text_in[78]), .E(ld), .CK(divclk), .Q(
        text_in_r[78]) );
  EDFFX1 text_in_r_reg_77_ ( .D(text_in[77]), .E(ld), .CK(divclk), .Q(
        text_in_r[77]) );
  EDFFX1 text_in_r_reg_76_ ( .D(text_in[76]), .E(ld), .CK(divclk), .Q(
        text_in_r[76]) );
  EDFFX1 text_in_r_reg_75_ ( .D(text_in[75]), .E(ld), .CK(divclk), .Q(
        text_in_r[75]) );
  EDFFX1 text_in_r_reg_74_ ( .D(text_in[74]), .E(ld), .CK(divclk), .Q(
        text_in_r[74]) );
  EDFFX1 text_in_r_reg_73_ ( .D(text_in[73]), .E(ld), .CK(divclk), .Q(
        text_in_r[73]) );
  EDFFX1 text_in_r_reg_72_ ( .D(text_in[72]), .E(ld), .CK(divclk), .Q(
        text_in_r[72]) );
  EDFFX1 text_in_r_reg_71_ ( .D(text_in[71]), .E(ld), .CK(divclk), .Q(
        text_in_r[71]) );
  EDFFX1 text_in_r_reg_70_ ( .D(text_in[70]), .E(ld), .CK(divclk), .Q(
        text_in_r[70]) );
  EDFFX1 text_in_r_reg_69_ ( .D(text_in[69]), .E(ld), .CK(divclk), .Q(
        text_in_r[69]) );
  EDFFX1 text_in_r_reg_68_ ( .D(text_in[68]), .E(ld), .CK(divclk), .Q(
        text_in_r[68]) );
  EDFFX1 text_in_r_reg_67_ ( .D(text_in[67]), .E(ld), .CK(divclk), .Q(
        text_in_r[67]) );
  EDFFX1 text_in_r_reg_66_ ( .D(text_in[66]), .E(ld), .CK(divclk), .Q(
        text_in_r[66]) );
  EDFFX1 text_in_r_reg_65_ ( .D(text_in[65]), .E(ld), .CK(divclk), .Q(
        text_in_r[65]) );
  EDFFX1 text_in_r_reg_64_ ( .D(text_in[64]), .E(ld), .CK(divclk), .Q(
        text_in_r[64]) );
  EDFFX1 text_in_r_reg_63_ ( .D(text_in[63]), .E(ld), .CK(divclk), .Q(
        text_in_r[63]) );
  EDFFX1 text_in_r_reg_62_ ( .D(text_in[62]), .E(ld), .CK(divclk), .Q(
        text_in_r[62]) );
  EDFFX1 text_in_r_reg_61_ ( .D(text_in[61]), .E(ld), .CK(divclk), .Q(
        text_in_r[61]) );
  EDFFX1 text_in_r_reg_60_ ( .D(text_in[60]), .E(ld), .CK(divclk), .Q(
        text_in_r[60]) );
  EDFFX1 text_in_r_reg_59_ ( .D(text_in[59]), .E(ld), .CK(divclk), .Q(
        text_in_r[59]) );
  EDFFX1 text_in_r_reg_58_ ( .D(text_in[58]), .E(ld), .CK(divclk), .Q(
        text_in_r[58]) );
  EDFFX1 text_in_r_reg_57_ ( .D(text_in[57]), .E(ld), .CK(divclk), .Q(
        text_in_r[57]) );
  EDFFX1 text_in_r_reg_56_ ( .D(text_in[56]), .E(ld), .CK(divclk), .Q(
        text_in_r[56]) );
  EDFFX1 text_in_r_reg_55_ ( .D(text_in[55]), .E(ld), .CK(divclk), .Q(
        text_in_r[55]) );
  EDFFX1 text_in_r_reg_54_ ( .D(text_in[54]), .E(ld), .CK(divclk), .Q(
        text_in_r[54]) );
  EDFFX1 text_in_r_reg_53_ ( .D(text_in[53]), .E(ld), .CK(divclk), .Q(
        text_in_r[53]) );
  EDFFX1 text_in_r_reg_52_ ( .D(text_in[52]), .E(ld), .CK(divclk), .Q(
        text_in_r[52]) );
  EDFFX1 text_in_r_reg_51_ ( .D(text_in[51]), .E(ld), .CK(divclk), .Q(
        text_in_r[51]) );
  EDFFX1 text_in_r_reg_50_ ( .D(text_in[50]), .E(ld), .CK(divclk), .Q(
        text_in_r[50]) );
  EDFFX1 text_in_r_reg_49_ ( .D(text_in[49]), .E(ld), .CK(divclk), .Q(
        text_in_r[49]) );
  EDFFX1 text_in_r_reg_48_ ( .D(text_in[48]), .E(ld), .CK(divclk), .Q(
        text_in_r[48]) );
  EDFFX1 text_in_r_reg_47_ ( .D(text_in[47]), .E(ld), .CK(divclk), .Q(
        text_in_r[47]) );
  EDFFX1 text_in_r_reg_46_ ( .D(text_in[46]), .E(ld), .CK(divclk), .Q(
        text_in_r[46]) );
  EDFFX1 text_in_r_reg_45_ ( .D(text_in[45]), .E(ld), .CK(divclk), .Q(
        text_in_r[45]) );
  EDFFX1 text_in_r_reg_44_ ( .D(text_in[44]), .E(ld), .CK(divclk), .Q(
        text_in_r[44]) );
  EDFFX1 text_in_r_reg_43_ ( .D(text_in[43]), .E(ld), .CK(divclk), .Q(
        text_in_r[43]) );
  EDFFX1 text_in_r_reg_42_ ( .D(text_in[42]), .E(ld), .CK(divclk), .Q(
        text_in_r[42]) );
  EDFFX1 text_in_r_reg_41_ ( .D(text_in[41]), .E(ld), .CK(divclk), .Q(
        text_in_r[41]) );
  EDFFX1 text_in_r_reg_40_ ( .D(text_in[40]), .E(ld), .CK(divclk), .Q(
        text_in_r[40]) );
  EDFFX1 text_in_r_reg_39_ ( .D(text_in[39]), .E(ld), .CK(divclk), .Q(
        text_in_r[39]) );
  EDFFX1 text_in_r_reg_38_ ( .D(text_in[38]), .E(ld), .CK(divclk), .Q(
        text_in_r[38]) );
  EDFFX1 text_in_r_reg_37_ ( .D(text_in[37]), .E(ld), .CK(divclk), .Q(
        text_in_r[37]) );
  EDFFX1 text_in_r_reg_36_ ( .D(text_in[36]), .E(ld), .CK(divclk), .Q(
        text_in_r[36]) );
  EDFFX1 text_in_r_reg_7_ ( .D(text_in[7]), .E(ld), .CK(divclk), .Q(text_in_r[7])
         );
  EDFFX1 text_in_r_reg_6_ ( .D(text_in[6]), .E(ld), .CK(divclk), .Q(text_in_r[6])
         );
  EDFFX1 text_in_r_reg_5_ ( .D(text_in[5]), .E(ld), .CK(divclk), .Q(text_in_r[5])
         );
  EDFFX1 text_in_r_reg_4_ ( .D(text_in[4]), .E(ld), .CK(divclk), .Q(text_in_r[4])
         );
  EDFFX1 text_in_r_reg_3_ ( .D(text_in[3]), .E(ld), .CK(divclk), .Q(text_in_r[3])
         );
  EDFFX1 text_in_r_reg_2_ ( .D(text_in[2]), .E(ld), .CK(divclk), .Q(text_in_r[2])
         );
  EDFFX1 text_in_r_reg_1_ ( .D(text_in[1]), .E(ld), .CK(divclk), .Q(text_in_r[1])
         );
  EDFFX1 text_in_r_reg_0_ ( .D(text_in[0]), .E(ld), .CK(divclk), .Q(text_in_r[0])
         );
  EDFFX1 text_in_r_reg_35_ ( .D(text_in[35]), .E(ld), .CK(divclk), .Q(
        text_in_r[35]) );
  EDFFX1 text_in_r_reg_34_ ( .D(text_in[34]), .E(ld), .CK(divclk), .Q(
        text_in_r[34]) );
  EDFFX1 text_in_r_reg_33_ ( .D(text_in[33]), .E(ld), .CK(divclk), .Q(
        text_in_r[33]) );
  EDFFX1 text_in_r_reg_32_ ( .D(text_in[32]), .E(ld), .CK(divclk), .Q(
        text_in_r[32]) );
  EDFFX1 text_in_r_reg_31_ ( .D(text_in[31]), .E(ld), .CK(divclk), .Q(
        text_in_r[31]) );
  EDFFX1 text_in_r_reg_30_ ( .D(text_in[30]), .E(ld), .CK(divclk), .Q(
        text_in_r[30]) );
  EDFFX1 text_in_r_reg_29_ ( .D(text_in[29]), .E(ld), .CK(divclk), .Q(
        text_in_r[29]) );
  EDFFX1 text_in_r_reg_28_ ( .D(text_in[28]), .E(ld), .CK(divclk), .Q(
        text_in_r[28]) );
  EDFFX1 text_in_r_reg_27_ ( .D(text_in[27]), .E(ld), .CK(divclk), .Q(
        text_in_r[27]) );
  EDFFX1 text_in_r_reg_26_ ( .D(text_in[26]), .E(ld), .CK(divclk), .Q(
        text_in_r[26]) );
  EDFFX1 text_in_r_reg_25_ ( .D(text_in[25]), .E(ld), .CK(divclk), .Q(
        text_in_r[25]) );
  EDFFX1 text_in_r_reg_24_ ( .D(text_in[24]), .E(ld), .CK(divclk), .Q(
        text_in_r[24]) );
  EDFFX1 text_in_r_reg_23_ ( .D(text_in[23]), .E(ld), .CK(divclk), .Q(
        text_in_r[23]) );
  EDFFX1 text_in_r_reg_22_ ( .D(text_in[22]), .E(ld), .CK(divclk), .Q(
        text_in_r[22]) );
  EDFFX1 text_in_r_reg_21_ ( .D(text_in[21]), .E(ld), .CK(divclk), .Q(
        text_in_r[21]) );
  EDFFX1 text_in_r_reg_20_ ( .D(text_in[20]), .E(ld), .CK(divclk), .Q(
        text_in_r[20]) );
  EDFFX1 text_in_r_reg_19_ ( .D(text_in[19]), .E(ld), .CK(divclk), .Q(
        text_in_r[19]) );
  EDFFX1 text_in_r_reg_18_ ( .D(text_in[18]), .E(ld), .CK(divclk), .Q(
        text_in_r[18]) );
  EDFFX1 text_in_r_reg_17_ ( .D(text_in[17]), .E(ld), .CK(divclk), .Q(
        text_in_r[17]) );
  EDFFX1 text_in_r_reg_16_ ( .D(text_in[16]), .E(ld), .CK(divclk), .Q(
        text_in_r[16]) );
  EDFFX1 text_in_r_reg_15_ ( .D(text_in[15]), .E(ld), .CK(divclk), .Q(
        text_in_r[15]) );
  EDFFX1 text_in_r_reg_14_ ( .D(text_in[14]), .E(ld), .CK(divclk), .Q(
        text_in_r[14]) );
  EDFFX1 text_in_r_reg_13_ ( .D(text_in[13]), .E(ld), .CK(divclk), .Q(
        text_in_r[13]) );
  EDFFX1 text_in_r_reg_12_ ( .D(text_in[12]), .E(ld), .CK(divclk), .Q(
        text_in_r[12]) );
  EDFFX1 text_in_r_reg_11_ ( .D(text_in[11]), .E(ld), .CK(divclk), .Q(
        text_in_r[11]) );
  EDFFX1 text_in_r_reg_10_ ( .D(text_in[10]), .E(ld), .CK(divclk), .Q(
        text_in_r[10]) );
  EDFFX1 text_in_r_reg_9_ ( .D(text_in[9]), .E(ld), .CK(divclk), .Q(text_in_r[9])
         );
  EDFFX1 text_in_r_reg_8_ ( .D(text_in[8]), .E(ld), .CK(divclk), .Q(text_in_r[8])
         );
  DFFX1 dcnt_reg_1_ ( .D(n399), .CK(divclk), .QN(n3) );
  DFFHQX1 dcnt_reg_2_ ( .D(n398), .CK(divclk), .Q(dcnt_2_) );
WDDLDFFMS  sa21_reg_6_ ( .D(N182), .CK(clk), .Q(sa21[6]) );
WDDLDFFMS  sa11_reg_6_ ( .D(N198), .CK(clk), .Q(sa11[6]) );
WDDLDFFMS  sa01_reg_6_ ( .D(N214), .CK(clk), .Q(sa01[6]) );
WDDLDFFMS  sa12_reg_6_ ( .D(N134), .CK(clk), .Q(sa12[6]) );
WDDLDFFMS  sa02_reg_6_ ( .D(N150), .CK(clk), .Q(sa02[6]) );
WDDLDFFMS  sa22_reg_6_ ( .D(N118), .CK(clk), .Q(sa22[6]) );
WDDLDFFMS  sa13_reg_6_ ( .D(N70), .CK(clk), .Q(sa13[6]) );
WDDLDFFMS  sa03_reg_6_ ( .D(N86), .CK(clk), .Q(sa03[6]) );
WDDLDFFMS  sa23_reg_6_ ( .D(N54), .CK(clk), .Q(sa23[6]) );
WDDLDFFMS  sa10_reg_6_ ( .D(N262), .CK(clk), .Q(sa10[6]) );
WDDLDFFMS  sa00_reg_6_ ( .D(N278), .CK(clk), .Q(sa00[6]) );
WDDLDFFMS  sa20_reg_6_ ( .D(N246), .CK(clk), .Q(sa20[6]) );
WDDLDFFMS  sa00_reg_0_ ( .D(N272), .CK(clk), .Q(sa00[0]) );
WDDLDFFMS  sa22_reg_0_ ( .D(N112), .CK(clk), .Q(sa22[0]) );
WDDLDFFMS  sa21_reg_0_ ( .D(N176), .CK(clk), .Q(sa21[0]) );
WDDLDFFMS  sa23_reg_0_ ( .D(N48), .CK(clk), .Q(sa23[0]) );
WDDLDFFMS  sa31_reg_0_ ( .D(N160), .CK(clk), .Q(sa31[0]) );
WDDLDFFMS  sa01_reg_0_ ( .D(N208), .CK(clk), .Q(sa01[0]) );
WDDLDFFMS  sa02_reg_0_ ( .D(N144), .CK(clk), .Q(sa02[0]) );
WDDLDFFMS  sa32_reg_0_ ( .D(N96), .CK(clk), .Q(sa32[0]) );
WDDLDFFMS  sa03_reg_0_ ( .D(N80), .CK(clk), .Q(sa03[0]) );
WDDLDFFMS  sa33_reg_0_ ( .D(N32), .CK(clk), .Q(sa33[0]) );
WDDLDFFMS  sa30_reg_0_ ( .D(N224), .CK(clk), .Q(sa30[0]) );
WDDLDFFMS  sa11_reg_0_ ( .D(N192), .CK(clk), .Q(sa11[0]) );
WDDLDFFMS  sa13_reg_0_ ( .D(N64), .CK(clk), .Q(sa13[0]) );
WDDLDFFMS  sa20_reg_0_ ( .D(N240), .CK(clk), .Q(sa20[0]) );
WDDLDFFMS  sa12_reg_0_ ( .D(N128), .CK(clk), .Q(sa12[0]) );
WDDLDFFMS  sa10_reg_0_ ( .D(N256), .CK(clk), .Q(sa10[0]) );
WDDLDFFMS  sa31_reg_6_ ( .D(N166), .CK(clk), .Q(sa31[6]) );
WDDLDFFMS  sa32_reg_6_ ( .D(N102), .CK(clk), .Q(sa32[6]) );
WDDLDFFMS  sa33_reg_6_ ( .D(N38), .CK(clk), .Q(sa33[6]) );
WDDLDFFMS  sa30_reg_6_ ( .D(N230), .CK(clk), .Q(sa30[6]) );
WDDLDFFMS  sa21_reg_5_ ( .D(N181), .CK(clk), .Q(sa21[5]) );
WDDLDFFMS  sa22_reg_5_ ( .D(N117), .CK(clk), .Q(sa22[5]) );
WDDLDFFMS  sa23_reg_5_ ( .D(N53), .CK(clk), .Q(sa23[5]) );
WDDLDFFMS  sa20_reg_5_ ( .D(N245), .CK(clk), .Q(sa20[5]) );
WDDLDFFMS  sa21_reg_2_ ( .D(N178), .CK(clk), .Q(sa21[2]) );
WDDLDFFMS  sa11_reg_2_ ( .D(N194), .CK(clk), .Q(sa11[2]) );
WDDLDFFMS  sa12_reg_2_ ( .D(N130), .CK(clk), .Q(sa12[2]) );
WDDLDFFMS  sa22_reg_2_ ( .D(N114), .CK(clk), .Q(sa22[2]) );
WDDLDFFMS  sa13_reg_2_ ( .D(N66), .CK(clk), .Q(sa13[2]) );
WDDLDFFMS  sa23_reg_2_ ( .D(N50), .CK(clk), .Q(sa23[2]) );
WDDLDFFMS  sa10_reg_2_ ( .D(N258), .CK(clk), .Q(sa10[2]) );
WDDLDFFMS  sa20_reg_2_ ( .D(N242), .CK(clk), .Q(sa20[2]) );
WDDLDFFMS  sa10_reg_7_ ( .D(N263), .CK(clk), .Q(sa10[7]) );
WDDLDFFMS  sa03_reg_7_ ( .D(N87), .CK(clk), .Q(sa03[7]) );
WDDLDFFMS  sa13_reg_7_ ( .D(N71), .CK(clk), .Q(sa13[7]) );
WDDLDFFMS  sa02_reg_7_ ( .D(N151), .CK(clk), .Q(sa02[7]) );
WDDLDFFMS  sa12_reg_7_ ( .D(N135), .CK(clk), .Q(sa12[7]) );
WDDLDFFMS  sa01_reg_7_ ( .D(N215), .CK(clk), .Q(sa01[7]) );
WDDLDFFMS  sa11_reg_7_ ( .D(N199), .CK(clk), .Q(sa11[7]) );
WDDLDFFMS  sa20_reg_7_ ( .D(N247), .CK(clk), .Q(sa20[7]) );
WDDLDFFMS  sa21_reg_7_ ( .D(N183), .CK(clk), .Q(sa21[7]) );
WDDLDFFMS  sa23_reg_7_ ( .D(N55), .CK(clk), .Q(sa23[7]) );
WDDLDFFMS  sa22_reg_7_ ( .D(N119), .CK(clk), .Q(sa22[7]) );
WDDLDFFMS  sa00_reg_7_ ( .D(N279), .CK(clk), .Q(sa00[7]) );
WDDLDFFMS  sa31_reg_5_ ( .D(N165), .CK(clk), .Q(sa31[5]) );
WDDLDFFMS  sa11_reg_5_ ( .D(N197), .CK(clk), .Q(sa11[5]) );
WDDLDFFMS  sa01_reg_5_ ( .D(N213), .CK(clk), .Q(sa01[5]) );
WDDLDFFMS  sa32_reg_5_ ( .D(N101), .CK(clk), .Q(sa32[5]) );
WDDLDFFMS  sa12_reg_5_ ( .D(N133), .CK(clk), .Q(sa12[5]) );
WDDLDFFMS  sa02_reg_5_ ( .D(N149), .CK(clk), .Q(sa02[5]) );
WDDLDFFMS  sa33_reg_5_ ( .D(N37), .CK(clk), .Q(sa33[5]) );
WDDLDFFMS  sa13_reg_5_ ( .D(N69), .CK(clk), .Q(sa13[5]) );
WDDLDFFMS  sa03_reg_5_ ( .D(N85), .CK(clk), .Q(sa03[5]) );
WDDLDFFMS  sa30_reg_5_ ( .D(N229), .CK(clk), .Q(sa30[5]) );
WDDLDFFMS  sa10_reg_5_ ( .D(N261), .CK(clk), .Q(sa10[5]) );
WDDLDFFMS  sa00_reg_5_ ( .D(N277), .CK(clk), .Q(sa00[5]) );
WDDLDFFMS  sa21_reg_4_ ( .D(N180), .CK(clk), .Q(sa21[4]) );
WDDLDFFMS  sa22_reg_4_ ( .D(N116), .CK(clk), .Q(sa22[4]) );
WDDLDFFMS  sa23_reg_4_ ( .D(N52), .CK(clk), .Q(sa23[4]) );
WDDLDFFMS  sa11_reg_4_ ( .D(N196), .CK(clk), .Q(sa11[4]) );
WDDLDFFMS  sa13_reg_4_ ( .D(N68), .CK(clk), .Q(sa13[4]) );
WDDLDFFMS  sa20_reg_4_ ( .D(N244), .CK(clk), .Q(sa20[4]) );
WDDLDFFMS  sa12_reg_4_ ( .D(N132), .CK(clk), .Q(sa12[4]) );
WDDLDFFMS  sa10_reg_4_ ( .D(N260), .CK(clk), .Q(sa10[4]) );
WDDLDFFMS  sa21_reg_3_ ( .D(N179), .CK(clk), .Q(sa21[3]) );
WDDLDFFMS  sa31_reg_3_ ( .D(N163), .CK(clk), .Q(sa31[3]) );
WDDLDFFMS  sa01_reg_3_ ( .D(N211), .CK(clk), .Q(sa01[3]) );
WDDLDFFMS  sa02_reg_3_ ( .D(N147), .CK(clk), .Q(sa02[3]) );
WDDLDFFMS  sa22_reg_3_ ( .D(N115), .CK(clk), .Q(sa22[3]) );
WDDLDFFMS  sa32_reg_3_ ( .D(N99), .CK(clk), .Q(sa32[3]) );
WDDLDFFMS  sa03_reg_3_ ( .D(N83), .CK(clk), .Q(sa03[3]) );
WDDLDFFMS  sa23_reg_3_ ( .D(N51), .CK(clk), .Q(sa23[3]) );
WDDLDFFMS  sa33_reg_3_ ( .D(N35), .CK(clk), .Q(sa33[3]) );
WDDLDFFMS  sa30_reg_3_ ( .D(N227), .CK(clk), .Q(sa30[3]) );
WDDLDFFMS  sa11_reg_3_ ( .D(N195), .CK(clk), .Q(sa11[3]) );
WDDLDFFMS  sa13_reg_3_ ( .D(N67), .CK(clk), .Q(sa13[3]) );
WDDLDFFMS  sa20_reg_3_ ( .D(N243), .CK(clk), .Q(sa20[3]) );
WDDLDFFMS  sa12_reg_3_ ( .D(N131), .CK(clk), .Q(sa12[3]) );
WDDLDFFMS  sa00_reg_3_ ( .D(N275), .CK(clk), .Q(sa00[3]) );
WDDLDFFMS  sa10_reg_3_ ( .D(N259), .CK(clk), .Q(sa10[3]) );
WDDLDFFMS  sa31_reg_2_ ( .D(N162), .CK(clk), .Q(sa31[2]) );
WDDLDFFMS  sa01_reg_2_ ( .D(N210), .CK(clk), .Q(sa01[2]) );
WDDLDFFMS  sa32_reg_2_ ( .D(N98), .CK(clk), .Q(sa32[2]) );
WDDLDFFMS  sa02_reg_2_ ( .D(N146), .CK(clk), .Q(sa02[2]) );
WDDLDFFMS  sa33_reg_2_ ( .D(N34), .CK(clk), .Q(sa33[2]) );
WDDLDFFMS  sa03_reg_2_ ( .D(N82), .CK(clk), .Q(sa03[2]) );
WDDLDFFMS  sa30_reg_2_ ( .D(N226), .CK(clk), .Q(sa30[2]) );
WDDLDFFMS  sa00_reg_2_ ( .D(N274), .CK(clk), .Q(sa00[2]) );
WDDLDFFMS  sa30_reg_7_ ( .D(N231), .CK(clk), .Q(sa30[7]) );
WDDLDFFMS  sa31_reg_7_ ( .D(N167), .CK(clk), .Q(sa31[7]) );
WDDLDFFMS  sa32_reg_7_ ( .D(N103), .CK(clk), .Q(sa32[7]) );
WDDLDFFMS  sa33_reg_7_ ( .D(N39), .CK(clk), .Q(sa33[7]) );
WDDLDFFMS  sa31_reg_4_ ( .D(N164), .CK(clk), .Q(sa31[4]) );
WDDLDFFMS  sa01_reg_4_ ( .D(N212), .CK(clk), .Q(sa01[4]) );
WDDLDFFMS  sa02_reg_4_ ( .D(N148), .CK(clk), .Q(sa02[4]) );
WDDLDFFMS  sa32_reg_4_ ( .D(N100), .CK(clk), .Q(sa32[4]) );
WDDLDFFMS  sa03_reg_4_ ( .D(N84), .CK(clk), .Q(sa03[4]) );
WDDLDFFMS  sa33_reg_4_ ( .D(N36), .CK(clk), .Q(sa33[4]) );
WDDLDFFMS  sa30_reg_4_ ( .D(N228), .CK(clk), .Q(sa30[4]) );
WDDLDFFMS  sa00_reg_4_ ( .D(N276), .CK(clk), .Q(sa00[4]) );
  XOR2XL U1091 ( .A(w3[28]), .B(sa13_sr[4]), .Y(n480) );
  XOR2XL U671 ( .A(w0[28]), .B(sa10_sr[4]), .Y(n750) );
  XOR2XL U811 ( .A(w1[28]), .B(sa11_sr[4]), .Y(n660) );
  XOR2XL U951 ( .A(w2[28]), .B(sa12_sr[4]), .Y(n570) );
  XOR2XL U1022 ( .A(w2[13]), .B(sa32_sr[5]), .Y(n522) );
  XOR2XL U1066 ( .A(sa02_sr[5]), .B(sa12_sr[5]), .Y(n784) );
  XOR2XL U1162 ( .A(w3[13]), .B(sa33_sr[5]), .Y(n432) );
  XOR2XL U1206 ( .A(sa03_sr[5]), .B(sa13_sr[5]), .Y(n766) );
  XOR2XL U1016 ( .A(w2[12]), .B(sa32_sr[4]), .Y(n525) );
  XOR2XL U736 ( .A(w0[12]), .B(sa30_sr[4]), .Y(n705) );
  XOR2XL U876 ( .A(w1[12]), .B(sa31_sr[4]), .Y(n615) );
  XOR2XL U1161 ( .A(sa23_sr[7]), .B(sa33_sr[7]), .Y(n764) );
  XOR2XL U1156 ( .A(w3[12]), .B(sa33_sr[4]), .Y(n435) );
  XOR2XL U986 ( .A(sa12_sr[7]), .B(sa22_sr[7]), .Y(n780) );
  XOR2XL U981 ( .A(w2[20]), .B(sa02_sr[4]), .Y(n548) );
  XOR2XL U982 ( .A(sa12_sr[3]), .B(sa22_sr[3]), .Y(n547) );
  XOR2XL U706 ( .A(sa10_sr[7]), .B(sa20_sr[7]), .Y(n816) );
  XOR2XL U701 ( .A(w0[20]), .B(sa00_sr[4]), .Y(n728) );
  XOR2XL U702 ( .A(sa10_sr[3]), .B(sa20_sr[3]), .Y(n727) );
  XOR2XL U846 ( .A(sa11_sr[7]), .B(sa21_sr[7]), .Y(n798) );
  XOR2XL U841 ( .A(w1[20]), .B(sa01_sr[4]), .Y(n638) );
  XOR2XL U842 ( .A(sa11_sr[3]), .B(sa21_sr[3]), .Y(n637) );
  XOR2XL U1126 ( .A(sa13_sr[7]), .B(sa23_sr[7]), .Y(n762) );
  XOR2XL U1121 ( .A(w3[20]), .B(sa03_sr[4]), .Y(n458) );
  XOR2XL U1122 ( .A(sa13_sr[3]), .B(sa23_sr[3]), .Y(n457) );
  XOR2XL U815 ( .A(w1[29]), .B(sa11_sr[5]), .Y(n657) );
  XOR2XL U889 ( .A(sa21_sr[5]), .B(sa31_sr[5]), .Y(n803) );
  XOR2XL U675 ( .A(w0[29]), .B(sa10_sr[5]), .Y(n747) );
  XOR2XL U749 ( .A(sa20_sr[5]), .B(sa30_sr[5]), .Y(n821) );
  XOR2XL U800 ( .A(w1[25]), .B(sa11_sr[1]), .Y(n668) );
  XOR2XL U940 ( .A(w2[25]), .B(sa12_sr[1]), .Y(n578) );
  XOR2XL U660 ( .A(w0[25]), .B(sa10_sr[1]), .Y(n758) );
  XOR2XL U1080 ( .A(w3[25]), .B(sa13_sr[1]), .Y(n488) );
  XOR2XL U727 ( .A(w0[10]), .B(sa30_sr[2]), .Y(n710) );
  XOR2XL U768 ( .A(sa00_sr[2]), .B(sa10_sr[2]), .Y(n826) );
  XOR2XL U1007 ( .A(w2[10]), .B(sa32_sr[2]), .Y(n530) );
  XOR2XL U1147 ( .A(w3[10]), .B(sa33_sr[2]), .Y(n440) );
  XOR2XL U804 ( .A(w1[26]), .B(sa11_sr[2]), .Y(n665) );
  XOR2XL U875 ( .A(sa21_sr[2]), .B(sa31_sr[2]), .Y(n809) );
  XOR2XL U1084 ( .A(w3[26]), .B(sa13_sr[2]), .Y(n485) );
  XOR2XL U944 ( .A(w2[26]), .B(sa12_sr[2]), .Y(n575) );
  XOR2XL U992 ( .A(sa12_sr[5]), .B(sa22_sr[5]), .Y(n540) );
  XOR2XL U1033 ( .A(sa22_sr[6]), .B(sa32_sr[6]), .Y(n783) );
  XOR2XL U991 ( .A(w2[22]), .B(sa02_sr[6]), .Y(n541) );
  XOR2XL U712 ( .A(sa10_sr[5]), .B(sa20_sr[5]), .Y(n720) );
  XOR2XL U711 ( .A(w0[22]), .B(sa00_sr[6]), .Y(n721) );
  XOR2XL U852 ( .A(sa11_sr[5]), .B(sa21_sr[5]), .Y(n630) );
  XOR2XL U893 ( .A(sa21_sr[6]), .B(sa31_sr[6]), .Y(n801) );
  XOR2XL U851 ( .A(w1[22]), .B(sa01_sr[6]), .Y(n631) );
  XOR2XL U862 ( .A(w1[9]), .B(sa31_sr[1]), .Y(n623) );
  XOR2XL U722 ( .A(w0[9]), .B(sa30_sr[1]), .Y(n713) );
  XOR2XL U1142 ( .A(w3[9]), .B(sa33_sr[1]), .Y(n443) );
  XOR2XL U1002 ( .A(w2[9]), .B(sa32_sr[1]), .Y(n533) );
  XOR2XL U1132 ( .A(sa13_sr[5]), .B(sa23_sr[5]), .Y(n450) );
  XOR2XL U1173 ( .A(sa23_sr[6]), .B(sa33_sr[6]), .Y(n765) );
  XOR2XL U1131 ( .A(w3[22]), .B(sa03_sr[6]), .Y(n451) );
  XOR2XL U921 ( .A(sa01_sr[7]), .B(sa31_sr[7]), .Y(n797) );
  XOR2XL U781 ( .A(sa00_sr[7]), .B(sa30_sr[7]), .Y(n815) );
  XOR2XL U775 ( .A(w0[4]), .B(sa00_sr[3]), .Y(n683) );
  XOR2XL U776 ( .A(sa20_sr[4]), .B(sa30_sr[3]), .Y(n682) );
  XOR2XL U1061 ( .A(sa02_sr[7]), .B(sa32_sr[7]), .Y(n779) );
  XOR2XL U1055 ( .A(w2[4]), .B(sa02_sr[3]), .Y(n503) );
  XOR2XL U1056 ( .A(sa22_sr[4]), .B(sa32_sr[3]), .Y(n502) );
  XOR2XL U1195 ( .A(w3[4]), .B(sa03_sr[3]), .Y(n413) );
  XOR2XL U1196 ( .A(sa23_sr[4]), .B(sa33_sr[3]), .Y(n412) );
  XOR2XL U958 ( .A(w2[30]), .B(sa12_sr[6]), .Y(n565) );
  XOR2XL U890 ( .A(w1[15]), .B(sa31_sr[7]), .Y(n608) );
  XOR2XL U1030 ( .A(w2[15]), .B(sa32_sr[7]), .Y(n518) );
  XOR2XL U750 ( .A(w0[15]), .B(sa30_sr[7]), .Y(n698) );
  XOR2XL U1170 ( .A(w3[15]), .B(sa33_sr[7]), .Y(n428) );
  XOR2XL U687 ( .A(w0[17]), .B(sa00_sr[1]), .Y(n739) );
  XOR2XL U827 ( .A(w1[17]), .B(sa01_sr[1]), .Y(n649) );
  XOR2XL U1107 ( .A(w3[17]), .B(sa03_sr[1]), .Y(n469) );
  XOR2XL U967 ( .A(w2[17]), .B(sa02_sr[1]), .Y(n559) );
  XOR2XL U899 ( .A(sa21_sr[1]), .B(sa31_sr[0]), .Y(n603) );
  XOR2XL U1179 ( .A(sa23_sr[1]), .B(sa33_sr[0]), .Y(n423) );
  XOR2XL U759 ( .A(sa20_sr[1]), .B(sa30_sr[0]), .Y(n693) );
  XOR2XL U1039 ( .A(sa22_sr[1]), .B(sa32_sr[0]), .Y(n513) );
  XOR2XL U1087 ( .A(w3[27]), .B(sa13_sr[3]), .Y(n483) );
  XOR2XL U807 ( .A(w1[27]), .B(sa11_sr[3]), .Y(n663) );
  XOR2XL U667 ( .A(w0[27]), .B(sa10_sr[3]), .Y(n753) );
  XOR2XL U947 ( .A(w2[27]), .B(sa12_sr[3]), .Y(n573) );
  XOR2XL U923 ( .A(sa21_sr[5]), .B(sa31_sr[4]), .Y(n588) );
  XOR2XL U922 ( .A(w1[5]), .B(sa01_sr[4]), .Y(n589) );
  XOR2XL U1203 ( .A(sa23_sr[5]), .B(sa33_sr[4]), .Y(n408) );
  XOR2XL U1202 ( .A(w3[5]), .B(sa03_sr[4]), .Y(n409) );
  XOR2XL U1063 ( .A(sa22_sr[5]), .B(sa32_sr[4]), .Y(n498) );
  XOR2XL U1062 ( .A(w2[5]), .B(sa02_sr[4]), .Y(n499) );
  XOR2XL U783 ( .A(sa20_sr[5]), .B(sa30_sr[4]), .Y(n678) );
  XOR2XL U782 ( .A(w0[5]), .B(sa00_sr[4]), .Y(n679) );
  XOR2XL U1208 ( .A(sa23_sr[6]), .B(sa33_sr[5]), .Y(n405) );
  XOR2XL U1211 ( .A(sa03_sr[6]), .B(sa13_sr[6]), .Y(n763) );
  XOR2XL U1207 ( .A(w3[6]), .B(sa03_sr[5]), .Y(n406) );
  XOR2XL U788 ( .A(sa20_sr[6]), .B(sa30_sr[5]), .Y(n675) );
  XOR2XL U791 ( .A(sa00_sr[6]), .B(sa10_sr[6]), .Y(n817) );
  XOR2XL U787 ( .A(w0[6]), .B(sa00_sr[5]), .Y(n676) );
  XOR2XL U746 ( .A(w0[14]), .B(sa30_sr[6]), .Y(n700) );
  XOR2XL U1026 ( .A(w2[14]), .B(sa32_sr[6]), .Y(n520) );
  XOR2XL U1068 ( .A(sa22_sr[6]), .B(sa32_sr[5]), .Y(n495) );
  XOR2XL U1067 ( .A(w2[6]), .B(sa02_sr[5]), .Y(n496) );
  XOR2XL U886 ( .A(w1[14]), .B(sa31_sr[6]), .Y(n610) );
  XOR2XL U931 ( .A(sa01_sr[6]), .B(sa11_sr[6]), .Y(n799) );
  XOR2XL U928 ( .A(sa21_sr[6]), .B(sa31_sr[5]), .Y(n585) );
  XOR2XL U927 ( .A(w1[6]), .B(sa01_sr[5]), .Y(n586) );
  XOR2XL U681 ( .A(w0[31]), .B(sa10_sr[7]), .Y(n743) );
  XOR2XL U961 ( .A(w2[31]), .B(sa12_sr[7]), .Y(n563) );
  XOR2XL U1101 ( .A(w3[31]), .B(sa13_sr[7]), .Y(n473) );
  XOR2XL U821 ( .A(w1[31]), .B(sa11_sr[7]), .Y(n653) );
  XOR2XL U1011 ( .A(w2[11]), .B(sa32_sr[3]), .Y(n528) );
  XOR2XL U871 ( .A(w1[11]), .B(sa31_sr[3]), .Y(n618) );
  XOR2XL U1166 ( .A(w3[14]), .B(sa33_sr[6]), .Y(n430) );
  XOR2XL U731 ( .A(w0[11]), .B(sa30_sr[3]), .Y(n708) );
  XOR2XL U1151 ( .A(w3[11]), .B(sa33_sr[3]), .Y(n438) );
  XOR2XL U856 ( .A(sa11_sr[6]), .B(sa21_sr[6]), .Y(n627) );
  XOR2XL U855 ( .A(w1[23]), .B(sa01_sr[7]), .Y(n628) );
  XOR2XL U1136 ( .A(sa13_sr[6]), .B(sa23_sr[6]), .Y(n447) );
  XOR2XL U1135 ( .A(w3[23]), .B(sa03_sr[7]), .Y(n448) );
  XOR2XL U996 ( .A(sa12_sr[6]), .B(sa22_sr[6]), .Y(n537) );
  XOR2XL U995 ( .A(w2[23]), .B(sa02_sr[7]), .Y(n538) );
  XOR2XL U1045 ( .A(sa22_sr[2]), .B(sa32_sr[1]), .Y(n509) );
  XOR2XL U1044 ( .A(w2[2]), .B(sa02_sr[1]), .Y(n510) );
  XOR2XL U905 ( .A(sa21_sr[2]), .B(sa31_sr[1]), .Y(n599) );
  XOR2XL U904 ( .A(w1[2]), .B(sa01_sr[1]), .Y(n600) );
  XOR2XL U1185 ( .A(sa23_sr[2]), .B(sa33_sr[1]), .Y(n419) );
  XOR2XL U1184 ( .A(w3[2]), .B(sa03_sr[1]), .Y(n420) );
  XOR2XL U765 ( .A(sa20_sr[2]), .B(sa30_sr[1]), .Y(n689) );
  XOR2XL U764 ( .A(w0[2]), .B(sa00_sr[1]), .Y(n690) );
  XOR2XL U716 ( .A(sa10_sr[6]), .B(sa20_sr[6]), .Y(n717) );
  XOR2XL U715 ( .A(w0[23]), .B(sa00_sr[7]), .Y(n718) );
  XOR2XL U696 ( .A(w0[19]), .B(sa00_sr[3]), .Y(n732) );
  XOR2XL U697 ( .A(sa10_sr[2]), .B(sa20_sr[2]), .Y(n731) );
  XOR2XL U836 ( .A(w1[19]), .B(sa01_sr[3]), .Y(n642) );
  XOR2XL U837 ( .A(sa11_sr[2]), .B(sa21_sr[2]), .Y(n641) );
  XOR2XL U976 ( .A(w2[19]), .B(sa02_sr[3]), .Y(n552) );
  XOR2XL U977 ( .A(sa12_sr[2]), .B(sa22_sr[2]), .Y(n551) );
  XOR2XL U1116 ( .A(w3[19]), .B(sa03_sr[3]), .Y(n462) );
  XOR2XL U1117 ( .A(sa13_sr[2]), .B(sa23_sr[2]), .Y(n461) );
  XOR2XL U988 ( .A(sa12_sr[4]), .B(sa22_sr[4]), .Y(n543) );
  XOR2XL U987 ( .A(w2[21]), .B(sa02_sr[5]), .Y(n544) );
  XOR2XL U708 ( .A(sa10_sr[4]), .B(sa20_sr[4]), .Y(n723) );
  XOR2XL U707 ( .A(w0[21]), .B(sa00_sr[5]), .Y(n724) );
  XOR2XL U848 ( .A(sa11_sr[4]), .B(sa21_sr[4]), .Y(n633) );
  XOR2XL U847 ( .A(w1[21]), .B(sa01_sr[5]), .Y(n634) );
  XOR2XL U1128 ( .A(sa13_sr[4]), .B(sa23_sr[4]), .Y(n453) );
  XOR2XL U1127 ( .A(w3[21]), .B(sa03_sr[5]), .Y(n454) );
  XOR2XL U909 ( .A(w1[3]), .B(sa01_sr[2]), .Y(n597) );
  XOR2XL U910 ( .A(sa21_sr[3]), .B(sa31_sr[2]), .Y(n596) );
  XOR2XL U1189 ( .A(w3[3]), .B(sa03_sr[2]), .Y(n417) );
  XOR2XL U1190 ( .A(sa23_sr[3]), .B(sa33_sr[2]), .Y(n416) );
  XOR2XL U1072 ( .A(w2[7]), .B(sa02_sr[6]), .Y(n493) );
  XOR2XL U793 ( .A(sa20_sr[7]), .B(sa30_sr[6]), .Y(n672) );
  XOR2XL U792 ( .A(w0[7]), .B(sa00_sr[6]), .Y(n673) );
  XOR2XL U932 ( .A(w1[7]), .B(sa01_sr[6]), .Y(n583) );
  XOR2XL U1212 ( .A(w3[7]), .B(sa03_sr[6]), .Y(n403) );
  XOR2XL U833 ( .A(sa11_sr[1]), .B(sa21_sr[1]), .Y(n644) );
  XOR2XL U832 ( .A(w1[18]), .B(sa01_sr[2]), .Y(n645) );
  XOR2XL U693 ( .A(sa10_sr[1]), .B(sa20_sr[1]), .Y(n734) );
  XOR2XL U692 ( .A(w0[18]), .B(sa00_sr[2]), .Y(n735) );
  XOR2XL U973 ( .A(sa12_sr[1]), .B(sa22_sr[1]), .Y(n554) );
  XOR2XL U972 ( .A(w2[18]), .B(sa02_sr[2]), .Y(n555) );
  XOR2XL U1113 ( .A(sa13_sr[1]), .B(sa23_sr[1]), .Y(n464) );
  XOR2XL U1112 ( .A(w3[18]), .B(sa03_sr[2]), .Y(n465) );
  DFFX4 ld_r_reg ( .D(ld), .CK(divclk), .Q(n960), .QN(n4) );
WDDLDFFMS sa32_reg_1_ ( .D(N97), .CK(clk), .Q(sa32[1]) );
WDDLDFFMS sa31_reg_1_ ( .D(N161), .CK(clk), .Q(sa31[1]) );
WDDLDFFMS sa30_reg_1_ ( .D(N225), .CK(clk), .Q(sa30[1]) );
WDDLDFFMS sa33_reg_1_ ( .D(N33), .CK(clk), .Q(sa33[1]) );
WDDLDFFMS sa21_reg_1_ ( .D(N177), .CK(clk), .Q(sa21[1]) );
WDDLDFFMS sa20_reg_1_ ( .D(N241), .CK(clk), .Q(sa20[1]) );
  //wddl
  //DFFHQX2 sa23_reg_1_ ( .D(N49), .CK(divclk), .Q(sa23[1]) );
WDDLDFFHQX2 sa23_reg_1_ ( .D(N49), .Dinv(N49inv), .CLK(clk), .PRECLK(divclk), .Q(sa23[1]));
//DFFHQX1 sa23_reg_1_ ( .D(N49), .CK(divclk), .Q(sa23[1]) );
//WDDLDFFMS sa23_reg_1_ ( .D(N49), .CK(clk), .Q(sa23[1]) );
WDDLDFFMS sa22_reg_1_ ( .D(N113), .CK(clk), .Q(sa22[1]) );
WDDLDFFMS sa10_reg_1_ ( .D(N257), .CK(clk), .Q(sa10[1]) );
WDDLDFFMS sa13_reg_1_ ( .D(N65), .CK(clk), .Q(sa13[1]) );
WDDLDFFMS sa12_reg_1_ ( .D(N129), .CK(clk), .Q(sa12[1]) );
WDDLDFFMS sa11_reg_1_ ( .D(N193), .CK(clk), .Q(sa11[1]) );
WDDLDFFMS sa03_reg_1_ ( .D(N81), .CK(clk), .Q(sa03[1]) );
WDDLDFFMS sa02_reg_1_ ( .D(N145), .CK(clk), .Q(sa02[1]) );
WDDLDFFMS sa01_reg_1_ ( .D(N209), .CK(clk), .Q(sa01[1]) );
WDDLDFFMS sa00_reg_1_ ( .D(N273), .CK(clk), .Q(sa00[1]) );
  XOR2X1 U898 ( .A(w1[1]), .B(sa01_sr[0]), .Y(n604) );
  XOR2X1 U684 ( .A(w0[16]), .B(sa00_sr[0]), .Y(n741) );
  XOR2X1 U866 ( .A(sa21_sr[0]), .B(sa31_sr[0]), .Y(n813) );
  XOR2X1 U719 ( .A(w0[8]), .B(sa30_sr[0]), .Y(n715) );
  XOR2X1 U897 ( .A(sa01_sr[0]), .B(sa11_sr[0]), .Y(n812) );
  XOR2X1 U1177 ( .A(sa03_sr[0]), .B(sa13_sr[0]), .Y(n776) );
  XOR2X1 U1038 ( .A(w2[1]), .B(sa02_sr[0]), .Y(n514) );
  XOR2X1 U754 ( .A(w0[0]), .B(sa20_sr[0]), .Y(n696) );
  XOR2X1 U758 ( .A(w0[1]), .B(sa00_sr[0]), .Y(n694) );
  XOR2X1 U1037 ( .A(sa02_sr[0]), .B(sa12_sr[0]), .Y(n794) );
  XOR2X1 U1077 ( .A(w3[24]), .B(sa13_sr[0]), .Y(n490) );
  XOR2X1 U657 ( .A(w0[24]), .B(sa10_sr[0]), .Y(n760) );
  XOR2X1 U1146 ( .A(sa23_sr[0]), .B(sa33_sr[0]), .Y(n777) );
  XOR2X1 U726 ( .A(sa20_sr[0]), .B(sa30_sr[0]), .Y(n831) );
  XOR2X1 U1006 ( .A(sa22_sr[0]), .B(sa32_sr[0]), .Y(n795) );
  XOR2X1 U1178 ( .A(w3[1]), .B(sa03_sr[0]), .Y(n424) );
  XOR2X1 U757 ( .A(sa00_sr[0]), .B(sa10_sr[0]), .Y(n830) );
  XOR2X1 U1174 ( .A(w3[0]), .B(sa23_sr[0]), .Y(n426) );
  XOR2X1 U1139 ( .A(w3[8]), .B(sa33_sr[0]), .Y(n445) );
  XOR2X1 U1021 ( .A(sa22_sr[7]), .B(sa32_sr[7]), .Y(n782) );
  XOR2X1 U1025 ( .A(sa22_sr[4]), .B(sa32_sr[4]), .Y(n787) );
  XOR2X1 U1015 ( .A(sa22_sr[2]), .B(sa32_sr[2]), .Y(n791) );
  XOR2X1 U1048 ( .A(sa02_sr[2]), .B(sa12_sr[2]), .Y(n790) );
  XOR2X1 U1194 ( .A(sa03_sr[3]), .B(sa13_sr[3]), .Y(n770) );
  XOR2X1 U741 ( .A(sa20_sr[7]), .B(sa30_sr[7]), .Y(n818) );
  XOR2X1 U1201 ( .A(sa03_sr[7]), .B(sa33_sr[7]), .Y(n761) );
  XOR2X1 U1020 ( .A(sa22_sr[3]), .B(sa32_sr[3]), .Y(n789) );
  XOR2X1 U753 ( .A(sa20_sr[6]), .B(sa30_sr[6]), .Y(n819) );
  XOR2X1 U735 ( .A(sa20_sr[2]), .B(sa30_sr[2]), .Y(n827) );
  XOR2X1 U1160 ( .A(sa23_sr[3]), .B(sa33_sr[3]), .Y(n771) );
  XOR2X1 U786 ( .A(sa00_sr[5]), .B(sa10_sr[5]), .Y(n820) );
  XOR2X1 U1188 ( .A(sa03_sr[2]), .B(sa13_sr[2]), .Y(n772) );
  XOR2X1 U867 ( .A(w1[10]), .B(sa31_sr[2]), .Y(n620) );
  XOR2X1 U1060 ( .A(sa02_sr[4]), .B(sa12_sr[4]), .Y(n786) );
  XOR2X1 U1054 ( .A(sa02_sr[3]), .B(sa12_sr[3]), .Y(n788) );
  XOR2X1 U955 ( .A(w2[29]), .B(sa12_sr[5]), .Y(n567) );
  XOR2X1 U1071 ( .A(sa02_sr[6]), .B(sa12_sr[6]), .Y(n781) );
  XOR2X1 U1169 ( .A(sa23_sr[5]), .B(sa33_sr[5]), .Y(n767) );
  XOR2X1 U1029 ( .A(sa22_sr[5]), .B(sa32_sr[5]), .Y(n785) );
  XOR2X1 U1155 ( .A(sa23_sr[2]), .B(sa33_sr[2]), .Y(n773) );
  XOR2X1 U920 ( .A(sa01_sr[4]), .B(sa11_sr[4]), .Y(n804) );
  XOR2X1 U745 ( .A(sa20_sr[4]), .B(sa30_sr[4]), .Y(n823) );
  XOR2X1 U926 ( .A(sa01_sr[5]), .B(sa11_sr[5]), .Y(n802) );
  XOR2X1 U908 ( .A(sa01_sr[2]), .B(sa11_sr[2]), .Y(n808) );
  XOR2X1 U1076 ( .A(sa02_sr[7]), .B(sa12_sr[7]), .Y(n796) );
  XOR2X1 U1200 ( .A(sa03_sr[4]), .B(sa13_sr[4]), .Y(n768) );
  XOR2X1 U740 ( .A(sa20_sr[3]), .B(sa30_sr[3]), .Y(n825) );
  XOR2X1 U1216 ( .A(sa03_sr[7]), .B(sa13_sr[7]), .Y(n778) );
  XOR2X1 U880 ( .A(sa21_sr[3]), .B(sa31_sr[3]), .Y(n807) );
  XOR2X1 U774 ( .A(sa00_sr[3]), .B(sa10_sr[3]), .Y(n824) );
  XOR2X1 U881 ( .A(sa21_sr[7]), .B(sa31_sr[7]), .Y(n800) );
  XOR2X1 U796 ( .A(sa00_sr[7]), .B(sa10_sr[7]), .Y(n832) );
  XOR2X1 U936 ( .A(sa01_sr[7]), .B(sa11_sr[7]), .Y(n814) );
  XOR2X1 U914 ( .A(sa01_sr[3]), .B(sa11_sr[3]), .Y(n806) );
  XOR2X1 U1165 ( .A(sa23_sr[4]), .B(sa33_sr[4]), .Y(n769) );
  XOR2X1 U780 ( .A(sa00_sr[4]), .B(sa10_sr[4]), .Y(n822) );
  XOR2X1 U885 ( .A(sa21_sr[4]), .B(sa31_sr[4]), .Y(n805) );
  XOR2X1 U703 ( .A(n816), .B(n823), .Y(n726) );
  XOR2X1 U738 ( .A(n825), .B(n705), .Y(n703) );
  XOR2X1 U956 ( .A(n786), .B(n785), .Y(n566) );
  XOR2X1 U1140 ( .A(n764), .B(n776), .Y(n444) );
  XOR2X1 U1064 ( .A(n784), .B(n499), .Y(n497) );
  XOR2X1 U1089 ( .A(n771), .B(n483), .Y(n481) );
  XOR2X1 U1058 ( .A(n503), .B(n502), .Y(n500) );
  XOR2X1 U979 ( .A(n552), .B(n551), .Y(n549) );
  XOR2X1 U1133 ( .A(n765), .B(n451), .Y(n449) );
  XOR2X1 U1092 ( .A(n778), .B(n770), .Y(n479) );
  XOR2X1 U747 ( .A(n817), .B(n821), .Y(n699) );
  XOR2X1 U1175 ( .A(n761), .B(n776), .Y(n425) );
  XOR2X1 U1123 ( .A(n762), .B(n769), .Y(n456) );
  XOR2X1 U658 ( .A(n832), .B(n831), .Y(n759) );
  XOR2X1 U1057 ( .A(n779), .B(n786), .Y(n501) );
  XOR2X1 U997 ( .A(n782), .B(n538), .Y(n536) );
  XOR2X1 U1010 ( .A(sa22_sr[1]), .B(sa32_sr[1]), .Y(n793) );
  XOR2X1 U993 ( .A(n783), .B(n541), .Y(n539) );
  XOR2X1 U717 ( .A(n818), .B(n718), .Y(n716) );
  XOR2X1 U699 ( .A(n732), .B(n731), .Y(n729) );
  XOR2X1 U730 ( .A(sa20_sr[1]), .B(sa30_sr[1]), .Y(n829) );
  XOR2X1 U1191 ( .A(n761), .B(n770), .Y(n415) );
  XOR2X1 U704 ( .A(n728), .B(n727), .Y(n725) );
  XOR2X1 U989 ( .A(n785), .B(n544), .Y(n542) );
  XOR2X1 U1192 ( .A(n417), .B(n416), .Y(n414) );
  XOR2X1 U713 ( .A(n819), .B(n721), .Y(n719) );
  XOR2X1 U983 ( .A(n780), .B(n787), .Y(n546) );
  XOR2X1 U751 ( .A(n832), .B(n819), .Y(n697) );
  XOR2X1 U1114 ( .A(n773), .B(n465), .Y(n463) );
  XOR2X1 U1129 ( .A(n767), .B(n454), .Y(n452) );
  XOR2X1 U673 ( .A(n823), .B(n750), .Y(n748) );
  XOR2X1 U698 ( .A(n816), .B(n825), .Y(n730) );
  XOR2X1 U1078 ( .A(n778), .B(n777), .Y(n489) );
  XOR2X1 U1137 ( .A(n764), .B(n448), .Y(n446) );
  XOR2X1 U1209 ( .A(n763), .B(n406), .Y(n404) );
  XOR2X1 U1183 ( .A(sa03_sr[1]), .B(sa13_sr[1]), .Y(n774) );
  XOR2X1 U676 ( .A(n822), .B(n821), .Y(n746) );
  XOR2X1 U709 ( .A(n821), .B(n724), .Y(n722) );
  XOR2X1 U1214 ( .A(n778), .B(n403), .Y(n401) );
  XOR2X1 U682 ( .A(n818), .B(n817), .Y(n742) );
  XOR2X1 U984 ( .A(n548), .B(n547), .Y(n545) );
  XOR2X1 U1118 ( .A(n762), .B(n771), .Y(n460) );
  XOR2X1 U685 ( .A(n816), .B(n831), .Y(n740) );
  XOR2X1 U948 ( .A(n796), .B(n790), .Y(n572) );
  XOR2X1 U1197 ( .A(n761), .B(n768), .Y(n411) );
  XOR2X1 U763 ( .A(sa00_sr[1]), .B(sa10_sr[1]), .Y(n828) );
  XOR2X1 U949 ( .A(n789), .B(n573), .Y(n571) );
  XOR2X1 U959 ( .A(n784), .B(n783), .Y(n564) );
  XOR2X1 U952 ( .A(n796), .B(n788), .Y(n569) );
  XOR2X1 U1124 ( .A(n458), .B(n457), .Y(n455) );
  XOR2X1 U1198 ( .A(n413), .B(n412), .Y(n410) );
  XOR2X1 U1119 ( .A(n462), .B(n461), .Y(n459) );
  XOR2X1 U953 ( .A(n787), .B(n570), .Y(n568) );
  XOR2X1 U1069 ( .A(n781), .B(n496), .Y(n494) );
  XOR2X1 U668 ( .A(n832), .B(n826), .Y(n752) );
  XOR2X1 U962 ( .A(n782), .B(n781), .Y(n562) );
  XOR2X1 U694 ( .A(n827), .B(n735), .Y(n733) );
  XOR2X1 U1204 ( .A(n766), .B(n409), .Y(n407) );
  XOR2X1 U669 ( .A(n825), .B(n753), .Y(n751) );
  XOR2X1 U672 ( .A(n832), .B(n824), .Y(n749) );
  XOR2X1 U903 ( .A(sa01_sr[1]), .B(sa11_sr[1]), .Y(n810) );
  XOR2X1 U808 ( .A(n814), .B(n808), .Y(n662) );
  XOR2X1 U1074 ( .A(n796), .B(n493), .Y(n491) );
  XOR2X1 U870 ( .A(sa21_sr[1]), .B(sa31_sr[1]), .Y(n811) );
  XOR2X1 U801 ( .A(n814), .B(n812), .Y(n667) );
  XOR2X1 U809 ( .A(n807), .B(n663), .Y(n661) );
  XOR2X1 U1093 ( .A(n769), .B(n480), .Y(n478) );
  XOR2X1 U812 ( .A(n814), .B(n806), .Y(n659) );
  XOR2X1 U813 ( .A(n805), .B(n660), .Y(n658) );
  XOR2X1 U816 ( .A(n804), .B(n803), .Y(n656) );
  XOR2X1 U934 ( .A(n814), .B(n583), .Y(n581) );
  XOR2X1 U822 ( .A(n800), .B(n799), .Y(n652) );
  XOR2X1 U1088 ( .A(n778), .B(n772), .Y(n482) );
  XOR2X1 U857 ( .A(n800), .B(n628), .Y(n626) );
  XOR2X1 U872 ( .A(n800), .B(n806), .Y(n617) );
  XOR2X1 U755 ( .A(n815), .B(n830), .Y(n695) );
  XOR2X1 U873 ( .A(n809), .B(n618), .Y(n616) );
  XOR2X1 U1043 ( .A(sa02_sr[1]), .B(sa12_sr[1]), .Y(n792) );
  XOR2X1 U853 ( .A(n801), .B(n631), .Y(n629) );
  XOR2X1 U1012 ( .A(n782), .B(n788), .Y(n527) );
  XOR2X1 U929 ( .A(n799), .B(n586), .Y(n584) );
  XOR2X1 U1013 ( .A(n791), .B(n528), .Y(n526) );
  XOR2X1 U1152 ( .A(n764), .B(n770), .Y(n437) );
  XOR2X1 U877 ( .A(n800), .B(n804), .Y(n614) );
  XOR2X1 U1153 ( .A(n773), .B(n438), .Y(n436) );
  XOR2X1 U878 ( .A(n807), .B(n615), .Y(n613) );
  XOR2X1 U849 ( .A(n803), .B(n634), .Y(n632) );
  XOR2X1 U777 ( .A(n815), .B(n822), .Y(n681) );
  XOR2X1 U924 ( .A(n802), .B(n589), .Y(n587) );
  XOR2X1 U778 ( .A(n683), .B(n682), .Y(n680) );
  XOR2X1 U1150 ( .A(sa23_sr[1]), .B(sa33_sr[1]), .Y(n775) );
  XOR2X1 U1157 ( .A(n764), .B(n768), .Y(n434) );
  XOR2X1 U1017 ( .A(n782), .B(n786), .Y(n524) );
  XOR2X1 U1158 ( .A(n771), .B(n435), .Y(n433) );
  XOR2X1 U1018 ( .A(n789), .B(n525), .Y(n523) );
  XOR2X1 U844 ( .A(n638), .B(n637), .Y(n635) );
  XOR2X1 U784 ( .A(n820), .B(n679), .Y(n677) );
  XOR2X1 U887 ( .A(n799), .B(n803), .Y(n609) );
  XOR2X1 U1163 ( .A(n766), .B(n769), .Y(n431) );
  XOR2X1 U1023 ( .A(n784), .B(n787), .Y(n521) );
  XOR2X1 U789 ( .A(n817), .B(n676), .Y(n674) );
  XOR2X1 U1031 ( .A(n796), .B(n783), .Y(n517) );
  XOR2X1 U891 ( .A(n814), .B(n801), .Y(n607) );
  XOR2X1 U1027 ( .A(n781), .B(n785), .Y(n519) );
  XOR2X1 U794 ( .A(n832), .B(n673), .Y(n671) );
  XOR2X1 U1171 ( .A(n778), .B(n765), .Y(n427) );
  XOR2X1 U737 ( .A(n818), .B(n822), .Y(n704) );
  XOR2X1 U839 ( .A(n642), .B(n641), .Y(n639) );
  XOR2X1 U838 ( .A(n798), .B(n807), .Y(n640) );
  XOR2X1 U733 ( .A(n827), .B(n708), .Y(n706) );
  XOR2X1 U843 ( .A(n798), .B(n805), .Y(n636) );
  XOR2X1 U834 ( .A(n809), .B(n645), .Y(n643) );
  XOR2X1 U978 ( .A(n780), .B(n789), .Y(n550) );
  XOR2X1 U974 ( .A(n791), .B(n555), .Y(n553) );
  XOR2X1 U720 ( .A(n818), .B(n830), .Y(n714) );
  XOR2X1 U1081 ( .A(n778), .B(n776), .Y(n487) );
  XOR2X1 U912 ( .A(n597), .B(n596), .Y(n594) );
  XOR2X1 U911 ( .A(n797), .B(n806), .Y(n595) );
  XOR2X1 U732 ( .A(n818), .B(n824), .Y(n707) );
  XOR2X1 U1167 ( .A(n763), .B(n767), .Y(n429) );
  XOR2X1 U1075 ( .A(n492), .B(n491), .Y(sa32_next[7]) );
  XOR2X1 U1024 ( .A(n522), .B(n521), .Y(sa22_next[5]) );
  XOR2X1 U970 ( .A(n559), .B(n558), .Y(n556) );
  XOR2X1 U990 ( .A(n543), .B(n542), .Y(sa12_next[5]) );
  XOR2X1 U1085 ( .A(n774), .B(n773), .Y(n484) );
  XOR2X1 U1014 ( .A(n527), .B(n526), .Y(sa22_next[3]) );
  XOR2X1 U1028 ( .A(n520), .B(n519), .Y(sa22_next[6]) );
  XOR2X1 U969 ( .A(n780), .B(n793), .Y(n557) );
  XOR2X1 U1003 ( .A(n782), .B(n792), .Y(n532) );
  XOR2X1 U985 ( .A(n546), .B(n545), .Y(sa12_next[4]) );
  XOR2X1 U1070 ( .A(n495), .B(n494), .Y(sa32_next[6]) );
  XOR2X1 U975 ( .A(n554), .B(n553), .Y(sa12_next[2]) );
  XOR2X1 U1103 ( .A(n473), .B(n472), .Y(sa03_next[7]) );
  XOR2X1 U1065 ( .A(n498), .B(n497), .Y(sa32_next[5]) );
  XOR2X1 U1046 ( .A(n790), .B(n510), .Y(n508) );
  XOR2X1 U1082 ( .A(n775), .B(n488), .Y(n486) );
  XOR2X1 U998 ( .A(n537), .B(n536), .Y(sa12_next[7]) );
  XOR2X1 U1004 ( .A(n795), .B(n533), .Y(n531) );
  XOR2X1 U1059 ( .A(n501), .B(n500), .Y(sa32_next[4]) );
  XOR2X1 U994 ( .A(n540), .B(n539), .Y(sa12_next[6]) );
  XOR2X1 U1019 ( .A(n524), .B(n523), .Y(sa22_next[4]) );
  XOR2X1 U1032 ( .A(n518), .B(n517), .Y(sa22_next[7]) );
  XOR2X1 U1215 ( .A(n402), .B(n401), .Y(sa33_next[7]) );
  XOR2X1 U1008 ( .A(n790), .B(n793), .Y(n529) );
  XOR2X1 U980 ( .A(n550), .B(n549), .Y(sa12_next[3]) );
  XOR2X1 U901 ( .A(n604), .B(n603), .Y(n601) );
  XOR2X1 U1115 ( .A(n464), .B(n463), .Y(sa13_next[2]) );
  XOR2X1 U674 ( .A(n749), .B(n748), .Y(sa00_next[4]) );
  XOR2X1 U1110 ( .A(n469), .B(n468), .Y(n466) );
  XOR2X1 U670 ( .A(n752), .B(n751), .Y(sa00_next[3]) );
  XOR2X1 U1109 ( .A(n762), .B(n775), .Y(n467) );
  XOR2X1 U892 ( .A(n608), .B(n607), .Y(sa21_next[7]) );
  XOR2X1 U888 ( .A(n610), .B(n609), .Y(sa21_next[6]) );
  XOR2X1 U662 ( .A(n829), .B(n758), .Y(n756) );
  XOR2X1 U879 ( .A(n614), .B(n613), .Y(sa21_next[4]) );
  XOR2X1 U906 ( .A(n808), .B(n600), .Y(n598) );
  XOR2X1 U913 ( .A(n595), .B(n594), .Y(sa31_next[3]) );
  XOR2X1 U814 ( .A(n659), .B(n658), .Y(sa01_next[4]) );
  XOR2X1 U1172 ( .A(n428), .B(n427), .Y(sa23_next[7]) );
  XOR2X1 U817 ( .A(n657), .B(n656), .Y(sa01_next[5]) );
  XOR2X1 U659 ( .A(n760), .B(n759), .Y(sa00_next[0]) );
  XOR2X1 U718 ( .A(n717), .B(n716), .Y(sa10_next[7]) );
  XOR2X1 U823 ( .A(n653), .B(n652), .Y(sa01_next[7]) );
  XOR2X1 U714 ( .A(n720), .B(n719), .Y(sa10_next[6]) );
  XOR2X1 U756 ( .A(n696), .B(n695), .Y(sa30_next[0]) );
  XOR2X1 U710 ( .A(n723), .B(n722), .Y(sa10_next[5]) );
  XOR2X1 U760 ( .A(n815), .B(n828), .Y(n692) );
  XOR2X1 U1168 ( .A(n430), .B(n429), .Y(sa23_next[6]) );
  XOR2X1 U1164 ( .A(n432), .B(n431), .Y(sa23_next[5]) );
  XOR2X1 U761 ( .A(n694), .B(n693), .Y(n691) );
  XOR2X1 U874 ( .A(n617), .B(n616), .Y(sa21_next[3]) );
  XOR2X1 U868 ( .A(n808), .B(n811), .Y(n619) );
  XOR2X1 U864 ( .A(n813), .B(n623), .Y(n621) );
  XOR2X1 U863 ( .A(n800), .B(n810), .Y(n622) );
  XOR2X1 U925 ( .A(n588), .B(n587), .Y(sa31_next[5]) );
  XOR2X1 U1159 ( .A(n434), .B(n433), .Y(sa23_next[4]) );
  XOR2X1 U766 ( .A(n826), .B(n690), .Y(n688) );
  XOR2X1 U779 ( .A(n681), .B(n680), .Y(sa30_next[4]) );
  XOR2X1 U785 ( .A(n678), .B(n677), .Y(sa30_next[5]) );
  XOR2X1 U1041 ( .A(n514), .B(n513), .Y(n511) );
  XOR2X1 U790 ( .A(n675), .B(n674), .Y(sa30_next[6]) );
  XOR2X1 U795 ( .A(n672), .B(n671), .Y(sa30_next[7]) );
  XOR2X1 U1154 ( .A(n437), .B(n436), .Y(sa23_next[3]) );
  XOR2X1 U930 ( .A(n585), .B(n584), .Y(sa31_next[6]) );
  XOR2X1 U721 ( .A(n715), .B(n714), .Y(sa20_next[0]) );
  XOR2X1 U935 ( .A(n582), .B(n581), .Y(sa31_next[7]) );
  XOR2X1 U705 ( .A(n726), .B(n725), .Y(sa10_next[4]) );
  XOR2X1 U1148 ( .A(n772), .B(n775), .Y(n439) );
  XOR2X1 U723 ( .A(n818), .B(n828), .Y(n712) );
  XOR2X1 U724 ( .A(n831), .B(n713), .Y(n711) );
  XOR2X1 U728 ( .A(n826), .B(n829), .Y(n709) );
  XOR2X1 U700 ( .A(n730), .B(n729), .Y(sa10_next[3]) );
  XOR2X1 U695 ( .A(n734), .B(n733), .Y(sa10_next[2]) );
  XOR2X1 U734 ( .A(n707), .B(n706), .Y(sa20_next[3]) );
  XOR2X1 U690 ( .A(n739), .B(n738), .Y(n736) );
  XOR2X1 U739 ( .A(n704), .B(n703), .Y(sa20_next[4]) );
  XOR2X1 U689 ( .A(n816), .B(n829), .Y(n737) );
  XOR2X1 U748 ( .A(n700), .B(n699), .Y(sa20_next[6]) );
  XOR2X1 U752 ( .A(n698), .B(n697), .Y(sa20_next[7]) );
  XOR2X1 U1210 ( .A(n405), .B(n404), .Y(sa33_next[6]) );
  XOR2X1 U686 ( .A(n741), .B(n740), .Y(sa10_next[0]) );
  XOR2X1 U1040 ( .A(n779), .B(n792), .Y(n512) );
  XOR2X1 U1193 ( .A(n415), .B(n414), .Y(sa33_next[3]) );
  XOR2X1 U1138 ( .A(n447), .B(n446), .Y(sa13_next[7]) );
  XOR2X1 U1186 ( .A(n772), .B(n420), .Y(n418) );
  XOR2X1 U802 ( .A(n811), .B(n668), .Y(n666) );
  XOR2X1 U957 ( .A(n567), .B(n566), .Y(sa02_next[5]) );
  XOR2X1 U954 ( .A(n569), .B(n568), .Y(sa02_next[4]) );
  XOR2X1 U683 ( .A(n743), .B(n742), .Y(sa00_next[7]) );
  XOR2X1 U805 ( .A(n810), .B(n809), .Y(n664) );
  XOR2X1 U1199 ( .A(n411), .B(n410), .Y(sa33_next[4]) );
  XOR2X1 U1134 ( .A(n450), .B(n449), .Y(sa13_next[6]) );
  XOR2X1 U845 ( .A(n636), .B(n635), .Y(sa11_next[4]) );
  XOR2X1 U840 ( .A(n640), .B(n639), .Y(sa11_next[3]) );
  XOR2X1 U1090 ( .A(n482), .B(n481), .Y(sa03_next[3]) );
  XOR2X1 U835 ( .A(n644), .B(n643), .Y(sa11_next[2]) );
  XOR2X1 U850 ( .A(n633), .B(n632), .Y(sa11_next[5]) );
  XOR2X1 U858 ( .A(n627), .B(n626), .Y(sa11_next[7]) );
  XOR2X1 U960 ( .A(n565), .B(n564), .Y(sa02_next[6]) );
  XOR2X1 U1130 ( .A(n453), .B(n452), .Y(sa13_next[5]) );
  XOR2X1 U950 ( .A(n572), .B(n571), .Y(sa02_next[3]) );
  XOR2X1 U1205 ( .A(n408), .B(n407), .Y(sa33_next[5]) );
  XOR2X1 U830 ( .A(n649), .B(n648), .Y(n646) );
  XOR2X1 U942 ( .A(n793), .B(n578), .Y(n576) );
  XOR2X1 U1144 ( .A(n777), .B(n443), .Y(n441) );
  XOR2X1 U963 ( .A(n563), .B(n562), .Y(sa02_next[7]) );
  XOR2X1 U829 ( .A(n798), .B(n811), .Y(n647) );
  XOR2X1 U1141 ( .A(n445), .B(n444), .Y(sa23_next[0]) );
  XOR2X1 U1143 ( .A(n764), .B(n774), .Y(n442) );
  XOR2X1 U1180 ( .A(n761), .B(n774), .Y(n422) );
  XOR2X1 U945 ( .A(n792), .B(n791), .Y(n574) );
  XOR2X1 U677 ( .A(n747), .B(n746), .Y(sa00_next[5]) );
  XOR2X1 U1125 ( .A(n456), .B(n455), .Y(sa13_next[4]) );
  XOR2X1 U854 ( .A(n630), .B(n629), .Y(sa11_next[6]) );
  XOR2X1 U1120 ( .A(n460), .B(n459), .Y(sa13_next[3]) );
  XOR2X1 U1176 ( .A(n426), .B(n425), .Y(sa33_next[0]) );
  XOR2X1 U1094 ( .A(n479), .B(n478), .Y(sa03_next[4]) );
  XOR2X1 U1181 ( .A(n424), .B(n423), .Y(n421) );
  XOR2X1 U900 ( .A(n797), .B(n810), .Y(n602) );
  XOR2X1 U1079 ( .A(n490), .B(n489), .Y(sa03_next[0]) );
  XOR2X1 U810 ( .A(n662), .B(n661), .Y(sa01_next[3]) );
  XOR2X1 U1009 ( .A(n530), .B(n529), .Y(sa22_next[2]) );
  XOR2X1 U1047 ( .A(n509), .B(n508), .Y(sa32_next[2]) );
  XOR2X1 U1005 ( .A(n532), .B(n531), .Y(sa22_next[1]) );
  XOR2X1 U803 ( .A(n667), .B(n666), .Y(sa01_next[1]) );
  XOR2X1 U806 ( .A(n665), .B(n664), .Y(sa01_next[2]) );
  XOR2X1 U1086 ( .A(n485), .B(n484), .Y(sa03_next[2]) );
  XOR2X1 U1042 ( .A(n512), .B(n511), .Y(sa32_next[1]) );
  XOR2X1 U1187 ( .A(n419), .B(n418), .Y(sa33_next[2]) );
  XOR2X1 U1182 ( .A(n422), .B(n421), .Y(sa33_next[1]) );
  XOR2X1 U663 ( .A(n757), .B(n756), .Y(sa00_next[1]) );
  XOR2X1 U762 ( .A(n692), .B(n691), .Y(sa30_next[1]) );
  XOR2X1 U767 ( .A(n689), .B(n688), .Y(sa30_next[2]) );
  XOR2X1 U725 ( .A(n712), .B(n711), .Y(sa20_next[1]) );
  XOR2X1 U729 ( .A(n710), .B(n709), .Y(sa20_next[2]) );
  XOR2X1 U691 ( .A(n737), .B(n736), .Y(sa10_next[1]) );
  XOR2X1 U971 ( .A(n557), .B(n556), .Y(sa12_next[1]) );
  XOR2X1 U1083 ( .A(n487), .B(n486), .Y(sa03_next[1]) );
  XOR2X1 U1149 ( .A(n440), .B(n439), .Y(sa23_next[2]) );
  XOR2X1 U907 ( .A(n599), .B(n598), .Y(sa31_next[2]) );
  XOR2X1 U1111 ( .A(n467), .B(n466), .Y(sa13_next[1]) );
  XOR2X1 U831 ( .A(n647), .B(n646), .Y(sa11_next[1]) );
  XOR2X1 U902 ( .A(n602), .B(n601), .Y(sa31_next[1]) );
  XOR2X1 U869 ( .A(n620), .B(n619), .Y(sa21_next[2]) );
  XOR2X1 U865 ( .A(n622), .B(n621), .Y(sa21_next[1]) );
  XOR2X1 U946 ( .A(n575), .B(n574), .Y(sa02_next[2]) );
  XOR2X1 U1145 ( .A(n442), .B(n441), .Y(sa23_next[1]) );
  XOR2X1 U943 ( .A(n577), .B(n576), .Y(sa02_next[1]) );
  XOR2X1 U688 ( .A(sa10_sr[0]), .B(sa20_sr[0]), .Y(n738) );
  XOR2X1 U1108 ( .A(sa13_sr[0]), .B(sa23_sr[0]), .Y(n468) );
  XOR2X1 U968 ( .A(sa12_sr[0]), .B(sa22_sr[0]), .Y(n558) );
  XOR2X1 U828 ( .A(sa11_sr[0]), .B(sa21_sr[0]), .Y(n648) );
  XOR2XL U1213 ( .A(sa23_sr[7]), .B(sa33_sr[6]), .Y(n402) );
  XOR2XL U933 ( .A(sa21_sr[7]), .B(sa31_sr[6]), .Y(n582) );
  XOR2XL U1073 ( .A(sa22_sr[7]), .B(sa32_sr[6]), .Y(n492) );
  XOR2X1 U941 ( .A(n796), .B(n794), .Y(n577) );
  XOR2X1 U1102 ( .A(n764), .B(n763), .Y(n472) );
  XOR2X1 U661 ( .A(n832), .B(n830), .Y(n757) );
  DFFTRXL dcnt_reg_3_ ( .D(n1187), .RN(rst), .CK(divclk), .QN(n2) );
  AOI21X1 U1217 ( .A0(w1[4]), .A1(text_in_r[68]), .B0(n4), .Y(n833) );
  OAI21XL U1218 ( .A0(w1[4]), .A1(text_in_r[68]), .B0(n833), .Y(n834) );
  AOI2BB2X1 U1219 ( .B0(w1[4]), .B1(sa01_sr[3]), .A0N(sa01_sr[3]), .A1N(w1[4]), 
        .Y(n835) );
  INVX1 U1220 ( .A(sa31_sr[3]), .Y(n836) );
  AOI2BB2X1 U1221 ( .B0(sa21_sr[4]), .B1(n836), .A0N(n836), .A1N(sa21_sr[4]), 
        .Y(n837) );
  XOR2X1 U1222 ( .A(n835), .B(n837), .Y(n838) );
  NAND2X1 U1223 ( .A(n838), .B(n804), .Y(n839) );
  OAI21XL U1224 ( .A0(n838), .A1(n804), .B0(n839), .Y(n840) );
  INVX1 U1225 ( .A(n4), .Y(n841) );
  AOI21X1 U1226 ( .A0(n797), .A1(n840), .B0(n841), .Y(n842) );
  OAI21XL U1227 ( .A0(n797), .A1(n840), .B0(n842), .Y(n843) );
  NAND2X1 U1228 ( .A(n834), .B(n843), .Y(N164) );
  AOI2BB2X1 U1229 ( .B0(w2[3]), .B1(sa02_sr[2]), .A0N(sa02_sr[2]), .A1N(w2[3]), 
        .Y(n844) );
  INVX1 U1230 ( .A(sa32_sr[2]), .Y(n845) );
  AOI2BB2X1 U1231 ( .B0(sa22_sr[3]), .B1(n845), .A0N(n845), .A1N(sa22_sr[3]), 
        .Y(n846) );
  XOR2X1 U1232 ( .A(n844), .B(n846), .Y(n847) );
  NAND2X1 U1233 ( .A(n847), .B(n788), .Y(n848) );
  OAI21XL U1234 ( .A0(n847), .A1(n788), .B0(n848), .Y(n849) );
  OAI21XL U1235 ( .A0(n779), .A1(n849), .B0(n4), .Y(n850) );
  AOI21X1 U1236 ( .A0(n779), .A1(n849), .B0(n850), .Y(n851) );
  NOR2X1 U1237 ( .A(text_in_r[35]), .B(w2[3]), .Y(n852) );
  AOI211X1 U1238 ( .A0(text_in_r[35]), .A1(w2[3]), .B0(n965), .C0(n852), .Y(
        n853) );
  OR2X1 U1239 ( .A(n851), .B(n853), .Y(N99) );
  AOI2BB2X1 U1240 ( .B0(w2[16]), .B1(n780), .A0N(n780), .A1N(w2[16]), .Y(n854)
         );
  AOI2BB2X1 U1241 ( .B0(sa02_sr[0]), .B1(n795), .A0N(n795), .A1N(sa02_sr[0]), 
        .Y(n855) );
  NAND2X1 U1242 ( .A(n854), .B(n855), .Y(n856) );
  OAI211X1 U1243 ( .A0(n854), .A1(n855), .B0(n4), .C0(n856), .Y(n857) );
  AOI21XL U1244 ( .A0(w2[16]), .A1(text_in_r[48]), .B0(n964), .Y(n858) );
  OAI21XL U1245 ( .A0(w2[16]), .A1(text_in_r[48]), .B0(n858), .Y(n859) );
  NAND2X1 U1246 ( .A(n857), .B(n859), .Y(N128) );
  AOI2BB2X1 U1247 ( .B0(w1[16]), .B1(n798), .A0N(n798), .A1N(w1[16]), .Y(n860)
         );
  AOI2BB2X1 U1248 ( .B0(sa01_sr[0]), .B1(n813), .A0N(n813), .A1N(sa01_sr[0]), 
        .Y(n861) );
  NAND2X1 U1249 ( .A(n860), .B(n861), .Y(n862) );
  OAI211X1 U1250 ( .A0(n860), .A1(n861), .B0(n4), .C0(n862), .Y(n863) );
  AOI21XL U1251 ( .A0(w1[16]), .A1(text_in_r[80]), .B0(n963), .Y(n864) );
  OAI21XL U1252 ( .A0(w1[16]), .A1(text_in_r[80]), .B0(n864), .Y(n865) );
  NAND2X1 U1253 ( .A(n863), .B(n865), .Y(N192) );
  AOI2BB2X1 U1254 ( .B0(w2[0]), .B1(n779), .A0N(n779), .A1N(w2[0]), .Y(n866)
         );
  AOI2BB2X1 U1255 ( .B0(sa22_sr[0]), .B1(n794), .A0N(n794), .A1N(sa22_sr[0]), 
        .Y(n867) );
  NAND2X1 U1256 ( .A(n866), .B(n867), .Y(n868) );
  OAI211X1 U1257 ( .A0(n866), .A1(n867), .B0(n4), .C0(n868), .Y(n869) );
  AOI21X1 U1258 ( .A0(w2[0]), .A1(text_in_r[32]), .B0(n965), .Y(n870) );
  OAI21XL U1259 ( .A0(w2[0]), .A1(text_in_r[32]), .B0(n870), .Y(n871) );
  NAND2X1 U1260 ( .A(n869), .B(n871), .Y(N96) );
  AOI2BB2X1 U1261 ( .B0(w1[24]), .B1(n814), .A0N(n814), .A1N(w1[24]), .Y(n872)
         );
  AOI2BB2X1 U1262 ( .B0(sa11_sr[0]), .B1(n813), .A0N(n813), .A1N(sa11_sr[0]), 
        .Y(n873) );
  NAND2X1 U1263 ( .A(n872), .B(n873), .Y(n874) );
  OAI211X1 U1264 ( .A0(n872), .A1(n873), .B0(n4), .C0(n874), .Y(n875) );
  AOI21XL U1265 ( .A0(w1[24]), .A1(text_in_r[88]), .B0(n963), .Y(n876) );
  OAI21XL U1266 ( .A0(w1[24]), .A1(text_in_r[88]), .B0(n876), .Y(n877) );
  NAND2X1 U1267 ( .A(n875), .B(n877), .Y(N208) );
  INVX1 U1268 ( .A(n4), .Y(n878) );
  AOI2BB2X1 U1269 ( .B0(n795), .B1(sa12_sr[0]), .A0N(sa12_sr[0]), .A1N(n795), 
        .Y(n879) );
  OAI21XL U1270 ( .A0(n796), .A1(n879), .B0(n4), .Y(n880) );
  AOI21X1 U1271 ( .A0(n796), .A1(n879), .B0(n880), .Y(n881) );
  AOI21X1 U1272 ( .A0(text_in_r[56]), .A1(n878), .B0(n881), .Y(n882) );
  XNOR2X1 U1273 ( .A(n882), .B(w2[24]), .Y(N144) );
  AOI2BB2X1 U1274 ( .B0(w1[0]), .B1(n797), .A0N(n797), .A1N(w1[0]), .Y(n883)
         );
  AOI2BB2X1 U1275 ( .B0(sa21_sr[0]), .B1(n812), .A0N(n812), .A1N(sa21_sr[0]), 
        .Y(n884) );
  NAND2X1 U1276 ( .A(n883), .B(n884), .Y(n885) );
  OAI211X1 U1277 ( .A0(n883), .A1(n884), .B0(n4), .C0(n885), .Y(n886) );
  AOI21XL U1278 ( .A0(w1[0]), .A1(text_in_r[64]), .B0(n963), .Y(n887) );
  OAI21XL U1279 ( .A0(w1[0]), .A1(text_in_r[64]), .B0(n887), .Y(n888) );
  NAND2X1 U1280 ( .A(n886), .B(n888), .Y(N160) );
  AOI2BB2X1 U1281 ( .B0(w0[26]), .B1(n828), .A0N(n828), .A1N(w0[26]), .Y(n889)
         );
  AOI2BB2X1 U1282 ( .B0(sa10_sr[2]), .B1(n827), .A0N(n827), .A1N(sa10_sr[2]), 
        .Y(n890) );
  NAND2X1 U1283 ( .A(n889), .B(n890), .Y(n891) );
  OAI211X1 U1284 ( .A0(n889), .A1(n890), .B0(n4), .C0(n891), .Y(n892) );
  AOI21XL U1285 ( .A0(w0[26]), .A1(text_in_r[122]), .B0(n961), .Y(n893) );
  OAI21XL U1286 ( .A0(w0[26]), .A1(text_in_r[122]), .B0(n893), .Y(n894) );
  NAND2X1 U1287 ( .A(n892), .B(n894), .Y(N274) );
  AOI2BB2X1 U1288 ( .B0(w3[29]), .B1(n768), .A0N(n768), .A1N(w3[29]), .Y(n895)
         );
  AOI2BB2X1 U1289 ( .B0(sa13_sr[5]), .B1(n767), .A0N(n767), .A1N(sa13_sr[5]), 
        .Y(n896) );
  NAND2X1 U1290 ( .A(n895), .B(n896), .Y(n897) );
  OAI211X1 U1291 ( .A0(n895), .A1(n896), .B0(n965), .C0(n897), .Y(n898) );
  AOI21XL U1292 ( .A0(w3[29]), .A1(text_in_r[29]), .B0(n964), .Y(n899) );
  OAI21XL U1293 ( .A0(w3[29]), .A1(text_in_r[29]), .B0(n899), .Y(n900) );
  NAND2X1 U1294 ( .A(n898), .B(n900), .Y(N85) );
  AOI2BB2X1 U1295 ( .B0(w0[13]), .B1(n820), .A0N(n820), .A1N(w0[13]), .Y(n901)
         );
  AOI2BB2X1 U1296 ( .B0(sa30_sr[5]), .B1(n823), .A0N(n823), .A1N(sa30_sr[5]), 
        .Y(n902) );
  NAND2X1 U1297 ( .A(n901), .B(n902), .Y(n903) );
  OAI211X1 U1298 ( .A0(n901), .A1(n902), .B0(n4), .C0(n903), .Y(n904) );
  AOI21XL U1299 ( .A0(w0[13]), .A1(text_in_r[109]), .B0(n961), .Y(n905) );
  OAI21XL U1300 ( .A0(w0[13]), .A1(text_in_r[109]), .B0(n905), .Y(n906) );
  NAND2X1 U1301 ( .A(n904), .B(n906), .Y(N245) );
  AOI2BB2X1 U1302 ( .B0(w1[13]), .B1(n802), .A0N(n802), .A1N(w1[13]), .Y(n907)
         );
  AOI2BB2X1 U1303 ( .B0(sa31_sr[5]), .B1(n805), .A0N(n805), .A1N(sa31_sr[5]), 
        .Y(n908) );
  NAND2X1 U1304 ( .A(n907), .B(n908), .Y(n909) );
  OAI211X1 U1305 ( .A0(n907), .A1(n908), .B0(n4), .C0(n909), .Y(n910) );
  AOI21XL U1306 ( .A0(w1[13]), .A1(text_in_r[77]), .B0(n963), .Y(n911) );
  OAI21XL U1307 ( .A0(w1[13]), .A1(text_in_r[77]), .B0(n911), .Y(n912) );
  NAND2X1 U1308 ( .A(n910), .B(n912), .Y(N181) );
  INVX1 U1309 ( .A(n4), .Y(n913) );
  AOI2BB2X1 U1310 ( .B0(n812), .B1(sa31_sr[0]), .A0N(sa31_sr[0]), .A1N(n812), 
        .Y(n914) );
  OAI21XL U1311 ( .A0(n800), .A1(n914), .B0(n4), .Y(n915) );
  AOI21X1 U1312 ( .A0(n800), .A1(n914), .B0(n915), .Y(n916) );
  AOI21X1 U1313 ( .A0(text_in_r[72]), .A1(n913), .B0(n916), .Y(n917) );
  XNOR2X1 U1314 ( .A(n917), .B(w1[8]), .Y(N176) );
  AOI21X1 U1315 ( .A0(w0[3]), .A1(text_in_r[99]), .B0(n4), .Y(n918) );
  OAI21XL U1316 ( .A0(w0[3]), .A1(text_in_r[99]), .B0(n918), .Y(n919) );
  INVX1 U1317 ( .A(n4), .Y(n920) );
  AOI2BB2X1 U1318 ( .B0(w0[3]), .B1(sa00_sr[2]), .A0N(sa00_sr[2]), .A1N(w0[3]), 
        .Y(n921) );
  AOI2BB2X1 U1319 ( .B0(sa20_sr[3]), .B1(n922), .A0N(n922), .A1N(sa20_sr[3]), 
        .Y(n923) );
  XOR2X1 U1320 ( .A(n921), .B(n923), .Y(n924) );
  NAND2X1 U1321 ( .A(n924), .B(n824), .Y(n925) );
  OAI21XL U1322 ( .A0(n924), .A1(n824), .B0(n925), .Y(n926) );
  AOI21X1 U1323 ( .A0(n815), .A1(n926), .B0(n920), .Y(n927) );
  OAI21XL U1324 ( .A0(n815), .A1(n926), .B0(n927), .Y(n928) );
  NAND2X1 U1325 ( .A(n919), .B(n928), .Y(N227) );
  INVX1 U1326 ( .A(sa30_sr[2]), .Y(n922) );
  AOI2BB2X1 U1327 ( .B0(w3[16]), .B1(n762), .A0N(n762), .A1N(w3[16]), .Y(n929)
         );
  AOI2BB2X1 U1328 ( .B0(sa03_sr[0]), .B1(n777), .A0N(n777), .A1N(sa03_sr[0]), 
        .Y(n930) );
  NAND2X1 U1329 ( .A(n929), .B(n930), .Y(n931) );
  OAI211X1 U1330 ( .A0(n929), .A1(n930), .B0(n965), .C0(n931), .Y(n932) );
  AOI21X1 U1331 ( .A0(w3[16]), .A1(text_in_r[16]), .B0(n963), .Y(n933) );
  OAI21XL U1332 ( .A0(w3[16]), .A1(text_in_r[16]), .B0(n933), .Y(n934) );
  NAND2X1 U1333 ( .A(n932), .B(n934), .Y(N64) );
  AOI2BB2X1 U1334 ( .B0(w2[8]), .B1(n782), .A0N(n782), .A1N(w2[8]), .Y(n935)
         );
  AOI2BB2X1 U1335 ( .B0(sa32_sr[0]), .B1(n794), .A0N(n794), .A1N(sa32_sr[0]), 
        .Y(n936) );
  NAND2X1 U1336 ( .A(n935), .B(n936), .Y(n937) );
  OAI211X1 U1337 ( .A0(n935), .A1(n936), .B0(n4), .C0(n937), .Y(n938) );
  AOI21X1 U1338 ( .A0(w2[8]), .A1(text_in_r[40]), .B0(n965), .Y(n939) );
  OAI21XL U1339 ( .A0(w2[8]), .A1(text_in_r[40]), .B0(n939), .Y(n940) );
  NAND2X1 U1340 ( .A(n938), .B(n940), .Y(N112) );
  AOI2BB2X1 U1341 ( .B0(w0[30]), .B1(n820), .A0N(n820), .A1N(w0[30]), .Y(n941)
         );
  AOI2BB2X1 U1342 ( .B0(sa10_sr[6]), .B1(n819), .A0N(n819), .A1N(sa10_sr[6]), 
        .Y(n942) );
  NAND2X1 U1343 ( .A(n941), .B(n942), .Y(n943) );
  OAI211X1 U1344 ( .A0(n941), .A1(n942), .B0(n4), .C0(n943), .Y(n944) );
  AOI21X1 U1345 ( .A0(w0[30]), .A1(text_in_r[126]), .B0(n961), .Y(n945) );
  OAI21XL U1346 ( .A0(w0[30]), .A1(text_in_r[126]), .B0(n945), .Y(n946) );
  NAND2X1 U1347 ( .A(n944), .B(n946), .Y(N278) );
  AOI2BB2X1 U1348 ( .B0(w3[30]), .B1(n766), .A0N(n766), .A1N(w3[30]), .Y(n947)
         );
  AOI2BB2X1 U1349 ( .B0(sa13_sr[6]), .B1(n765), .A0N(n765), .A1N(sa13_sr[6]), 
        .Y(n948) );
  NAND2X1 U1350 ( .A(n947), .B(n948), .Y(n949) );
  OAI211X1 U1351 ( .A0(n947), .A1(n948), .B0(n965), .C0(n949), .Y(n950) );
  AOI21X1 U1352 ( .A0(w3[30]), .A1(text_in_r[30]), .B0(n964), .Y(n951) );
  OAI21XL U1353 ( .A0(w3[30]), .A1(text_in_r[30]), .B0(n951), .Y(n952) );
  NAND2X1 U1354 ( .A(n950), .B(n952), .Y(N86) );
  AOI2BB2X1 U1355 ( .B0(w1[30]), .B1(n802), .A0N(n802), .A1N(w1[30]), .Y(n953)
         );
  AOI2BB2X1 U1356 ( .B0(sa11_sr[6]), .B1(n801), .A0N(n801), .A1N(sa11_sr[6]), 
        .Y(n954) );
  NAND2X1 U1357 ( .A(n953), .B(n954), .Y(n955) );
  OAI211X1 U1358 ( .A0(n953), .A1(n954), .B0(n4), .C0(n955), .Y(n956) );
  AOI21X1 U1359 ( .A0(w1[30]), .A1(text_in_r[94]), .B0(n962), .Y(n957) );
  OAI21XL U1360 ( .A0(w1[30]), .A1(text_in_r[94]), .B0(n957), .Y(n958) );
  NAND2X1 U1361 ( .A(n956), .B(n958), .Y(N214) );
  OAI2BB1XL U1362 ( .A0N(n4), .A1N(sa00_next[1]), .B0(n1115), .Y(N273) );
  OAI2BB1XL U1363 ( .A0N(n4), .A1N(sa22_next[1]), .B0(n976), .Y(N113) );
  OAI2BB1XL U1364 ( .A0N(n4), .A1N(sa02_next[1]), .B0(n1004), .Y(N145) );
  OAI2BB1XL U1365 ( .A0N(n4), .A1N(sa20_next[2]), .B0(n1087), .Y(N242) );
  OAI2BB1XL U1366 ( .A0N(n4), .A1N(sa20_next[1]), .B0(n1085), .Y(N241) );
  OAI2BB1XL U1367 ( .A0N(n4), .A1N(sa21_next[1]), .B0(n1030), .Y(N177) );
  OAI2BB1XL U1368 ( .A0N(n4), .A1N(sa12_next[1]), .B0(n990), .Y(N129) );
  OAI2BB1XL U1369 ( .A0N(n4), .A1N(sa32_next[2]), .B0(n1185), .Y(N98) );
  OAI2BB1XL U1370 ( .A0N(n4), .A1N(sa02_next[2]), .B0(n1006), .Y(N146) );
  OAI2BB1XL U1371 ( .A0N(n4), .A1N(sa21_next[2]), .B0(n1032), .Y(N178) );
  OAI2BB1XL U1372 ( .A0N(n4), .A1N(sa03_next[2]), .B0(n1175), .Y(N82) );
//wddl
 
//  OAI2BB1XL U1373 ( .A0N(n4), .A1N(sa23_next[1]), .B0(n1143), .Y(N49) );
  CLKINVX3 Uwddlclk ( .A(divclk), .Y(clk_bar));
  WDDLNANDCOMP U1373 ( .A(n4), .B(sa23_next[1]) , .C(n1143), .clkinv(clk_bar), .Y(N49) , .Y_bar(N49inv));  
  OAI2BB1XL U1374 ( .A0N(n4), .A1N(sa01_next[2]), .B0(n1059), .Y(N210) );
  OAI2BB1XL U1375 ( .A0N(n4), .A1N(sa30_next[1]), .B0(n1071), .Y(N225) );
  OAI2BB1XL U1376 ( .A0N(n4), .A1N(sa31_next[1]), .B0(n1018), .Y(N161) );
  OAI2BB1XL U1377 ( .A0N(n4), .A1N(sa10_next[1]), .B0(n1099), .Y(N257) );
  OAI2BB1XL U1378 ( .A0N(n4), .A1N(sa22_next[2]), .B0(n978), .Y(N114) );
  OAI2BB1XL U1379 ( .A0N(n4), .A1N(sa30_next[2]), .B0(n1073), .Y(N226) );
  OAI2BB1XL U1380 ( .A0N(n4), .A1N(sa01_next[1]), .B0(n1056), .Y(N209) );
  OAI2BB1XL U1381 ( .A0N(n4), .A1N(sa31_next[2]), .B0(n1020), .Y(N162) );
  OAI2BB1XL U1382 ( .A0N(n4), .A1N(sa33_next[2]), .B0(n1129), .Y(N34) );
  OAI2BB1XL U1383 ( .A0N(n4), .A1N(sa11_next[1]), .B0(n1042), .Y(N193) );
  OAI2BB1XL U1384 ( .A0N(n4), .A1N(sa11_next[7]), .B0(n1054), .Y(N199) );
  OAI2BB1XL U1385 ( .A0N(n4), .A1N(sa03_next[3]), .B0(n1177), .Y(N83) );
  OAI2BB1XL U1386 ( .A0N(n4), .A1N(sa00_next[7]), .B0(n1123), .Y(N279) );
  OAI2BB1XL U1387 ( .A0N(n4), .A1N(sa22_next[5]), .B0(n984), .Y(N117) );
  OAI2BB1XL U1388 ( .A0N(n4), .A1N(sa11_next[3]), .B0(n1046), .Y(N195) );
  OAI2BB1XL U1389 ( .A0N(n4), .A1N(sa32_next[7]), .B0(n974), .Y(N103) );
  OAI2BB1XL U1390 ( .A0N(n4), .A1N(sa01_next[5]), .B0(n1065), .Y(N213) );
  OAI2BB1XL U1391 ( .A0N(n4), .A1N(sa22_next[7]), .B0(n988), .Y(N119) );
  OAI2BB1XL U1392 ( .A0N(n4), .A1N(sa00_next[5]), .B0(n1121), .Y(N277) );
  OAI2BB1XL U1393 ( .A0N(n4), .A1N(sa21_next[7]), .B0(n1040), .Y(N183) );
  OAI2BB1XL U1394 ( .A0N(n4), .A1N(sa00_next[4]), .B0(n1119), .Y(N276) );
  OAI2BB1XL U1395 ( .A0N(n4), .A1N(sa12_next[4]), .B0(n996), .Y(N132) );
  OAI2BB1XL U1396 ( .A0N(n4), .A1N(sa13_next[7]), .B0(n1169), .Y(N71) );
  OAI2BB1XL U1397 ( .A0N(n4), .A1N(sa01_next[3]), .B0(n1061), .Y(N211) );
  OAI2BB1XL U1398 ( .A0N(n4), .A1N(sa23_next[0]), .B0(n1141), .Y(N48) );
  OAI2BB1XL U1399 ( .A0N(n4), .A1N(sa12_next[3]), .B0(n994), .Y(N131) );
  OAI2BB1XL U1400 ( .A0N(n4), .A1N(sa11_next[2]), .B0(n1044), .Y(N194) );
  OAI2BB1XL U1401 ( .A0N(n4), .A1N(sa22_next[3]), .B0(n980), .Y(N115) );
  OAI2BB1XL U1402 ( .A0N(n4), .A1N(sa01_next[7]), .B0(n1067), .Y(N215) );
  OAI2BB1XL U1403 ( .A0N(n4), .A1N(sa22_next[4]), .B0(n982), .Y(N116) );
  OAI2BB1XL U1404 ( .A0N(n4), .A1N(sa01_next[4]), .B0(n1063), .Y(N212) );
  OAI2BB1XL U1405 ( .A0N(n4), .A1N(sa03_next[4]), .B0(n1179), .Y(N84) );
  OAI2BB1XL U1406 ( .A0N(n4), .A1N(sa12_next[7]), .B0(n1002), .Y(N135) );
  OAI2BB1XL U1407 ( .A0N(n4), .A1N(sa20_next[0]), .B0(n1083), .Y(N240) );
  OAI2BB1XL U1408 ( .A0N(n4), .A1N(sa31_next[7]), .B0(n1028), .Y(N167) );
  OAI2BB1XL U1409 ( .A0N(n4), .A1N(sa02_next[3]), .B0(n1008), .Y(N147) );
  OAI2BB1XL U1410 ( .A0N(n4), .A1N(sa30_next[7]), .B0(n1081), .Y(N231) );
  OAI2BB1XL U1411 ( .A0N(n4), .A1N(sa20_next[7]), .B0(n1095), .Y(N247) );
  OAI2BB1XL U1412 ( .A0N(n4), .A1N(sa21_next[3]), .B0(n1034), .Y(N179) );
  OAI2BB1XL U1413 ( .A0N(n4), .A1N(sa10_next[0]), .B0(n1097), .Y(N256) );
  OAI2BB1XL U1414 ( .A0N(n4), .A1N(sa21_next[4]), .B0(n1036), .Y(N180) );
  OAI2BB1XL U1415 ( .A0N(n4), .A1N(sa10_next[7]), .B0(n1111), .Y(N263) );
  OAI2BB1XL U1416 ( .A0N(n4), .A1N(sa00_next[3]), .B0(n1117), .Y(N275) );
  OAI2BB1XL U1417 ( .A0N(n4), .A1N(sa31_next[5]), .B0(n1024), .Y(N165) );
  OAI2BB1XL U1418 ( .A0N(n4), .A1N(sa10_next[4]), .B0(n1105), .Y(N260) );
  OAI2BB1XL U1419 ( .A0N(n4), .A1N(sa02_next[4]), .B0(n1010), .Y(N148) );
  OAI2BB1XL U1420 ( .A0N(n4), .A1N(sa11_next[4]), .B0(n1048), .Y(N196) );
  OAI2BB1XL U1421 ( .A0N(n4), .A1N(sa20_next[3]), .B0(n1089), .Y(N243) );
  OAI2BB1XL U1422 ( .A0N(n4), .A1N(sa02_next[7]), .B0(n1016), .Y(N151) );
  OAI2BB1XL U1423 ( .A0N(n4), .A1N(sa32_next[5]), .B0(n970), .Y(N101) );
  OAI2BB1XL U1424 ( .A0N(n4), .A1N(sa30_next[5]), .B0(n1077), .Y(N229) );
  OAI2BB1XL U1425 ( .A0N(n4), .A1N(sa02_next[5]), .B0(n1012), .Y(N149) );
  OAI2BB1XL U1426 ( .A0N(n4), .A1N(sa00_next[0]), .B0(n1113), .Y(N272) );
  OAI2BB1XL U1427 ( .A0N(n4), .A1N(sa20_next[4]), .B0(n1091), .Y(N244) );
  OAI2BB1XL U1428 ( .A0N(n4), .A1N(sa10_next[3]), .B0(n1103), .Y(N259) );
  OAI2BB1XL U1429 ( .A0N(n4), .A1N(sa30_next[6]), .B0(n1079), .Y(N230) );
  OAI2BB1XL U1430 ( .A0N(n4), .A1N(sa10_next[5]), .B0(n1107), .Y(N261) );
  OAI2BB1XL U1431 ( .A0N(n4), .A1N(sa20_next[6]), .B0(n1093), .Y(N246) );
  OAI2BB1XL U1432 ( .A0N(n4), .A1N(sa12_next[6]), .B0(n1000), .Y(N134) );
  OAI2BB1XL U1433 ( .A0N(n4), .A1N(sa21_next[6]), .B0(n1038), .Y(N182) );
  OAI2BB1XL U1434 ( .A0N(n4), .A1N(sa31_next[6]), .B0(n1026), .Y(N166) );
  OAI2BB1XL U1435 ( .A0N(n4), .A1N(sa11_next[5]), .B0(n1050), .Y(N197) );
  OAI2BB1XL U1436 ( .A0N(n4), .A1N(sa11_next[6]), .B0(n1052), .Y(N198) );
  OAI2BB1XL U1437 ( .A0N(n4), .A1N(sa02_next[6]), .B0(n1014), .Y(N150) );
  OAI2BB1XL U1438 ( .A0N(n4), .A1N(sa31_next[3]), .B0(n1022), .Y(N163) );
  OAI2BB1XL U1439 ( .A0N(n4), .A1N(sa32_next[4]), .B0(n968), .Y(N100) );
  OAI2BB1XL U1440 ( .A0N(n4), .A1N(sa03_next[7]), .B0(n1181), .Y(N87) );
  OAI2BB1XL U1441 ( .A0N(n4), .A1N(sa30_next[0]), .B0(n1069), .Y(N224) );
  OAI2BB1XL U1442 ( .A0N(n4), .A1N(sa30_next[4]), .B0(n1075), .Y(N228) );
  CLKINVX3 U1443 ( .A(n960), .Y(n965) );
  OAI2BB1XL U1444 ( .A0N(n965), .A1N(sa23_next[2]), .B0(n1145), .Y(N50) );
  OAI2BB1XL U1445 ( .A0N(n965), .A1N(sa03_next[1]), .B0(n1173), .Y(N81) );
  OAI2BB1XL U1446 ( .A0N(n965), .A1N(sa32_next[1]), .B0(n1183), .Y(N97) );
  OAI2BB1XL U1447 ( .A0N(n965), .A1N(sa13_next[6]), .B0(n1167), .Y(N70) );
  OAI2BB1XL U1448 ( .A0N(n965), .A1N(sa13_next[5]), .B0(n1165), .Y(N69) );
  OAI2BB1XL U1449 ( .A0N(n965), .A1N(sa23_next[3]), .B0(n1147), .Y(N51) );
  OAI2BB1XL U1450 ( .A0N(n965), .A1N(sa13_next[4]), .B0(n1163), .Y(N68) );
  OAI2BB1XL U1451 ( .A0N(n965), .A1N(sa23_next[4]), .B0(n1149), .Y(N52) );
  OAI2BB1XL U1452 ( .A0N(n965), .A1N(sa13_next[3]), .B0(n1161), .Y(N67) );
  OAI2BB1XL U1453 ( .A0N(n965), .A1N(sa13_next[2]), .B0(n1159), .Y(N66) );
  OAI2BB1XL U1454 ( .A0N(n965), .A1N(sa23_next[7]), .B0(n1155), .Y(N55) );
  OAI2BB1XL U1455 ( .A0N(n965), .A1N(sa23_next[6]), .B0(n1153), .Y(N54) );
  AOI2BB2XL U1456 ( .B0(w1[1]), .B1(sa31_sr[1]), .A0N(sa31_sr[1]), .A1N(w1[1]), 
        .Y(N486) );
  AOI2BB2XL U1457 ( .B0(w0[9]), .B1(sa20_sr[1]), .A0N(sa20_sr[1]), .A1N(w0[9]), 
        .Y(N446) );
  AOI2BB2XL U1458 ( .B0(w0[25]), .B1(sa00_sr[1]), .A0N(sa00_sr[1]), .A1N(
        w0[25]), .Y(N382) );
  AOI2BB2XL U1459 ( .B0(w1[17]), .B1(sa11_sr[1]), .A0N(sa11_sr[1]), .A1N(
        w1[17]), .Y(N422) );
  AOI2BB2XL U1460 ( .B0(w2[25]), .B1(sa02_sr[1]), .A0N(sa02_sr[1]), .A1N(
        w2[25]), .Y(N398) );
  AOI2BB2XL U1461 ( .B0(w3[1]), .B1(sa33_sr[1]), .A0N(sa33_sr[1]), .A1N(w3[1]), 
        .Y(N502) );
  AOI2BB2XL U1462 ( .B0(w2[9]), .B1(sa22_sr[1]), .A0N(sa22_sr[1]), .A1N(w2[9]), 
        .Y(N462) );
  AOI2BB2XL U1463 ( .B0(w3[25]), .B1(sa03_sr[1]), .A0N(sa03_sr[1]), .A1N(
        w3[25]), .Y(N406) );
  AOI2BB2XL U1464 ( .B0(w3[9]), .B1(sa23_sr[1]), .A0N(sa23_sr[1]), .A1N(w3[9]), 
        .Y(N470) );
  AOI2BB2XL U1465 ( .B0(w2[1]), .B1(sa32_sr[1]), .A0N(sa32_sr[1]), .A1N(w2[1]), 
        .Y(N494) );
  AOI2BB2XL U1466 ( .B0(w0[17]), .B1(sa10_sr[1]), .A0N(sa10_sr[1]), .A1N(
        w0[17]), .Y(N414) );
  AOI2BB2XL U1467 ( .B0(w1[25]), .B1(sa01_sr[1]), .A0N(sa01_sr[1]), .A1N(
        w1[25]), .Y(N390) );
  AOI2BB2XL U1468 ( .B0(w2[17]), .B1(sa12_sr[1]), .A0N(sa12_sr[1]), .A1N(
        w2[17]), .Y(N430) );
  AOI2BB2XL U1469 ( .B0(w3[17]), .B1(sa13_sr[1]), .A0N(sa13_sr[1]), .A1N(
        w3[17]), .Y(N438) );
  AOI2BB2XL U1470 ( .B0(w1[9]), .B1(sa21_sr[1]), .A0N(sa21_sr[1]), .A1N(w1[9]), 
        .Y(N454) );
  AOI2BB2XL U1471 ( .B0(w0[1]), .B1(sa30_sr[1]), .A0N(sa30_sr[1]), .A1N(w0[1]), 
        .Y(N478) );
  AOI2BB2XL U1472 ( .B0(w0[31]), .B1(sa00_sr[7]), .A0N(sa00_sr[7]), .A1N(
        w0[31]), .Y(N376) );
  AOI2BB2XL U1473 ( .B0(w2[20]), .B1(sa12_sr[4]), .A0N(sa12_sr[4]), .A1N(
        w2[20]), .Y(N427) );
  AOI2BB2XL U1474 ( .B0(w2[11]), .B1(sa22_sr[3]), .A0N(sa22_sr[3]), .A1N(
        w2[11]), .Y(N460) );
  AOI2BB2XL U1475 ( .B0(w0[23]), .B1(sa10_sr[7]), .A0N(sa10_sr[7]), .A1N(
        w0[23]), .Y(N408) );
  AOI2BB2XL U1476 ( .B0(w3[4]), .B1(sa33_sr[4]), .A0N(sa33_sr[4]), .A1N(w3[4]), 
        .Y(N499) );
  AOI2BB2XL U1477 ( .B0(w3[19]), .B1(sa13_sr[3]), .A0N(sa13_sr[3]), .A1N(
        w3[19]), .Y(N436) );
  AOI2BB2XL U1478 ( .B0(w1[27]), .B1(sa01_sr[3]), .A0N(sa01_sr[3]), .A1N(
        w1[27]), .Y(N388) );
  AOI2BB2XL U1479 ( .B0(w0[21]), .B1(sa10_sr[5]), .A0N(sa10_sr[5]), .A1N(
        w0[21]), .Y(N410) );
  AOI2BB2XL U1480 ( .B0(w0[30]), .B1(sa00_sr[6]), .A0N(sa00_sr[6]), .A1N(
        w0[30]), .Y(N377) );
  AOI2BB2XL U1481 ( .B0(w3[20]), .B1(sa13_sr[4]), .A0N(sa13_sr[4]), .A1N(
        w3[20]), .Y(N435) );
  AOI2BB2XL U1482 ( .B0(w0[6]), .B1(sa30_sr[6]), .A0N(sa30_sr[6]), .A1N(w0[6]), 
        .Y(N473) );
  AOI2BB2XL U1483 ( .B0(w2[29]), .B1(sa02_sr[5]), .A0N(sa02_sr[5]), .A1N(
        w2[29]), .Y(N394) );
  AOI2BB2XL U1484 ( .B0(w3[23]), .B1(sa13_sr[7]), .A0N(sa13_sr[7]), .A1N(
        w3[23]), .Y(N432) );
  AOI2BB2XL U1485 ( .B0(w0[11]), .B1(sa20_sr[3]), .A0N(sa20_sr[3]), .A1N(
        w0[11]), .Y(N444) );
  AOI2BB2XL U1486 ( .B0(w3[28]), .B1(sa03_sr[4]), .A0N(sa03_sr[4]), .A1N(
        w3[28]), .Y(N403) );
  AOI2BB2XL U1487 ( .B0(w2[10]), .B1(sa22_sr[2]), .A0N(sa22_sr[2]), .A1N(
        w2[10]), .Y(N461) );
  AOI2BB2XL U1488 ( .B0(w3[18]), .B1(sa13_sr[2]), .A0N(sa13_sr[2]), .A1N(
        w3[18]), .Y(N437) );
  AOI2BB2XL U1489 ( .B0(w3[2]), .B1(sa33_sr[2]), .A0N(sa33_sr[2]), .A1N(w3[2]), 
        .Y(N501) );
  AOI2BB2XL U1490 ( .B0(w3[27]), .B1(sa03_sr[3]), .A0N(sa03_sr[3]), .A1N(
        w3[27]), .Y(N404) );
  AOI2BB2XL U1491 ( .B0(w3[22]), .B1(sa13_sr[6]), .A0N(sa13_sr[6]), .A1N(
        w3[22]), .Y(N433) );
  AOI2BB2XL U1492 ( .B0(w2[21]), .B1(sa12_sr[5]), .A0N(sa12_sr[5]), .A1N(
        w2[21]), .Y(N426) );
  AOI2BB2XL U1493 ( .B0(w1[18]), .B1(sa11_sr[2]), .A0N(sa11_sr[2]), .A1N(
        w1[18]), .Y(N421) );
  AOI2BB2XL U1494 ( .B0(w1[28]), .B1(sa01_sr[4]), .A0N(sa01_sr[4]), .A1N(
        w1[28]), .Y(N387) );
  AOI2BB2XL U1495 ( .B0(w2[26]), .B1(sa02_sr[2]), .A0N(sa02_sr[2]), .A1N(
        w2[26]), .Y(N397) );
  AOI2BB2XL U1496 ( .B0(w2[28]), .B1(sa02_sr[4]), .A0N(sa02_sr[4]), .A1N(
        w2[28]), .Y(N395) );
  AOI2BB2XL U1497 ( .B0(w0[14]), .B1(sa20_sr[6]), .A0N(sa20_sr[6]), .A1N(
        w0[14]), .Y(N441) );
  AOI2BB2XL U1498 ( .B0(w1[26]), .B1(sa01_sr[2]), .A0N(sa01_sr[2]), .A1N(
        w1[26]), .Y(N389) );
  AOI2BB2XL U1499 ( .B0(w2[6]), .B1(sa32_sr[6]), .A0N(sa32_sr[6]), .A1N(w2[6]), 
        .Y(N489) );
  AOI2BB2XL U1500 ( .B0(w2[30]), .B1(sa02_sr[6]), .A0N(sa02_sr[6]), .A1N(
        w2[30]), .Y(N393) );
  AOI2BB2XL U1501 ( .B0(w3[21]), .B1(sa13_sr[5]), .A0N(sa13_sr[5]), .A1N(
        w3[21]), .Y(N434) );
  AOI2BB2XL U1502 ( .B0(w2[7]), .B1(sa32_sr[7]), .A0N(sa32_sr[7]), .A1N(w2[7]), 
        .Y(N488) );
  AOI2BB2XL U1503 ( .B0(w3[3]), .B1(sa33_sr[3]), .A0N(sa33_sr[3]), .A1N(w3[3]), 
        .Y(N500) );
  AOI2BB2XL U1504 ( .B0(w3[15]), .B1(sa23_sr[7]), .A0N(sa23_sr[7]), .A1N(
        w3[15]), .Y(N464) );
  AOI2BB2XL U1505 ( .B0(w0[26]), .B1(sa00_sr[2]), .A0N(sa00_sr[2]), .A1N(
        w0[26]), .Y(N381) );
  AOI2BB2XL U1506 ( .B0(w2[22]), .B1(sa12_sr[6]), .A0N(sa12_sr[6]), .A1N(
        w2[22]), .Y(N425) );
  AOI2BB2XL U1507 ( .B0(w3[14]), .B1(sa23_sr[6]), .A0N(sa23_sr[6]), .A1N(
        w3[14]), .Y(N465) );
  AOI2BB2XL U1508 ( .B0(w3[13]), .B1(sa23_sr[5]), .A0N(sa23_sr[5]), .A1N(
        w3[13]), .Y(N466) );
  AOI2BB2XL U1509 ( .B0(w0[13]), .B1(sa20_sr[5]), .A0N(sa20_sr[5]), .A1N(
        w0[13]), .Y(N442) );
  AOI2BB2XL U1510 ( .B0(w2[31]), .B1(sa02_sr[7]), .A0N(sa02_sr[7]), .A1N(
        w2[31]), .Y(N392) );
  AOI2BB2XL U1511 ( .B0(w1[19]), .B1(sa11_sr[3]), .A0N(sa11_sr[3]), .A1N(
        w1[19]), .Y(N420) );
  AOI2BB2XL U1512 ( .B0(w3[12]), .B1(sa23_sr[4]), .A0N(sa23_sr[4]), .A1N(
        w3[12]), .Y(N467) );
  AOI2BB2XL U1513 ( .B0(w2[27]), .B1(sa02_sr[3]), .A0N(sa02_sr[3]), .A1N(
        w2[27]), .Y(N396) );
  AOI2BB2XL U1514 ( .B0(w3[11]), .B1(sa23_sr[3]), .A0N(sa23_sr[3]), .A1N(
        w3[11]), .Y(N468) );
  AOI2BB2XL U1515 ( .B0(w2[2]), .B1(sa32_sr[2]), .A0N(sa32_sr[2]), .A1N(w2[2]), 
        .Y(N493) );
  AOI2BB2XL U1516 ( .B0(w3[5]), .B1(sa33_sr[5]), .A0N(sa33_sr[5]), .A1N(w3[5]), 
        .Y(N498) );
  AOI2BB2XL U1517 ( .B0(w3[10]), .B1(sa23_sr[2]), .A0N(sa23_sr[2]), .A1N(
        w3[10]), .Y(N469) );
  AOI2BB2XL U1518 ( .B0(w3[26]), .B1(sa03_sr[2]), .A0N(sa03_sr[2]), .A1N(
        w3[26]), .Y(N405) );
  AOI2BB2XL U1519 ( .B0(w1[3]), .B1(sa31_sr[3]), .A0N(sa31_sr[3]), .A1N(w1[3]), 
        .Y(N484) );
  AOI2BB2XL U1520 ( .B0(w1[5]), .B1(sa31_sr[5]), .A0N(sa31_sr[5]), .A1N(w1[5]), 
        .Y(N482) );
  AOI2BB2XL U1521 ( .B0(w0[3]), .B1(sa30_sr[3]), .A0N(sa30_sr[3]), .A1N(w0[3]), 
        .Y(N476) );
  AOI2BB2XL U1522 ( .B0(w3[7]), .B1(sa33_sr[7]), .A0N(sa33_sr[7]), .A1N(w3[7]), 
        .Y(N496) );
  AOI2BB2XL U1523 ( .B0(w3[6]), .B1(sa33_sr[6]), .A0N(sa33_sr[6]), .A1N(w3[6]), 
        .Y(N497) );
  AOI2BB2XL U1524 ( .B0(w0[7]), .B1(sa30_sr[7]), .A0N(sa30_sr[7]), .A1N(w0[7]), 
        .Y(N472) );
  AOI2BB2XL U1525 ( .B0(w0[27]), .B1(sa00_sr[3]), .A0N(sa00_sr[3]), .A1N(
        w0[27]), .Y(N380) );
  AOI2BB2XL U1526 ( .B0(w2[3]), .B1(sa32_sr[3]), .A0N(sa32_sr[3]), .A1N(w2[3]), 
        .Y(N492) );
  AOI2BB2XL U1527 ( .B0(w0[18]), .B1(sa10_sr[2]), .A0N(sa10_sr[2]), .A1N(
        w0[18]), .Y(N413) );
  AOI2BB2XL U1528 ( .B0(w1[4]), .B1(sa31_sr[4]), .A0N(sa31_sr[4]), .A1N(w1[4]), 
        .Y(N483) );
  AOI2BB2XL U1529 ( .B0(w0[12]), .B1(sa20_sr[4]), .A0N(sa20_sr[4]), .A1N(
        w0[12]), .Y(N443) );
  AOI2BB2XL U1530 ( .B0(w0[28]), .B1(sa00_sr[4]), .A0N(sa00_sr[4]), .A1N(
        w0[28]), .Y(N379) );
  AOI2BB2XL U1531 ( .B0(w1[15]), .B1(sa21_sr[7]), .A0N(sa21_sr[7]), .A1N(
        w1[15]), .Y(N448) );
  AOI2BB2XL U1532 ( .B0(w1[23]), .B1(sa11_sr[7]), .A0N(sa11_sr[7]), .A1N(
        w1[23]), .Y(N416) );
  AOI2BB2XL U1533 ( .B0(w0[22]), .B1(sa10_sr[6]), .A0N(sa10_sr[6]), .A1N(
        w0[22]), .Y(N409) );
  AOI2BB2XL U1534 ( .B0(w1[31]), .B1(sa01_sr[7]), .A0N(sa01_sr[7]), .A1N(
        w1[31]), .Y(N384) );
  AOI2BB2XL U1535 ( .B0(w2[14]), .B1(sa22_sr[6]), .A0N(sa22_sr[6]), .A1N(
        w2[14]), .Y(N457) );
  AOI2BB2XL U1536 ( .B0(w1[22]), .B1(sa11_sr[6]), .A0N(sa11_sr[6]), .A1N(
        w1[22]), .Y(N417) );
  AOI2BB2XL U1537 ( .B0(w1[13]), .B1(sa21_sr[5]), .A0N(sa21_sr[5]), .A1N(
        w1[13]), .Y(N450) );
  AOI2BB2XL U1538 ( .B0(w0[15]), .B1(sa20_sr[7]), .A0N(sa20_sr[7]), .A1N(
        w0[15]), .Y(N440) );
  AOI2BB2XL U1539 ( .B0(w0[20]), .B1(sa10_sr[4]), .A0N(sa10_sr[4]), .A1N(
        w0[20]), .Y(N411) );
  AOI2BB2XL U1540 ( .B0(w1[11]), .B1(sa21_sr[3]), .A0N(sa21_sr[3]), .A1N(
        w1[11]), .Y(N452) );
  AOI2BB2XL U1541 ( .B0(w2[23]), .B1(sa12_sr[7]), .A0N(sa12_sr[7]), .A1N(
        w2[23]), .Y(N424) );
  AOI2BB2XL U1542 ( .B0(w2[13]), .B1(sa22_sr[5]), .A0N(sa22_sr[5]), .A1N(
        w2[13]), .Y(N458) );
  AOI2BB2XL U1543 ( .B0(w1[30]), .B1(sa01_sr[6]), .A0N(sa01_sr[6]), .A1N(
        w1[30]), .Y(N385) );
  AOI2BB2XL U1544 ( .B0(w2[4]), .B1(sa32_sr[4]), .A0N(sa32_sr[4]), .A1N(w2[4]), 
        .Y(N491) );
  AOI2BB2XL U1545 ( .B0(w1[2]), .B1(sa31_sr[2]), .A0N(sa31_sr[2]), .A1N(w1[2]), 
        .Y(N485) );
  AOI2BB2XL U1546 ( .B0(w1[10]), .B1(sa21_sr[2]), .A0N(sa21_sr[2]), .A1N(
        w1[10]), .Y(N453) );
  AOI2BB2XL U1547 ( .B0(w0[10]), .B1(sa20_sr[2]), .A0N(sa20_sr[2]), .A1N(
        w0[10]), .Y(N445) );
  AOI2BB2XL U1548 ( .B0(w1[7]), .B1(sa31_sr[7]), .A0N(sa31_sr[7]), .A1N(w1[7]), 
        .Y(N480) );
  AOI2BB2XL U1549 ( .B0(w3[29]), .B1(sa03_sr[5]), .A0N(sa03_sr[5]), .A1N(
        w3[29]), .Y(N402) );
  AOI2BB2XL U1550 ( .B0(w1[20]), .B1(sa11_sr[4]), .A0N(sa11_sr[4]), .A1N(
        w1[20]), .Y(N419) );
  AOI2BB2XL U1551 ( .B0(w0[5]), .B1(sa30_sr[5]), .A0N(sa30_sr[5]), .A1N(w0[5]), 
        .Y(N474) );
  AOI2BB2XL U1552 ( .B0(w2[15]), .B1(sa22_sr[7]), .A0N(sa22_sr[7]), .A1N(
        w2[15]), .Y(N456) );
  AOI2BB2XL U1553 ( .B0(w1[12]), .B1(sa21_sr[4]), .A0N(sa21_sr[4]), .A1N(
        w1[12]), .Y(N451) );
  AOI2BB2XL U1554 ( .B0(w0[29]), .B1(sa00_sr[5]), .A0N(sa00_sr[5]), .A1N(
        w0[29]), .Y(N378) );
  AOI2BB2XL U1555 ( .B0(w0[2]), .B1(sa30_sr[2]), .A0N(sa30_sr[2]), .A1N(w0[2]), 
        .Y(N477) );
  AOI2BB2XL U1556 ( .B0(w1[14]), .B1(sa21_sr[6]), .A0N(sa21_sr[6]), .A1N(
        w1[14]), .Y(N449) );
  AOI2BB2XL U1557 ( .B0(w1[29]), .B1(sa01_sr[5]), .A0N(sa01_sr[5]), .A1N(
        w1[29]), .Y(N386) );
  AOI2BB2XL U1558 ( .B0(w1[6]), .B1(sa31_sr[6]), .A0N(sa31_sr[6]), .A1N(w1[6]), 
        .Y(N481) );
  AOI2BB2XL U1559 ( .B0(w0[4]), .B1(sa30_sr[4]), .A0N(sa30_sr[4]), .A1N(w0[4]), 
        .Y(N475) );
  AOI2BB2XL U1560 ( .B0(w2[18]), .B1(sa12_sr[2]), .A0N(sa12_sr[2]), .A1N(
        w2[18]), .Y(N429) );
  AOI2BB2XL U1561 ( .B0(w2[19]), .B1(sa12_sr[3]), .A0N(sa12_sr[3]), .A1N(
        w2[19]), .Y(N428) );
  AOI2BB2XL U1562 ( .B0(w3[30]), .B1(sa03_sr[6]), .A0N(sa03_sr[6]), .A1N(
        w3[30]), .Y(N401) );
  AOI2BB2XL U1563 ( .B0(w2[12]), .B1(sa22_sr[4]), .A0N(sa22_sr[4]), .A1N(
        w2[12]), .Y(N459) );
  AOI2BB2XL U1564 ( .B0(w1[21]), .B1(sa11_sr[5]), .A0N(sa11_sr[5]), .A1N(
        w1[21]), .Y(N418) );
  AOI2BB2XL U1565 ( .B0(w0[19]), .B1(sa10_sr[3]), .A0N(sa10_sr[3]), .A1N(
        w0[19]), .Y(N412) );
  AOI2BB2XL U1566 ( .B0(w3[31]), .B1(sa03_sr[7]), .A0N(sa03_sr[7]), .A1N(
        w3[31]), .Y(N400) );
  AOI2BB2XL U1567 ( .B0(w2[5]), .B1(sa32_sr[5]), .A0N(sa32_sr[5]), .A1N(w2[5]), 
        .Y(N490) );
  AOI2BB2XL U1568 ( .B0(w0[8]), .B1(sa20_sr[0]), .A0N(sa20_sr[0]), .A1N(w0[8]), 
        .Y(N447) );
  AOI2BB2XL U1569 ( .B0(w2[16]), .B1(sa12_sr[0]), .A0N(sa12_sr[0]), .A1N(
        w2[16]), .Y(N431) );
  AOI2BB2XL U1570 ( .B0(w3[16]), .B1(sa13_sr[0]), .A0N(sa13_sr[0]), .A1N(
        w3[16]), .Y(N439) );
  AOI2BB2XL U1571 ( .B0(w0[0]), .B1(sa30_sr[0]), .A0N(sa30_sr[0]), .A1N(w0[0]), 
        .Y(N479) );
  AOI2BB2XL U1572 ( .B0(w1[16]), .B1(sa11_sr[0]), .A0N(sa11_sr[0]), .A1N(
        w1[16]), .Y(N423) );
  AOI2BB2XL U1573 ( .B0(w2[24]), .B1(sa02_sr[0]), .A0N(sa02_sr[0]), .A1N(
        w2[24]), .Y(N399) );
  AOI2BB2XL U1574 ( .B0(w3[0]), .B1(sa33_sr[0]), .A0N(sa33_sr[0]), .A1N(w3[0]), 
        .Y(N503) );
  AOI2BB2XL U1575 ( .B0(w1[24]), .B1(sa01_sr[0]), .A0N(sa01_sr[0]), .A1N(
        w1[24]), .Y(N391) );
  AOI2BB2XL U1576 ( .B0(w0[24]), .B1(sa00_sr[0]), .A0N(sa00_sr[0]), .A1N(
        w0[24]), .Y(N383) );
  AOI2BB2XL U1577 ( .B0(w1[0]), .B1(sa31_sr[0]), .A0N(sa31_sr[0]), .A1N(w1[0]), 
        .Y(N487) );
  AOI2BB2XL U1578 ( .B0(w3[8]), .B1(sa23_sr[0]), .A0N(sa23_sr[0]), .A1N(w3[8]), 
        .Y(N471) );
  AOI2BB2XL U1579 ( .B0(w0[16]), .B1(sa10_sr[0]), .A0N(sa10_sr[0]), .A1N(
        w0[16]), .Y(N415) );
  AOI2BB2XL U1580 ( .B0(w2[0]), .B1(sa32_sr[0]), .A0N(sa32_sr[0]), .A1N(w2[0]), 
        .Y(N495) );
  AOI2BB2XL U1581 ( .B0(w2[8]), .B1(sa22_sr[0]), .A0N(sa22_sr[0]), .A1N(w2[8]), 
        .Y(N463) );
  AOI2BB2XL U1582 ( .B0(w3[24]), .B1(sa03_sr[0]), .A0N(sa03_sr[0]), .A1N(
        w3[24]), .Y(N407) );
  AOI2BB2XL U1583 ( .B0(w1[8]), .B1(sa21_sr[0]), .A0N(sa21_sr[0]), .A1N(w1[8]), 
        .Y(N455) );
  OAI2BB1XL U1584 ( .A0N(n1192), .A1N(n1188), .B0(n139), .Y(n399) );
  NAND2XL U1585 ( .A(n1192), .B(n959), .Y(n137) );
  NOR2BXL U1586 ( .AN(n1192), .B(n1191), .Y(n398) );
  NOR3XL U1587 ( .A(dcnt_2_), .B(n959), .C(n1057), .Y(N21) );
  NAND3XL U1588 ( .A(n3), .B(n2), .C(n966), .Y(n1057) );
  CLKINVX3 U1589 ( .A(n960), .Y(n964) );
  AOI21XL U1590 ( .A0(n1190), .A1(dcnt_2_), .B0(n1189), .Y(n1191) );
  AOI21XL U1591 ( .A0(text_in_r[18]), .A1(w3[18]), .B0(n964), .Y(n1158) );
  AOI21XL U1592 ( .A0(w2[18]), .A1(text_in_r[50]), .B0(n4), .Y(n991) );
  AOI21XL U1593 ( .A0(w0[18]), .A1(text_in_r[114]), .B0(n961), .Y(n1100) );
  AOI21XL U1594 ( .A0(w1[18]), .A1(text_in_r[82]), .B0(n963), .Y(n1043) );
  AOI21XL U1595 ( .A0(w0[24]), .A1(text_in_r[120]), .B0(n961), .Y(n1112) );
  AOI21XL U1596 ( .A0(text_in_r[24]), .A1(w3[24]), .B0(n964), .Y(n1170) );
  AOI21XL U1597 ( .A0(w3[7]), .A1(text_in_r[7]), .B0(n962), .Y(n1138) );
  AOI21XL U1598 ( .A0(w1[7]), .A1(text_in_r[71]), .B0(n4), .Y(n1027) );
  AOI21XL U1599 ( .A0(w0[7]), .A1(text_in_r[103]), .B0(n962), .Y(n1080) );
  AOI21XL U1600 ( .A0(w2[7]), .A1(text_in_r[39]), .B0(n965), .Y(n973) );
  AOI21XL U1601 ( .A0(w0[16]), .A1(text_in_r[112]), .B0(n961), .Y(n1096) );
  AOI21XL U1602 ( .A0(w3[3]), .A1(text_in_r[3]), .B0(n962), .Y(n1130) );
  AOI21XL U1603 ( .A0(w1[3]), .A1(text_in_r[67]), .B0(n961), .Y(n1021) );
  AOI21XL U1604 ( .A0(text_in_r[21]), .A1(w3[21]), .B0(n964), .Y(n1164) );
  AOI21XL U1605 ( .A0(w1[21]), .A1(text_in_r[85]), .B0(n963), .Y(n1049) );
  AOI21XL U1606 ( .A0(w0[21]), .A1(text_in_r[117]), .B0(n4), .Y(n1106) );
  AOI21XL U1607 ( .A0(w2[21]), .A1(text_in_r[53]), .B0(n4), .Y(n997) );
  AOI21XL U1608 ( .A0(w3[0]), .A1(text_in_r[0]), .B0(n961), .Y(n1124) );
  AOI21XL U1609 ( .A0(w0[0]), .A1(text_in_r[96]), .B0(n962), .Y(n1068) );
  AOI21XL U1610 ( .A0(text_in_r[19]), .A1(w3[19]), .B0(n964), .Y(n1160) );
  AOI21XL U1611 ( .A0(w2[19]), .A1(text_in_r[51]), .B0(n964), .Y(n993) );
  AOI21XL U1612 ( .A0(w1[19]), .A1(text_in_r[83]), .B0(n4), .Y(n1045) );
  AOI21XL U1613 ( .A0(w0[19]), .A1(text_in_r[115]), .B0(n961), .Y(n1102) );
  AOI21XL U1614 ( .A0(w0[23]), .A1(text_in_r[119]), .B0(n961), .Y(n1110) );
  AOI21XL U1615 ( .A0(w0[8]), .A1(text_in_r[104]), .B0(n962), .Y(n1082) );
  AOI21XL U1616 ( .A0(w0[2]), .A1(text_in_r[98]), .B0(n962), .Y(n1072) );
  AOI21XL U1617 ( .A0(w3[2]), .A1(text_in_r[2]), .B0(n962), .Y(n1128) );
  AOI21XL U1618 ( .A0(w1[2]), .A1(text_in_r[66]), .B0(n965), .Y(n1019) );
  AOI21XL U1619 ( .A0(text_in_r[34]), .A1(w2[2]), .B0(n964), .Y(n1184) );
  AOI21XL U1620 ( .A0(w2[23]), .A1(text_in_r[55]), .B0(n964), .Y(n1001) );
  AOI21XL U1621 ( .A0(text_in_r[23]), .A1(w3[23]), .B0(n965), .Y(n1168) );
  AOI21XL U1622 ( .A0(w1[23]), .A1(text_in_r[87]), .B0(n963), .Y(n1053) );
  AOI21XL U1623 ( .A0(text_in_r[8]), .A1(w3[8]), .B0(n962), .Y(n1140) );
  AOI21XL U1624 ( .A0(text_in_r[11]), .A1(w3[11]), .B0(n963), .Y(n1146) );
  AOI21XL U1625 ( .A0(w0[11]), .A1(text_in_r[107]), .B0(n961), .Y(n1088) );
  AOI21XL U1626 ( .A0(text_in_r[14]), .A1(w3[14]), .B0(n963), .Y(n1152) );
  AOI21XL U1627 ( .A0(w1[11]), .A1(text_in_r[75]), .B0(n963), .Y(n1033) );
  AOI21XL U1628 ( .A0(w2[11]), .A1(text_in_r[43]), .B0(n4), .Y(n979) );
  AOI21XL U1629 ( .A0(w1[31]), .A1(text_in_r[95]), .B0(n962), .Y(n1066) );
  AOI21XL U1630 ( .A0(text_in_r[31]), .A1(w3[31]), .B0(n964), .Y(n1180) );
  AOI21XL U1631 ( .A0(w2[31]), .A1(text_in_r[63]), .B0(n963), .Y(n1015) );
  AOI21XL U1632 ( .A0(w0[31]), .A1(text_in_r[127]), .B0(n961), .Y(n1122) );
  AOI21XL U1633 ( .A0(w1[6]), .A1(text_in_r[70]), .B0(n4), .Y(n1025) );
  AOI21XL U1634 ( .A0(w1[14]), .A1(text_in_r[78]), .B0(n963), .Y(n1037) );
  AOI21XL U1635 ( .A0(w2[6]), .A1(text_in_r[38]), .B0(n964), .Y(n971) );
  AOI21XL U1636 ( .A0(w2[14]), .A1(text_in_r[46]), .B0(n964), .Y(n985) );
  AOI21XL U1637 ( .A0(w0[14]), .A1(text_in_r[110]), .B0(n961), .Y(n1092) );
  AOI21XL U1638 ( .A0(w0[6]), .A1(text_in_r[102]), .B0(n962), .Y(n1078) );
  AOI21XL U1639 ( .A0(w3[6]), .A1(text_in_r[6]), .B0(n962), .Y(n1136) );
  AOI21XL U1640 ( .A0(w0[5]), .A1(text_in_r[101]), .B0(n962), .Y(n1076) );
  AOI21XL U1641 ( .A0(w2[5]), .A1(text_in_r[37]), .B0(n965), .Y(n969) );
  AOI21XL U1642 ( .A0(w3[5]), .A1(text_in_r[5]), .B0(n962), .Y(n1134) );
  AOI21XL U1643 ( .A0(w1[5]), .A1(text_in_r[69]), .B0(n4), .Y(n1023) );
  AOI21XL U1644 ( .A0(w2[27]), .A1(text_in_r[59]), .B0(n962), .Y(n1007) );
  AOI21XL U1645 ( .A0(w0[27]), .A1(text_in_r[123]), .B0(n961), .Y(n1116) );
  AOI21XL U1646 ( .A0(w1[27]), .A1(text_in_r[91]), .B0(n962), .Y(n1060) );
  AOI21XL U1647 ( .A0(text_in_r[27]), .A1(w3[27]), .B0(n964), .Y(n1176) );
  AOI21XL U1648 ( .A0(text_in_r[33]), .A1(w2[1]), .B0(n965), .Y(n1182) );
  AOI21XL U1649 ( .A0(w0[1]), .A1(text_in_r[97]), .B0(n962), .Y(n1070) );
  AOI21XL U1650 ( .A0(w3[1]), .A1(text_in_r[1]), .B0(n961), .Y(n1126) );
  AOI21XL U1651 ( .A0(w1[1]), .A1(text_in_r[65]), .B0(n964), .Y(n1017) );
  AOI21XL U1652 ( .A0(w2[17]), .A1(text_in_r[49]), .B0(n964), .Y(n989) );
  AOI21XL U1653 ( .A0(text_in_r[17]), .A1(w3[17]), .B0(n963), .Y(n1156) );
  AOI21XL U1654 ( .A0(w1[17]), .A1(text_in_r[81]), .B0(n963), .Y(n1041) );
  AOI21XL U1655 ( .A0(w0[17]), .A1(text_in_r[113]), .B0(n961), .Y(n1098) );
  AOI21XL U1656 ( .A0(text_in_r[15]), .A1(w3[15]), .B0(n963), .Y(n1154) );
  AOI21XL U1657 ( .A0(w0[15]), .A1(text_in_r[111]), .B0(n961), .Y(n1094) );
  AOI21XL U1658 ( .A0(w2[15]), .A1(text_in_r[47]), .B0(n964), .Y(n987) );
  AOI21XL U1659 ( .A0(w1[15]), .A1(text_in_r[79]), .B0(n963), .Y(n1039) );
  AOI21XL U1660 ( .A0(w2[30]), .A1(text_in_r[62]), .B0(n961), .Y(n1013) );
  AOI21XL U1661 ( .A0(w3[4]), .A1(text_in_r[4]), .B0(n962), .Y(n1132) );
  AOI21XL U1662 ( .A0(w2[4]), .A1(text_in_r[36]), .B0(n961), .Y(n967) );
  AOI21XL U1663 ( .A0(w0[4]), .A1(text_in_r[100]), .B0(n962), .Y(n1074) );
  AOI21XL U1664 ( .A0(text_in_r[22]), .A1(w3[22]), .B0(n964), .Y(n1166) );
  AOI21XL U1665 ( .A0(w2[9]), .A1(text_in_r[41]), .B0(n964), .Y(n975) );
  AOI21XL U1666 ( .A0(text_in_r[9]), .A1(w3[9]), .B0(n962), .Y(n1142) );
  AOI21XL U1667 ( .A0(w0[9]), .A1(text_in_r[105]), .B0(n962), .Y(n1084) );
  AOI21XL U1668 ( .A0(w1[9]), .A1(text_in_r[73]), .B0(n4), .Y(n1029) );
  AOI21XL U1669 ( .A0(w1[22]), .A1(text_in_r[86]), .B0(n963), .Y(n1051) );
  AOI21XL U1670 ( .A0(w0[22]), .A1(text_in_r[118]), .B0(n961), .Y(n1108) );
  AOI21XL U1671 ( .A0(w2[22]), .A1(text_in_r[54]), .B0(n964), .Y(n999) );
  AOI21XL U1672 ( .A0(w2[26]), .A1(text_in_r[58]), .B0(n4), .Y(n1005) );
  AOI21XL U1673 ( .A0(text_in_r[26]), .A1(w3[26]), .B0(n964), .Y(n1174) );
  AOI21XL U1674 ( .A0(w1[26]), .A1(text_in_r[90]), .B0(n962), .Y(n1058) );
  AOI21XL U1675 ( .A0(text_in_r[10]), .A1(w3[10]), .B0(n963), .Y(n1144) );
  AOI21XL U1676 ( .A0(w1[10]), .A1(text_in_r[74]), .B0(n963), .Y(n1031) );
  AOI21XL U1677 ( .A0(w2[10]), .A1(text_in_r[42]), .B0(n965), .Y(n977) );
  AOI21XL U1678 ( .A0(w0[10]), .A1(text_in_r[106]), .B0(n961), .Y(n1086) );
  AOI21XL U1679 ( .A0(text_in_r[25]), .A1(w3[25]), .B0(n964), .Y(n1172) );
  AOI21XL U1680 ( .A0(w0[25]), .A1(text_in_r[121]), .B0(n4), .Y(n1114) );
  AOI21XL U1681 ( .A0(w2[25]), .A1(text_in_r[57]), .B0(n4), .Y(n1003) );
  AOI21XL U1682 ( .A0(w1[25]), .A1(text_in_r[89]), .B0(n963), .Y(n1055) );
  AOI21XL U1683 ( .A0(w2[29]), .A1(text_in_r[61]), .B0(n962), .Y(n1011) );
  AOI21XL U1684 ( .A0(w0[29]), .A1(text_in_r[125]), .B0(n961), .Y(n1120) );
  AOI21XL U1685 ( .A0(w1[29]), .A1(text_in_r[93]), .B0(n962), .Y(n1064) );
  AOI21XL U1686 ( .A0(text_in_r[20]), .A1(w3[20]), .B0(n964), .Y(n1162) );
  AOI21XL U1687 ( .A0(w1[20]), .A1(text_in_r[84]), .B0(n963), .Y(n1047) );
  AOI21XL U1688 ( .A0(w0[20]), .A1(text_in_r[116]), .B0(n961), .Y(n1104) );
  AOI21XL U1689 ( .A0(w2[20]), .A1(text_in_r[52]), .B0(n964), .Y(n995) );
  AOI21XL U1690 ( .A0(text_in_r[12]), .A1(w3[12]), .B0(n963), .Y(n1148) );
  AOI21XL U1691 ( .A0(w1[12]), .A1(text_in_r[76]), .B0(n963), .Y(n1035) );
  AOI21XL U1692 ( .A0(w0[12]), .A1(text_in_r[108]), .B0(n961), .Y(n1090) );
  AOI21XL U1693 ( .A0(w2[12]), .A1(text_in_r[44]), .B0(n4), .Y(n981) );
  AOI21XL U1694 ( .A0(text_in_r[13]), .A1(w3[13]), .B0(n963), .Y(n1150) );
  CLKINVX3 U1695 ( .A(n960), .Y(n963) );
  AOI21XL U1696 ( .A0(w2[13]), .A1(text_in_r[45]), .B0(n965), .Y(n983) );
  AOI21XL U1697 ( .A0(w2[28]), .A1(text_in_r[60]), .B0(n965), .Y(n1009) );
  AOI21XL U1698 ( .A0(w1[28]), .A1(text_in_r[92]), .B0(n962), .Y(n1062) );
  CLKINVX3 U1699 ( .A(n960), .Y(n962) );
  AOI21XL U1700 ( .A0(w0[28]), .A1(text_in_r[124]), .B0(n961), .Y(n1118) );
  CLKINVX3 U1701 ( .A(n960), .Y(n961) );
  AOI21XL U1702 ( .A0(text_in_r[28]), .A1(w3[28]), .B0(n964), .Y(n1178) );
  INVX1 U1703 ( .A(ld), .Y(n966) );
  OAI21XL U1704 ( .A0(w2[4]), .A1(text_in_r[36]), .B0(n967), .Y(n968) );
  OAI21XL U1705 ( .A0(w2[5]), .A1(text_in_r[37]), .B0(n969), .Y(n970) );
  OAI21XL U1706 ( .A0(w2[6]), .A1(text_in_r[38]), .B0(n971), .Y(n972) );
  OAI2BB1X1 U1707 ( .A0N(n4), .A1N(sa32_next[6]), .B0(n972), .Y(N102) );
  OAI21XL U1708 ( .A0(w2[7]), .A1(text_in_r[39]), .B0(n973), .Y(n974) );
  OAI21XL U1709 ( .A0(w2[9]), .A1(text_in_r[41]), .B0(n975), .Y(n976) );
  OAI21XL U1710 ( .A0(w2[10]), .A1(text_in_r[42]), .B0(n977), .Y(n978) );
  OAI21XL U1711 ( .A0(w2[11]), .A1(text_in_r[43]), .B0(n979), .Y(n980) );
  OAI21XL U1712 ( .A0(w2[12]), .A1(text_in_r[44]), .B0(n981), .Y(n982) );
  OAI21XL U1713 ( .A0(w2[13]), .A1(text_in_r[45]), .B0(n983), .Y(n984) );
  OAI21XL U1714 ( .A0(w2[14]), .A1(text_in_r[46]), .B0(n985), .Y(n986) );
  OAI2BB1X1 U1715 ( .A0N(n4), .A1N(sa22_next[6]), .B0(n986), .Y(N118) );
  OAI21XL U1716 ( .A0(w2[15]), .A1(text_in_r[47]), .B0(n987), .Y(n988) );
  OAI21XL U1717 ( .A0(w2[17]), .A1(text_in_r[49]), .B0(n989), .Y(n990) );
  OAI21XL U1718 ( .A0(w2[18]), .A1(text_in_r[50]), .B0(n991), .Y(n992) );
  OAI2BB1X1 U1719 ( .A0N(n4), .A1N(sa12_next[2]), .B0(n992), .Y(N130) );
  OAI21XL U1720 ( .A0(w2[19]), .A1(text_in_r[51]), .B0(n993), .Y(n994) );
  OAI21XL U1721 ( .A0(w2[20]), .A1(text_in_r[52]), .B0(n995), .Y(n996) );
  OAI21XL U1722 ( .A0(w2[21]), .A1(text_in_r[53]), .B0(n997), .Y(n998) );
  OAI2BB1X1 U1723 ( .A0N(n4), .A1N(sa12_next[5]), .B0(n998), .Y(N133) );
  OAI21XL U1724 ( .A0(w2[22]), .A1(text_in_r[54]), .B0(n999), .Y(n1000) );
  OAI21XL U1725 ( .A0(w2[23]), .A1(text_in_r[55]), .B0(n1001), .Y(n1002) );
  OAI21XL U1726 ( .A0(w2[25]), .A1(text_in_r[57]), .B0(n1003), .Y(n1004) );
  OAI21XL U1727 ( .A0(w2[26]), .A1(text_in_r[58]), .B0(n1005), .Y(n1006) );
  OAI21XL U1728 ( .A0(w2[27]), .A1(text_in_r[59]), .B0(n1007), .Y(n1008) );
  OAI21XL U1729 ( .A0(w2[28]), .A1(text_in_r[60]), .B0(n1009), .Y(n1010) );
  OAI21XL U1730 ( .A0(w2[29]), .A1(text_in_r[61]), .B0(n1011), .Y(n1012) );
  OAI21XL U1731 ( .A0(w2[30]), .A1(text_in_r[62]), .B0(n1013), .Y(n1014) );
  OAI21XL U1732 ( .A0(w2[31]), .A1(text_in_r[63]), .B0(n1015), .Y(n1016) );
  OAI21XL U1733 ( .A0(w1[1]), .A1(text_in_r[65]), .B0(n1017), .Y(n1018) );
  OAI21XL U1734 ( .A0(w1[2]), .A1(text_in_r[66]), .B0(n1019), .Y(n1020) );
  OAI21XL U1735 ( .A0(w1[3]), .A1(text_in_r[67]), .B0(n1021), .Y(n1022) );
  OAI21XL U1736 ( .A0(w1[5]), .A1(text_in_r[69]), .B0(n1023), .Y(n1024) );
  OAI21XL U1737 ( .A0(w1[6]), .A1(text_in_r[70]), .B0(n1025), .Y(n1026) );
  OAI21XL U1738 ( .A0(w1[7]), .A1(text_in_r[71]), .B0(n1027), .Y(n1028) );
  OAI21XL U1739 ( .A0(w1[9]), .A1(text_in_r[73]), .B0(n1029), .Y(n1030) );
  OAI21XL U1740 ( .A0(w1[10]), .A1(text_in_r[74]), .B0(n1031), .Y(n1032) );
  OAI21XL U1741 ( .A0(w1[11]), .A1(text_in_r[75]), .B0(n1033), .Y(n1034) );
  OAI21XL U1742 ( .A0(w1[12]), .A1(text_in_r[76]), .B0(n1035), .Y(n1036) );
  OAI21XL U1743 ( .A0(w1[14]), .A1(text_in_r[78]), .B0(n1037), .Y(n1038) );
  OAI21XL U1744 ( .A0(w1[15]), .A1(text_in_r[79]), .B0(n1039), .Y(n1040) );
  OAI21XL U1745 ( .A0(w1[17]), .A1(text_in_r[81]), .B0(n1041), .Y(n1042) );
  OAI21XL U1746 ( .A0(w1[18]), .A1(text_in_r[82]), .B0(n1043), .Y(n1044) );
  OAI21XL U1747 ( .A0(w1[19]), .A1(text_in_r[83]), .B0(n1045), .Y(n1046) );
  OAI21XL U1748 ( .A0(w1[20]), .A1(text_in_r[84]), .B0(n1047), .Y(n1048) );
  OAI21XL U1749 ( .A0(w1[21]), .A1(text_in_r[85]), .B0(n1049), .Y(n1050) );
  OAI21XL U1750 ( .A0(w1[22]), .A1(text_in_r[86]), .B0(n1051), .Y(n1052) );
  OAI21XL U1751 ( .A0(w1[23]), .A1(text_in_r[87]), .B0(n1053), .Y(n1054) );
  OAI21XL U1752 ( .A0(w1[25]), .A1(text_in_r[89]), .B0(n1055), .Y(n1056) );
  OAI21XL U1753 ( .A0(w1[26]), .A1(text_in_r[90]), .B0(n1058), .Y(n1059) );
  OAI21XL U1754 ( .A0(w1[27]), .A1(text_in_r[91]), .B0(n1060), .Y(n1061) );
  OAI21XL U1755 ( .A0(w1[28]), .A1(text_in_r[92]), .B0(n1062), .Y(n1063) );
  OAI21XL U1756 ( .A0(w1[29]), .A1(text_in_r[93]), .B0(n1064), .Y(n1065) );
  OAI21XL U1757 ( .A0(w1[31]), .A1(text_in_r[95]), .B0(n1066), .Y(n1067) );
  OAI21XL U1758 ( .A0(w0[0]), .A1(text_in_r[96]), .B0(n1068), .Y(n1069) );
  OAI21XL U1759 ( .A0(w0[1]), .A1(text_in_r[97]), .B0(n1070), .Y(n1071) );
  OAI21XL U1760 ( .A0(w0[2]), .A1(text_in_r[98]), .B0(n1072), .Y(n1073) );
  OAI21XL U1761 ( .A0(w0[4]), .A1(text_in_r[100]), .B0(n1074), .Y(n1075) );
  OAI21XL U1762 ( .A0(w0[5]), .A1(text_in_r[101]), .B0(n1076), .Y(n1077) );
  OAI21XL U1763 ( .A0(w0[6]), .A1(text_in_r[102]), .B0(n1078), .Y(n1079) );
  OAI21XL U1764 ( .A0(w0[7]), .A1(text_in_r[103]), .B0(n1080), .Y(n1081) );
  OAI21XL U1765 ( .A0(w0[8]), .A1(text_in_r[104]), .B0(n1082), .Y(n1083) );
  OAI21XL U1766 ( .A0(w0[9]), .A1(text_in_r[105]), .B0(n1084), .Y(n1085) );
  OAI21XL U1767 ( .A0(w0[10]), .A1(text_in_r[106]), .B0(n1086), .Y(n1087) );
  OAI21XL U1768 ( .A0(w0[11]), .A1(text_in_r[107]), .B0(n1088), .Y(n1089) );
  OAI21XL U1769 ( .A0(w0[12]), .A1(text_in_r[108]), .B0(n1090), .Y(n1091) );
  OAI21XL U1770 ( .A0(w0[14]), .A1(text_in_r[110]), .B0(n1092), .Y(n1093) );
  OAI21XL U1771 ( .A0(w0[15]), .A1(text_in_r[111]), .B0(n1094), .Y(n1095) );
  OAI21XL U1772 ( .A0(w0[16]), .A1(text_in_r[112]), .B0(n1096), .Y(n1097) );
  OAI21XL U1773 ( .A0(w0[17]), .A1(text_in_r[113]), .B0(n1098), .Y(n1099) );
  OAI21XL U1774 ( .A0(w0[18]), .A1(text_in_r[114]), .B0(n1100), .Y(n1101) );
  OAI2BB1X1 U1775 ( .A0N(n4), .A1N(sa10_next[2]), .B0(n1101), .Y(N258) );
  OAI21XL U1776 ( .A0(w0[19]), .A1(text_in_r[115]), .B0(n1102), .Y(n1103) );
  OAI21XL U1777 ( .A0(w0[20]), .A1(text_in_r[116]), .B0(n1104), .Y(n1105) );
  OAI21XL U1778 ( .A0(w0[21]), .A1(text_in_r[117]), .B0(n1106), .Y(n1107) );
  OAI21XL U1779 ( .A0(w0[22]), .A1(text_in_r[118]), .B0(n1108), .Y(n1109) );
  OAI2BB1X1 U1780 ( .A0N(n4), .A1N(sa10_next[6]), .B0(n1109), .Y(N262) );
  OAI21XL U1781 ( .A0(w0[23]), .A1(text_in_r[119]), .B0(n1110), .Y(n1111) );
  OAI21XL U1782 ( .A0(w0[24]), .A1(text_in_r[120]), .B0(n1112), .Y(n1113) );
  OAI21XL U1783 ( .A0(w0[25]), .A1(text_in_r[121]), .B0(n1114), .Y(n1115) );
  OAI21XL U1784 ( .A0(w0[27]), .A1(text_in_r[123]), .B0(n1116), .Y(n1117) );
  OAI21XL U1785 ( .A0(w0[28]), .A1(text_in_r[124]), .B0(n1118), .Y(n1119) );
  OAI21XL U1786 ( .A0(w0[29]), .A1(text_in_r[125]), .B0(n1120), .Y(n1121) );
  OAI21XL U1787 ( .A0(w0[31]), .A1(text_in_r[127]), .B0(n1122), .Y(n1123) );
  OAI21XL U1788 ( .A0(w3[0]), .A1(text_in_r[0]), .B0(n1124), .Y(n1125) );
  OAI2BB1X1 U1789 ( .A0N(n4), .A1N(sa33_next[0]), .B0(n1125), .Y(N32) );
  OAI21XL U1790 ( .A0(w3[1]), .A1(text_in_r[1]), .B0(n1126), .Y(n1127) );
  OAI2BB1X1 U1791 ( .A0N(n4), .A1N(sa33_next[1]), .B0(n1127), .Y(N33) );
  OAI21XL U1792 ( .A0(w3[2]), .A1(text_in_r[2]), .B0(n1128), .Y(n1129) );
  OAI21XL U1793 ( .A0(w3[3]), .A1(text_in_r[3]), .B0(n1130), .Y(n1131) );
  OAI2BB1X1 U1794 ( .A0N(n4), .A1N(sa33_next[3]), .B0(n1131), .Y(N35) );
  OAI21XL U1795 ( .A0(w3[4]), .A1(text_in_r[4]), .B0(n1132), .Y(n1133) );
  OAI2BB1X1 U1796 ( .A0N(n4), .A1N(sa33_next[4]), .B0(n1133), .Y(N36) );
  OAI21XL U1797 ( .A0(w3[5]), .A1(text_in_r[5]), .B0(n1134), .Y(n1135) );
  OAI2BB1X1 U1798 ( .A0N(n4), .A1N(sa33_next[5]), .B0(n1135), .Y(N37) );
  OAI21XL U1799 ( .A0(w3[6]), .A1(text_in_r[6]), .B0(n1136), .Y(n1137) );
  OAI2BB1X1 U1800 ( .A0N(n4), .A1N(sa33_next[6]), .B0(n1137), .Y(N38) );
  OAI21XL U1801 ( .A0(w3[7]), .A1(text_in_r[7]), .B0(n1138), .Y(n1139) );
  OAI2BB1X1 U1802 ( .A0N(n4), .A1N(sa33_next[7]), .B0(n1139), .Y(N39) );
  OAI21XL U1803 ( .A0(text_in_r[8]), .A1(w3[8]), .B0(n1140), .Y(n1141) );
  OAI21XL U1804 ( .A0(text_in_r[9]), .A1(w3[9]), .B0(n1142), .Y(n1143) );
  OAI21XL U1805 ( .A0(text_in_r[10]), .A1(w3[10]), .B0(n1144), .Y(n1145) );
  OAI21XL U1806 ( .A0(text_in_r[11]), .A1(w3[11]), .B0(n1146), .Y(n1147) );
  OAI21XL U1807 ( .A0(text_in_r[12]), .A1(w3[12]), .B0(n1148), .Y(n1149) );
  OAI21XL U1808 ( .A0(text_in_r[13]), .A1(w3[13]), .B0(n1150), .Y(n1151) );
  OAI2BB1X1 U1809 ( .A0N(n4), .A1N(sa23_next[5]), .B0(n1151), .Y(N53) );
  OAI21XL U1810 ( .A0(text_in_r[14]), .A1(w3[14]), .B0(n1152), .Y(n1153) );
  OAI21XL U1811 ( .A0(text_in_r[15]), .A1(w3[15]), .B0(n1154), .Y(n1155) );
  OAI21XL U1812 ( .A0(text_in_r[17]), .A1(w3[17]), .B0(n1156), .Y(n1157) );
  OAI2BB1X1 U1813 ( .A0N(n4), .A1N(sa13_next[1]), .B0(n1157), .Y(N65) );
  OAI21XL U1814 ( .A0(text_in_r[18]), .A1(w3[18]), .B0(n1158), .Y(n1159) );
  OAI21XL U1815 ( .A0(text_in_r[19]), .A1(w3[19]), .B0(n1160), .Y(n1161) );
  OAI21XL U1816 ( .A0(text_in_r[20]), .A1(w3[20]), .B0(n1162), .Y(n1163) );
  OAI21XL U1817 ( .A0(text_in_r[21]), .A1(w3[21]), .B0(n1164), .Y(n1165) );
  OAI21XL U1818 ( .A0(text_in_r[22]), .A1(w3[22]), .B0(n1166), .Y(n1167) );
  OAI21XL U1819 ( .A0(text_in_r[23]), .A1(w3[23]), .B0(n1168), .Y(n1169) );
  OAI21XL U1820 ( .A0(text_in_r[24]), .A1(w3[24]), .B0(n1170), .Y(n1171) );
  OAI2BB1X1 U1821 ( .A0N(n4), .A1N(sa03_next[0]), .B0(n1171), .Y(N80) );
  OAI21XL U1822 ( .A0(text_in_r[25]), .A1(w3[25]), .B0(n1172), .Y(n1173) );
  OAI21XL U1823 ( .A0(text_in_r[26]), .A1(w3[26]), .B0(n1174), .Y(n1175) );
  OAI21XL U1824 ( .A0(text_in_r[27]), .A1(w3[27]), .B0(n1176), .Y(n1177) );
  OAI21XL U1825 ( .A0(text_in_r[28]), .A1(w3[28]), .B0(n1178), .Y(n1179) );
  OAI21XL U1826 ( .A0(text_in_r[31]), .A1(w3[31]), .B0(n1180), .Y(n1181) );
  OAI21XL U1827 ( .A0(text_in_r[33]), .A1(w2[1]), .B0(n1182), .Y(n1183) );
  OAI21XL U1828 ( .A0(text_in_r[34]), .A1(w2[2]), .B0(n1184), .Y(n1185) );
  NAND2X1 U1829 ( .A(ld), .B(rst), .Y(n139) );
  NAND2X1 U1830 ( .A(n3), .B(n959), .Y(n1190) );
  NOR2X1 U1831 ( .A(dcnt_2_), .B(n1190), .Y(n1189) );
  INVX1 U1832 ( .A(rst), .Y(n1186) );
  AOI211X1 U1833 ( .A0(n1189), .A1(n2), .B0(ld), .C0(n1186), .Y(n1192) );
  OAI21XL U1834 ( .A0(n1189), .A1(n2), .B0(n966), .Y(n1187) );
  OAI21XL U1835 ( .A0(n3), .A1(n959), .B0(n1190), .Y(n1188) );
endmodule

//------------------------------------------------//
// LMDPL implementaiton for NOR
//-----------------------------------------------//

/*module nor_tablegen ( m_in0, m_in1, m_out, \t[7]_BAR , \t[3] , \t[2] , \t[1] , 
        \t[0] , \t[6]_BAR , \t[5]_BAR , \t[4]_BAR  );
  input m_in0, m_in1, m_out;
  output \t[7]_BAR , \t[3] , \t[2] , \t[1] , \t[0] , \t[6]_BAR , \t[5]_BAR ,
         \t[4]_BAR ;
  wire   \t[4]_BAR , \t[6]_BAR , \t[5]_BAR , \t[7]_BAR , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10;
  assign \t[0]  = \t[4]_BAR ;
  assign \t[2]  = \t[6]_BAR ;
  assign \t[1]  = \t[5]_BAR ;
  assign \t[3]  = \t[7]_BAR ;

  INVX1 U1 ( .A(m_out), .Y(n5) );
  NAND2X1 U2 ( .A(m_in1), .B(m_in0), .Y(n2) );
  NAND2X1 U3 ( .A(n5), .B(n2), .Y(n1) );
  OAI21XL U4 ( .A0(n5), .A1(n2), .B0(n1), .Y(\t[7]_BAR ) );
  INVX1 U5 ( .A(m_in1), .Y(n6) );
  NAND2X1 U6 ( .A(n6), .B(m_in0), .Y(n4) );
  NAND2X1 U7 ( .A(n5), .B(n4), .Y(n3) );
  OAI21XL U8 ( .A0(n5), .A1(n4), .B0(n3), .Y(\t[5]_BAR ) );
  NOR2X1 U9 ( .A(n6), .B(m_in0), .Y(n8) );
  NAND2X1 U10 ( .A(n8), .B(m_out), .Y(n7) );
  OAI21XL U11 ( .A0(n8), .A1(m_out), .B0(n7), .Y(\t[6]_BAR ) );
  NOR2X1 U12 ( .A(m_in1), .B(m_in0), .Y(n10) );
  NAND2X1 U13 ( .A(n10), .B(m_out), .Y(n9) );
  OAI21XL U14 ( .A0(n10), .A1(m_out), .B0(n9), .Y(\t[4]_BAR ) );
endmodule


module boolean_mask_dualrail_1 ( in, mask, in_m, in_m_bar );
  input in, mask;
  output in_m, in_m_bar;


  XNOR2X1 U1 ( .A(in), .B(mask), .Y(in_m_bar) );
  INVX1 U2 ( .A(in_m_bar), .Y(in_m) );
endmodule


module and3_lib ( in0, in1, in2, out );
  input in0, in1, in2;
  output out;


  AND3X1 and3_inst ( .A(in0), .B(in1), .C(in2), .Y(out) );
endmodule


module or4_lib ( in0, in1, in2, in3, out );
  input in0, in1, in2, in3;
  output out;


  OR4X1 or4_inst ( .A(in0), .B(in1), .C(in2), .D(in3), .Y(out) );
endmodule


module lmdpl_nl_gate ( t, a_m, a_m_bar, b_m, b_m_bar, q_m, q_m_bar );
  input [7:0] t;
  input a_m, a_m_bar, b_m, b_m_bar;
  output q_m, q_m_bar;

  wire   [7:0] and_out;

  and3_lib and3_inst_0 ( .in0(t[0]), .in1(a_m_bar), .in2(b_m_bar), .out(
        and_out[0]) );
  and3_lib and3_inst_1 ( .in0(t[1]), .in1(a_m), .in2(b_m_bar), .out(and_out[1]) );
  and3_lib and3_inst_2 ( .in0(t[2]), .in1(a_m_bar), .in2(b_m), .out(and_out[2]) );
  and3_lib and3_inst_3 ( .in0(t[3]), .in1(a_m), .in2(b_m), .out(and_out[3]) );
  and3_lib and3_inst_4 ( .in0(t[4]), .in1(a_m_bar), .in2(b_m_bar), .out(
        and_out[4]) );
  and3_lib and3_inst_5 ( .in0(t[5]), .in1(a_m), .in2(b_m_bar), .out(and_out[5]) );
  and3_lib and3_inst_6 ( .in0(t[6]), .in1(a_m_bar), .in2(b_m), .out(and_out[6]) );
  and3_lib and3_inst_7 ( .in0(t[7]), .in1(a_m), .in2(b_m), .out(and_out[7]) );
  or4_lib or4_inst_0 ( .in0(and_out[0]), .in1(and_out[1]), .in2(and_out[2]), 
        .in3(and_out[3]), .out(q_m_bar) );
  or4_lib or4_inst_1 ( .in0(and_out[4]), .in1(and_out[5]), .in2(and_out[6]), 
        .in3(and_out[7]), .out(q_m) );
endmodule


module boolean_mask_dualrail_0 ( in, mask, in_m, in_m_bar );
  input in, mask;
  output in_m, in_m_bar;


  XNOR2X1 U1 ( .A(in), .B(mask), .Y(in_m_bar) );
  INVX1 U2 ( .A(in_m_bar), .Y(in_m) );
endmodule


module nor_lmdpl ( clk, rst_n, precharge, in0, in1, m_in0, m_in1, m_out, out
 );
  input clk, rst_n, precharge, in0, in1, m_in0, m_in1, m_out;
  output out;
  wire   in0_m, in0_m_bar, in1_m, in1_m_bar, in0_m_pre_reg, in0_m_bar_pre_reg,
         in1_m_pre_reg, in1_m_bar_pre_reg, out_m, N16, n3, n4, n5, n6, n7, n8;
  wire   [7:0] t;
  wire   [7:0] t_reg;

  nor_tablegen nor_tablegen_inst ( .m_in0(m_in0), .m_in1(m_in1), .m_out(m_out), 
        .\t[7]_BAR (t[7]), .\t[3] (t[3]), .\t[2] (t[2]), .\t[1] (t[1]), 
        .\t[0] (t[0]), .\t[6]_BAR (t[6]), .\t[5]_BAR (t[5]), .\t[4]_BAR (t[4])
         );
  boolean_mask_dualrail_1 boolean_mask_dualrail_inst0 ( .in(in0), .mask(m_in0), 
        .in_m(in0_m), .in_m_bar(in0_m_bar) );
  boolean_mask_dualrail_0 boolean_mask_dualrail_inst1 ( .in(in1), .mask(m_in1), 
        .in_m(in1_m), .in_m_bar(in1_m_bar) );
  lmdpl_nl_gate lmdpl_nl_gate_inst ( .t(t_reg), .a_m(in0_m_pre_reg), .a_m_bar(
        in0_m_bar_pre_reg), .b_m(in1_m_pre_reg), .b_m_bar(in1_m_bar_pre_reg), 
        .q_m(out_m) );
  DFFHQX1 out_reg_reg ( .D(N16), .CK(clk), .Q(out) );
  DFFTRX1 t_reg_reg_3_ ( .D(t[3]), .RN(rst_n), .CK(clk), .Q(t_reg[3]) );
  DFFTRX1 t_reg_reg_2_ ( .D(t[2]), .RN(rst_n), .CK(clk), .Q(t_reg[2]) );
  DFFTRX1 t_reg_reg_1_ ( .D(t[1]), .RN(rst_n), .CK(clk), .Q(t_reg[1]) );
  DFFTRX1 t_reg_reg_0_ ( .D(t[0]), .RN(rst_n), .CK(clk), .Q(t_reg[0]) );
  DFFTRX1 t_reg_reg_7_ ( .D(n8), .RN(rst_n), .CK(clk), .Q(t_reg[7]) );
  DFFTRX1 t_reg_reg_6_ ( .D(n7), .RN(rst_n), .CK(clk), .Q(t_reg[6]) );
  DFFTRX1 t_reg_reg_5_ ( .D(n6), .RN(rst_n), .CK(clk), .Q(t_reg[5]) );
  DFFTRX1 t_reg_reg_4_ ( .D(n5), .RN(rst_n), .CK(clk), .Q(t_reg[4]) );
  DFFTRX1 in1_m_pre_reg_reg ( .D(n3), .RN(in1_m), .CK(clk), .Q(in1_m_pre_reg)
         );
  DFFTRX1 in1_m_bar_pre_reg_reg ( .D(n3), .RN(in1_m_bar), .CK(clk), .Q(
        in1_m_bar_pre_reg) );
  DFFTRX1 in0_m_pre_reg_reg ( .D(n3), .RN(in0_m), .CK(clk), .Q(in0_m_pre_reg)
         );
  DFFTRX1 in0_m_bar_pre_reg_reg ( .D(in0_m_bar), .RN(rst_n), .CK(clk), .Q(
        in0_m_bar_pre_reg) );
  AOI21XL U7 ( .A0(m_out), .A1(out_m), .B0(n4), .Y(N16) );
  INVX1 U8 ( .A(t[4]), .Y(n5) );
  INVX1 U9 ( .A(t[5]), .Y(n6) );
  INVX1 U10 ( .A(t[6]), .Y(n7) );
  INVX1 U11 ( .A(t[7]), .Y(n8) );
  NOR2BX1 U12 ( .AN(rst_n), .B(precharge), .Y(n3) );
  OAI21XL U13 ( .A0(m_out), .A1(out_m), .B0(rst_n), .Y(n4) );
endmodule
*/

//--------------------------------------------//
// combinational implemenent lmdpl
//--------------------------------------------//

module nor_tablegen ( m_in0, m_in1, m_out, t );
  output [7:0] t;
  input m_in0, m_in1, m_out;
  wire   N13, N15, N18, N21, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  assign t[7] = N13;
  assign t[6] = N15;
  assign t[5] = N18;
  assign t[4] = N21;

  INVX1 U1 ( .A(m_out), .Y(n8) );
  NAND2X1 U2 ( .A(m_in1), .B(m_in0), .Y(n2) );
  NAND2X1 U3 ( .A(n8), .B(n2), .Y(n1) );
  OAI21XL U4 ( .A0(n8), .A1(n2), .B0(n1), .Y(t[3]) );
  INVX1 U5 ( .A(t[3]), .Y(N13) );
  INVX1 U6 ( .A(m_in1), .Y(n5) );
  NOR2X1 U7 ( .A(n5), .B(m_in0), .Y(n4) );
  NAND2X1 U8 ( .A(n4), .B(m_out), .Y(n3) );
  OAI21XL U9 ( .A0(n4), .A1(m_out), .B0(n3), .Y(t[2]) );
  INVX1 U10 ( .A(t[2]), .Y(N15) );
  NAND2X1 U11 ( .A(n5), .B(m_in0), .Y(n7) );
  NAND2X1 U12 ( .A(n8), .B(n7), .Y(n6) );
  OAI21XL U13 ( .A0(n8), .A1(n7), .B0(n6), .Y(t[1]) );
  INVX1 U14 ( .A(t[1]), .Y(N18) );
  NOR2X1 U15 ( .A(m_in1), .B(m_in0), .Y(n10) );
  NAND2X1 U16 ( .A(n10), .B(m_out), .Y(n9) );
  OAI21XL U17 ( .A0(n10), .A1(m_out), .B0(n9), .Y(t[0]) );
  INVX1 U18 ( .A(t[0]), .Y(N21) );
endmodule


module boolean_mask_dualrail_1 ( in, mask, in_m, in_m_bar );
  input in, mask;
  output in_m, in_m_bar;


  XNOR2X1 U1 ( .A(in), .B(mask), .Y(in_m_bar) );
endmodule


module and3_lib ( in0, in1, in2, out );
  input in0, in1, in2;
  output out;


  AND3X1 and3_inst ( .A(in0), .B(in1), .C(in2), .Y(out) );
endmodule


module or4_lib ( in0, in1, in2, in3, out );
  input in0, in1, in2, in3;
  output out;


  OR4X1 or4_inst ( .A(in0), .B(in1), .C(in2), .D(in3), .Y(out) );
endmodule


module lmdpl_nl_gate ( t, a_m, a_m_bar, b_m, b_m_bar, q_m, q_m_bar );
  input [7:0] t;
  input a_m, a_m_bar, b_m, b_m_bar;
  output q_m, q_m_bar;

  wire   [7:0] and_out;

  and3_lib and3_inst_0 ( .in0(t[0]), .in1(a_m_bar), .in2(b_m_bar), .out(
        and_out[0]) );
  and3_lib and3_inst_1 ( .in0(t[1]), .in1(a_m), .in2(b_m_bar), .out(and_out[1]) );
  and3_lib and3_inst_2 ( .in0(t[2]), .in1(a_m_bar), .in2(b_m), .out(and_out[2]) );
  and3_lib and3_inst_3 ( .in0(t[3]), .in1(a_m), .in2(b_m), .out(and_out[3]) );
  and3_lib and3_inst_4 ( .in0(t[4]), .in1(a_m_bar), .in2(b_m_bar), .out(
        and_out[4]) );
  and3_lib and3_inst_5 ( .in0(t[5]), .in1(a_m), .in2(b_m_bar), .out(and_out[5]) );
  and3_lib and3_inst_6 ( .in0(t[6]), .in1(a_m_bar), .in2(b_m), .out(and_out[6]) );
  and3_lib and3_inst_7 ( .in0(t[7]), .in1(a_m), .in2(b_m), .out(and_out[7]) );
  or4_lib or4_inst_0 ( .in0(and_out[0]), .in1(and_out[1]), .in2(and_out[2]), 
        .in3(and_out[3]), .out(q_m_bar) );
  or4_lib or4_inst_1 ( .in0(and_out[4]), .in1(and_out[5]), .in2(and_out[6]), 
        .in3(and_out[7]), .out(q_m) );
endmodule


module boolean_mask_dualrail_0 ( in, mask, in_m, in_m_bar );
  input in, mask;
  output in_m, in_m_bar;


  XNOR2X1 U1 ( .A(in), .B(mask), .Y(in_m_bar) );
endmodule


module nor_lmdpl ( clk, rst_n, precharge, in0, in1, m_in0, m_in1, m_out, out
 );
  input clk, rst_n, precharge, in0, in1, m_in0, m_in1, m_out;
  output out;
  wire   in0_m_bar, in1_m_bar, in0_m_pre, in0_m_bar_pre, in1_m_pre,
         in1_m_bar_pre, out_m, out_m_bar, n4, n5, n6;
  wire   [7:0] t;

  nor_tablegen nor_tablegen_inst ( .m_in0(m_in0), .m_in1(m_in1), .m_out(m_out), 
        .t(t) );
  boolean_mask_dualrail_1 boolean_mask_dualrail_inst0 ( .in(in0), .mask(m_in0), 
        .in_m_bar(in0_m_bar) );
  boolean_mask_dualrail_0 boolean_mask_dualrail_inst1 ( .in(in1), .mask(m_in1), 
        .in_m_bar(in1_m_bar) );
  lmdpl_nl_gate lmdpl_nl_gate_inst ( .t(t), .a_m(in0_m_pre), .a_m_bar(
        in0_m_bar_pre), .b_m(in1_m_pre), .b_m_bar(in1_m_bar_pre), .q_m(out_m), 
        .q_m_bar(out_m_bar) );
  NOR2BX1 U9 ( .AN(in0_m_bar), .B(precharge), .Y(in0_m_bar_pre) );
  NOR2X1 U10 ( .A(precharge), .B(in0_m_bar), .Y(in0_m_pre) );
  NOR2BX1 U11 ( .AN(in1_m_bar), .B(precharge), .Y(in1_m_bar_pre) );
  NOR2X1 U12 ( .A(precharge), .B(in1_m_bar), .Y(in1_m_pre) );
  INVX1 U13 ( .A(out_m_bar), .Y(n6) );
  INVX1 U14 ( .A(out_m), .Y(n5) );
  INVX1 U15 ( .A(m_out), .Y(n4) );
  AOI33X1 U16 ( .A0(m_out), .A1(out_m), .A2(n6), .B0(out_m_bar), .B1(n5), .B2(
        n4), .Y(out) );
endmodule




