library verilog;
use verilog.vl_types.all;
entity PVDD2POC is
    port(
        VDDPST          : inout  vl_logic
    );
end PVDD2POC;
