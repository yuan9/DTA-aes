library verilog;
use verilog.vl_types.all;
entity PRO16CDG is
    port(
        I               : in     vl_logic;
        PAD             : out    vl_logic
    );
end PRO16CDG;
