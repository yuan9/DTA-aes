library verilog;
use verilog.vl_types.all;
entity udp_rslat_out is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end udp_rslat_out;
