library verilog;
use verilog.vl_types.all;
entity PDO24CDG is
    port(
        I               : in     vl_logic;
        PAD             : out    vl_logic
    );
end PDO24CDG;
