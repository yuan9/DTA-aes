library verilog;
use verilog.vl_types.all;
entity PVSS1DGZ is
    port(
        VSS             : inout  vl_logic
    );
end PVSS1DGZ;
