library verilog;
use verilog.vl_types.all;
entity \udp_rslatn_out_\ is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end \udp_rslatn_out_\;
