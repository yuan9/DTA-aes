library verilog;
use verilog.vl_types.all;
entity boolean_mask_dualrail_1 is
    port(
        \in\            : in     vl_logic;
        mask            : in     vl_logic;
        in_m            : out    vl_logic;
        in_m_bar        : out    vl_logic
    );
end boolean_mask_dualrail_1;
