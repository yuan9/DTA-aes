library verilog;
use verilog.vl_types.all;
entity PDO08CDG is
    port(
        I               : in     vl_logic;
        PAD             : out    vl_logic
    );
end PDO08CDG;
