library verilog;
use verilog.vl_types.all;
entity PVSS2ANA is
    port(
        AVSS            : inout  vl_logic
    );
end PVSS2ANA;
