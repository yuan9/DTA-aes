library verilog;
use verilog.vl_types.all;
entity PVDD2ANA is
    port(
        AVDD            : inout  vl_logic
    );
end PVDD2ANA;
