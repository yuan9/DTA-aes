
module aes_sbox_4 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358;

  OAI32X1 U1 ( .A0(n210), .A1(n145), .A2(n18), .B0(n27), .B1(n211), .Y(n209)
         );
  AOI221X1 U2 ( .A0(n278), .A1(n40), .B0(n185), .B1(n2), .C0(n279), .Y(n273)
         );
  OAI32X1 U3 ( .A0(n18), .A1(a[1]), .A2(n159), .B0(a[4]), .B1(n182), .Y(n318)
         );
  AOI31XL U4 ( .A0(n79), .A1(n44), .A2(n2), .B0(n280), .Y(n339) );
  AOI31X1 U5 ( .A0(n44), .A1(n129), .A2(n130), .B0(n131), .Y(n128) );
  AOI222XL U6 ( .A0(n185), .A1(n43), .B0(n186), .B1(n187), .C0(n6), .C1(n188), 
        .Y(n164) );
  AOI221X1 U7 ( .A0(n40), .A1(n136), .B0(n33), .B1(n47), .C0(n156), .Y(n141)
         );
  AOI222XL U8 ( .A0(n59), .A1(n43), .B0(n6), .B1(n221), .C0(n222), .C1(n187), 
        .Y(n218) );
  AOI221X1 U9 ( .A0(n225), .A1(n226), .B0(n296), .B1(n6), .C0(n297), .Y(n291)
         );
  AOI221X1 U10 ( .A0(n313), .A1(n5), .B0(n23), .B1(n2), .C0(n328), .Y(n320) );
  AOI221XL U11 ( .A0(n314), .A1(n43), .B0(n160), .B1(n24), .C0(n315), .Y(n307)
         );
  AOI221XL U12 ( .A0(n5), .A1(n96), .B0(n43), .B1(n239), .C0(n340), .Y(n336)
         );
  AOI221X1 U13 ( .A0(n40), .A1(n136), .B0(n33), .B1(n178), .C0(n338), .Y(n337)
         );
  AOI31X1 U14 ( .A0(a[2]), .A1(n58), .A2(a[1]), .B0(n40), .Y(n350) );
  OR2X2 U15 ( .A(a[2]), .B(a[7]), .Y(n1) );
  AOI221X1 U16 ( .A0(n5), .A1(n19), .B0(n33), .B1(n34), .C0(n35), .Y(n11) );
  OAI222X1 U17 ( .A0(n4), .A1(n37), .B0(n38), .B1(n20), .C0(a[4]), .C1(n39), 
        .Y(n35) );
  OAI222X1 U18 ( .A0(n20), .A1(n99), .B0(n27), .B1(n101), .C0(n184), .C1(n4), 
        .Y(n250) );
  OAI222X1 U19 ( .A0(n27), .A1(n34), .B0(n69), .B1(n205), .C0(n20), .C1(n79), 
        .Y(n260) );
  NAND2X2 U20 ( .A(n58), .B(n226), .Y(n34) );
  NOR2BXL U21 ( .AN(n101), .B(n25), .Y(n172) );
  AOI221XL U22 ( .A0(n43), .A1(n151), .B0(n25), .B1(n69), .C0(n275), .Y(n274)
         );
  NAND2XL U23 ( .A(n111), .B(n121), .Y(n303) );
  NAND2XL U24 ( .A(n111), .B(n300), .Y(n187) );
  NAND2XL U25 ( .A(n111), .B(n101), .Y(n21) );
  OAI2BB2XL U26 ( .B0(n20), .B1(n111), .A0N(n125), .A1N(n24), .Y(n220) );
  NAND2XL U27 ( .A(n198), .B(n24), .Y(n132) );
  AOI22XL U28 ( .A0(n33), .A1(a[3]), .B0(n24), .B1(n58), .Y(n277) );
  AOI22XL U29 ( .A0(n23), .A1(n24), .B0(n25), .B1(a[2]), .Y(n22) );
  AOI21XL U30 ( .A0(n44), .A1(n111), .B0(n4), .Y(n177) );
  NOR2X2 U31 ( .A(n44), .B(a[1]), .Y(n137) );
  CLKINVX3 U32 ( .A(n259), .Y(n44) );
  NOR2X2 U33 ( .A(n259), .B(n278), .Y(n47) );
  NOR2X2 U34 ( .A(a[4]), .B(a[3]), .Y(n278) );
  NOR2X2 U35 ( .A(n136), .B(n58), .Y(n259) );
  NOR2X2 U36 ( .A(n58), .B(a[3]), .Y(n159) );
  CLKINVX3 U37 ( .A(a[4]), .Y(n58) );
  NOR2X2 U38 ( .A(n136), .B(a[4]), .Y(n145) );
  CLKINVX3 U39 ( .A(a[3]), .Y(n136) );
  NOR2X4 U40 ( .A(n226), .B(n4), .Y(n40) );
  INVX4 U41 ( .A(a[2]), .Y(n69) );
  AOI21XL U42 ( .A0(n18), .A1(n162), .B0(n25), .Y(n161) );
  INVX4 U43 ( .A(n6), .Y(n18) );
  INVXL U44 ( .A(n20), .Y(n2) );
  MXI2XL U45 ( .A(n2), .B(n6), .S0(n28), .Y(n311) );
  NOR2XL U46 ( .A(n33), .B(n2), .Y(n302) );
  AOI22XL U47 ( .A0(n184), .A1(n5), .B0(n198), .B1(n43), .Y(n197) );
  AOI22XL U48 ( .A0(n40), .A1(n94), .B0(n43), .B1(n187), .Y(n244) );
  AOI21XL U49 ( .A0(n159), .A1(n43), .B0(n40), .Y(n262) );
  AOI22XL U50 ( .A0(n43), .A1(n100), .B0(n24), .B1(n125), .Y(n124) );
  AOI22XL U51 ( .A0(n43), .A1(n303), .B0(n24), .B1(n96), .Y(n358) );
  AOI222X4 U52 ( .A0(n125), .A1(n33), .B0(n145), .B1(n40), .C0(n43), .C1(n184), 
        .Y(n183) );
  AOI222X4 U53 ( .A0(n278), .A1(n24), .B0(n42), .B1(n33), .C0(n43), .C1(n136), 
        .Y(n351) );
  AOI2BB2XL U54 ( .B0(n43), .B1(n94), .A0N(n120), .A1N(n4), .Y(n119) );
  AOI22XL U55 ( .A0(n82), .A1(n43), .B0(n83), .B1(n24), .Y(n81) );
  AOI22XL U56 ( .A0(n98), .A1(n43), .B0(n6), .B1(n99), .Y(n97) );
  AOI22XL U57 ( .A0(n217), .A1(n43), .B0(n33), .B1(n47), .Y(n216) );
  AOI221X4 U58 ( .A0(n43), .A1(n44), .B0(n45), .B1(n24), .C0(n46), .Y(n9) );
  AOI221X4 U59 ( .A0(n43), .A1(n205), .B0(n32), .B1(n6), .C0(n206), .Y(n201)
         );
  AOI221X4 U60 ( .A0(n43), .A1(n208), .B0(n76), .B1(n24), .C0(n209), .Y(n207)
         );
  AOI221X4 U61 ( .A0(n70), .A1(n43), .B0(n24), .B1(n71), .C0(n72), .Y(n53) );
  AOI222X4 U62 ( .A0(n123), .A1(n43), .B0(a[2]), .B1(n203), .C0(n6), .C1(n71), 
        .Y(n202) );
  AOI221X4 U63 ( .A0(n59), .A1(n33), .B0(n43), .B1(n126), .C0(n127), .Y(n113)
         );
  AOI221X4 U64 ( .A0(n24), .A1(n82), .B0(n43), .B1(n295), .C0(n173), .Y(n346)
         );
  INVX4 U65 ( .A(n43), .Y(n20) );
  INVXL U66 ( .A(n36), .Y(n3) );
  INVX4 U67 ( .A(n3), .Y(n4) );
  INVXL U68 ( .A(n24), .Y(n36) );
  CLKINVX3 U69 ( .A(n1), .Y(n5) );
  CLKINVX3 U70 ( .A(n1), .Y(n6) );
  INVX12 U71 ( .A(n33), .Y(n27) );
  NOR2X4 U72 ( .A(n69), .B(a[7]), .Y(n33) );
  CLKINVX3 U73 ( .A(a[0]), .Y(n234) );
  NOR2X2 U74 ( .A(n252), .B(a[0]), .Y(n89) );
  AOI22XL U75 ( .A0(n70), .A1(n24), .B0(n96), .B1(n129), .Y(n241) );
  NOR2X4 U76 ( .A(n129), .B(n69), .Y(n24) );
  CLKINVX3 U77 ( .A(a[7]), .Y(n129) );
  NOR2X2 U78 ( .A(n252), .B(n234), .Y(n55) );
  CLKINVX3 U79 ( .A(a[5]), .Y(n252) );
  AOI22XL U80 ( .A0(n225), .A1(n226), .B0(n6), .B1(n227), .Y(n224) );
  INVX4 U81 ( .A(a[1]), .Y(n226) );
  OAI22XL U82 ( .A0(n201), .A1(n52), .B0(n202), .B1(n114), .Y(n193) );
  CLKINVX3 U83 ( .A(n14), .Y(n52) );
  NOR2X4 U84 ( .A(n129), .B(a[2]), .Y(n43) );
  MX2X1 U85 ( .A(n7), .B(n8), .S0(a[6]), .Y(d[7]) );
  OAI221XL U86 ( .A0(n9), .A1(n10), .B0(n11), .B1(n12), .C0(n13), .Y(n8) );
  AOI22X1 U87 ( .A0(n14), .A1(n15), .B0(n16), .B1(n17), .Y(n13) );
  OAI221XL U88 ( .A0(n18), .A1(n19), .B0(n20), .B1(n21), .C0(n22), .Y(n17) );
  OAI221XL U89 ( .A0(n26), .A1(n27), .B0(n28), .B1(n20), .C0(n29), .Y(n15) );
  AOI21X1 U90 ( .A0(n5), .A1(n30), .B0(n31), .Y(n29) );
  INVX1 U91 ( .A(n32), .Y(n26) );
  INVX1 U92 ( .A(n40), .Y(n39) );
  NOR2X1 U93 ( .A(n41), .B(n42), .Y(n38) );
  OAI221XL U94 ( .A0(n47), .A1(n18), .B0(n27), .B1(n48), .C0(n49), .Y(n46) );
  INVX1 U95 ( .A(n50), .Y(n49) );
  OAI221XL U96 ( .A0(n51), .A1(n52), .B0(n53), .B1(n10), .C0(n54), .Y(n7) );
  AOI22X1 U97 ( .A0(n55), .A1(n56), .B0(n16), .B1(n57), .Y(n54) );
  OAI221XL U98 ( .A0(n58), .A1(n18), .B0(n59), .B1(n27), .C0(n60), .Y(n57) );
  AOI2BB2X1 U99 ( .B0(n61), .B1(n24), .A0N(n62), .A1N(n20), .Y(n60) );
  OAI221XL U100 ( .A0(n63), .A1(n64), .B0(n65), .B1(n27), .C0(n66), .Y(n56) );
  INVX1 U101 ( .A(n67), .Y(n66) );
  AOI21X1 U102 ( .A0(n68), .A1(n69), .B0(n6), .Y(n63) );
  OAI211X1 U103 ( .A0(n73), .A1(n27), .B0(n74), .C0(n75), .Y(n72) );
  AOI211X1 U104 ( .A0(n5), .A1(n76), .B0(n77), .C0(n78), .Y(n51) );
  AOI21X1 U105 ( .A0(n79), .A1(n80), .B0(n27), .Y(n78) );
  INVX1 U106 ( .A(n81), .Y(n77) );
  MX2X1 U107 ( .A(n84), .B(n85), .S0(a[6]), .Y(d[6]) );
  OAI221XL U108 ( .A0(n86), .A1(n52), .B0(n87), .B1(n12), .C0(n88), .Y(n85) );
  AOI22X1 U109 ( .A0(n89), .A1(n90), .B0(n16), .B1(n91), .Y(n88) );
  OAI221XL U110 ( .A0(n73), .A1(n27), .B0(n92), .B1(n20), .C0(n93), .Y(n91) );
  AOI31X1 U111 ( .A0(n79), .A1(n94), .A2(n6), .B0(n67), .Y(n93) );
  NOR3X1 U112 ( .A(n4), .B(n95), .C(n96), .Y(n67) );
  OAI221XL U113 ( .A0(n27), .A1(n62), .B0(n4), .B1(n21), .C0(n97), .Y(n90) );
  NAND2X1 U114 ( .A(n100), .B(n101), .Y(n62) );
  AOI211X1 U115 ( .A0(n33), .A1(n102), .B0(n103), .C0(n104), .Y(n87) );
  AOI21X1 U116 ( .A0(n105), .A1(n106), .B0(n20), .Y(n104) );
  OAI22X1 U117 ( .A0(n45), .A1(n4), .B0(a[4]), .B1(n18), .Y(n103) );
  AOI211X1 U118 ( .A0(n5), .A1(n107), .B0(n108), .C0(n109), .Y(n86) );
  AOI21X1 U119 ( .A0(a[1]), .A1(n58), .B0(n27), .Y(n109) );
  OAI22X1 U120 ( .A0(n110), .A1(n4), .B0(n20), .B1(n21), .Y(n108) );
  OAI221XL U121 ( .A0(n112), .A1(n52), .B0(n113), .B1(n114), .C0(n115), .Y(n84) );
  AOI22X1 U122 ( .A0(n89), .A1(n116), .B0(n55), .B1(n117), .Y(n115) );
  OAI221XL U123 ( .A0(n18), .A1(n118), .B0(n27), .B1(n30), .C0(n119), .Y(n117)
         );
  NAND2X1 U124 ( .A(n121), .B(n122), .Y(n30) );
  OAI221XL U125 ( .A0(n18), .A1(n105), .B0(n123), .B1(n27), .C0(n124), .Y(n116) );
  OAI21XL U126 ( .A0(n18), .A1(n37), .B0(n128), .Y(n127) );
  INVX1 U127 ( .A(n132), .Y(n131) );
  AOI211X1 U128 ( .A0(n133), .A1(n69), .B0(n134), .C0(n135), .Y(n112) );
  OAI22X1 U129 ( .A0(n4), .A1(n136), .B0(n137), .B1(n27), .Y(n134) );
  INVX1 U130 ( .A(n70), .Y(n133) );
  MX2X1 U131 ( .A(n138), .B(n139), .S0(a[6]), .Y(d[5]) );
  OAI221XL U132 ( .A0(n140), .A1(n12), .B0(n141), .B1(n114), .C0(n142), .Y(
        n139) );
  AOI22X1 U133 ( .A0(n89), .A1(n143), .B0(n14), .B1(n144), .Y(n142) );
  OAI221XL U134 ( .A0(n145), .A1(n20), .B0(n4), .B1(n34), .C0(n146), .Y(n144)
         );
  AOI2BB1X1 U135 ( .A0N(n147), .A1N(n27), .B0(n148), .Y(n146) );
  AOI21X1 U136 ( .A0(n149), .A1(n150), .B0(n18), .Y(n148) );
  OAI221XL U137 ( .A0(n110), .A1(n18), .B0(n20), .B1(n151), .C0(n152), .Y(n143) );
  MXI2X1 U138 ( .A(n153), .B(n154), .S0(n155), .Y(n152) );
  NOR2X1 U139 ( .A(n145), .B(n69), .Y(n154) );
  NOR2X1 U140 ( .A(n4), .B(n136), .Y(n153) );
  OAI21XL U141 ( .A0(n157), .A1(n20), .B0(n158), .Y(n156) );
  AOI221X1 U142 ( .A0(n159), .A1(n24), .B0(n160), .B1(n33), .C0(n161), .Y(n140) );
  OAI21XL U143 ( .A0(n41), .A1(n163), .B0(n69), .Y(n162) );
  OAI221XL U144 ( .A0(n164), .A1(n114), .B0(n165), .B1(n52), .C0(n166), .Y(
        n138) );
  AOI22X1 U145 ( .A0(n89), .A1(n167), .B0(n55), .B1(n168), .Y(n166) );
  OAI211X1 U146 ( .A0(n20), .A1(n169), .B0(n170), .C0(n171), .Y(n168) );
  AOI22X1 U147 ( .A0(n137), .A1(n24), .B0(n172), .B1(n6), .Y(n171) );
  MXI2X1 U148 ( .A(n40), .B(n173), .S0(n96), .Y(n170) );
  OAI221XL U149 ( .A0(n159), .A1(n27), .B0(n145), .B1(n20), .C0(n174), .Y(n167) );
  AOI211X1 U150 ( .A0(n175), .A1(n5), .B0(n176), .C0(n177), .Y(n174) );
  INVX1 U151 ( .A(n178), .Y(n175) );
  AOI211X1 U152 ( .A0(n179), .A1(n24), .B0(n180), .C0(n181), .Y(n165) );
  NAND2X1 U153 ( .A(n74), .B(n182), .Y(n181) );
  INVX1 U154 ( .A(n183), .Y(n180) );
  OAI21XL U155 ( .A0(n69), .A1(n189), .B0(n27), .Y(n186) );
  MXI2X1 U156 ( .A(n190), .B(n191), .S0(a[6]), .Y(d[4]) );
  AOI211X1 U157 ( .A0(n89), .A1(n192), .B0(n193), .C0(n194), .Y(n191) );
  AOI31X1 U158 ( .A0(n195), .A1(n196), .A2(n197), .B0(n12), .Y(n194) );
  INVX1 U159 ( .A(n55), .Y(n12) );
  OAI2BB1X1 U160 ( .A0N(n199), .A1N(n200), .B0(n33), .Y(n195) );
  NAND2X1 U161 ( .A(n94), .B(n79), .Y(n203) );
  INVX1 U162 ( .A(n118), .Y(n123) );
  NAND2X1 U163 ( .A(n204), .B(n80), .Y(n118) );
  OAI22X1 U164 ( .A0(n28), .A1(n4), .B0(n188), .B1(n27), .Y(n206) );
  NOR2X1 U165 ( .A(n25), .B(n98), .Y(n32) );
  INVX1 U166 ( .A(n207), .Y(n192) );
  AOI211X1 U167 ( .A0(n55), .A1(n212), .B0(n213), .C0(n214), .Y(n190) );
  AOI31X1 U168 ( .A0(n215), .A1(n196), .A2(n216), .B0(n52), .Y(n214) );
  INVX1 U169 ( .A(n31), .Y(n196) );
  NOR2X1 U170 ( .A(n4), .B(n159), .Y(n31) );
  INVX1 U171 ( .A(n135), .Y(n215) );
  OAI22X1 U172 ( .A0(n218), .A1(n10), .B0(n219), .B1(n114), .Y(n213) );
  AOI211X1 U173 ( .A0(n208), .A1(n5), .B0(n220), .C0(n173), .Y(n219) );
  NOR2X1 U174 ( .A(n217), .B(n42), .Y(n208) );
  OAI21XL U175 ( .A0(n69), .A1(n223), .B0(n27), .Y(n222) );
  NAND2X1 U176 ( .A(n34), .B(n204), .Y(n221) );
  OAI221XL U177 ( .A0(n27), .A1(n64), .B0(n4), .B1(n83), .C0(n224), .Y(n212)
         );
  INVX1 U178 ( .A(n110), .Y(n64) );
  NOR2BX1 U179 ( .AN(n204), .B(n137), .Y(n110) );
  MX2X1 U180 ( .A(n228), .B(n229), .S0(a[6]), .Y(d[3]) );
  MX4X1 U181 ( .A(n230), .B(n231), .C(n232), .D(n233), .S0(n234), .S1(a[5]), 
        .Y(n229) );
  OAI211X1 U182 ( .A0(n27), .A1(n122), .B0(n158), .C0(n235), .Y(n233) );
  AOI2BB2X1 U183 ( .B0(n24), .B1(n187), .A0N(n227), .A1N(n20), .Y(n235) );
  OAI221XL U184 ( .A0(n18), .A1(n76), .B0(n59), .B1(n27), .C0(n236), .Y(n232)
         );
  OAI21XL U185 ( .A0(n237), .A1(n43), .B0(n238), .Y(n236) );
  INVX1 U186 ( .A(n239), .Y(n238) );
  AOI21X1 U187 ( .A0(n122), .A1(n106), .B0(n129), .Y(n237) );
  NAND2X1 U188 ( .A(n101), .B(n240), .Y(n76) );
  OAI221XL U189 ( .A0(n159), .A1(n27), .B0(n20), .B1(n34), .C0(n241), .Y(n231)
         );
  NOR2X1 U190 ( .A(n242), .B(n137), .Y(n70) );
  OAI211X1 U191 ( .A0(n4), .A1(n149), .B0(n243), .C0(n244), .Y(n230) );
  MXI2X1 U192 ( .A(n245), .B(n246), .S0(n130), .Y(n243) );
  XNOR2X1 U193 ( .A(n69), .B(a[1]), .Y(n130) );
  NOR2X1 U194 ( .A(a[7]), .B(n145), .Y(n246) );
  OAI21XL U195 ( .A0(n58), .A1(n27), .B0(n247), .Y(n245) );
  MXI2X1 U196 ( .A(n248), .B(n249), .S0(n234), .Y(n228) );
  MXI2X1 U197 ( .A(n250), .B(n251), .S0(n252), .Y(n249) );
  OAI221XL U198 ( .A0(n172), .A1(n18), .B0(n27), .B1(n83), .C0(n253), .Y(n251)
         );
  AOI2BB2X1 U199 ( .B0(n65), .B1(n24), .A0N(n169), .A1N(n20), .Y(n253) );
  NAND2X1 U200 ( .A(n199), .B(n204), .Y(n169) );
  NAND2X1 U201 ( .A(n200), .B(n106), .Y(n83) );
  INVX1 U202 ( .A(n211), .Y(n106) );
  AOI221X1 U203 ( .A0(n211), .A1(n5), .B0(n40), .B1(a[4]), .C0(n254), .Y(n248)
         );
  MXI2X1 U204 ( .A(n255), .B(n256), .S0(n252), .Y(n254) );
  NOR3X1 U205 ( .A(n257), .B(n258), .C(n50), .Y(n256) );
  OAI22X1 U206 ( .A0(n20), .A1(n68), .B0(n27), .B1(n37), .Y(n257) );
  AOI211X1 U207 ( .A0(n259), .A1(n24), .B0(n260), .C0(n261), .Y(n255) );
  INVX1 U208 ( .A(n262), .Y(n261) );
  NOR2X1 U209 ( .A(n94), .B(a[1]), .Y(n211) );
  MXI2X1 U210 ( .A(n263), .B(n264), .S0(a[6]), .Y(d[2]) );
  AOI211X1 U211 ( .A0(n55), .A1(n265), .B0(n266), .C0(n267), .Y(n264) );
  INVX1 U212 ( .A(n268), .Y(n267) );
  OAI31X1 U213 ( .A0(n176), .A1(n269), .A2(n270), .B0(n16), .Y(n268) );
  OAI21XL U214 ( .A0(n4), .A1(n271), .B0(n272), .Y(n270) );
  NOR2X1 U215 ( .A(n20), .B(n226), .Y(n176) );
  OAI22X1 U216 ( .A0(n273), .A1(n10), .B0(n274), .B1(n52), .Y(n266) );
  MXI2X1 U217 ( .A(n276), .B(n277), .S0(n155), .Y(n275) );
  XNOR2X1 U218 ( .A(n129), .B(a[1]), .Y(n155) );
  NAND2X1 U219 ( .A(a[2]), .B(n149), .Y(n276) );
  OAI221XL U220 ( .A0(a[1]), .A1(n247), .B0(n4), .B1(n189), .C0(n272), .Y(n279) );
  NAND2X1 U221 ( .A(n41), .B(n33), .Y(n272) );
  INVX1 U222 ( .A(n280), .Y(n247) );
  OAI221XL U223 ( .A0(n281), .A1(n27), .B0(n4), .B1(n111), .C0(n282), .Y(n265)
         );
  AOI211X1 U224 ( .A0(n5), .A1(n125), .B0(n50), .C0(n283), .Y(n282) );
  AOI21X1 U225 ( .A0(n200), .A1(n223), .B0(n20), .Y(n283) );
  NOR2X1 U226 ( .A(n199), .B(n4), .Y(n50) );
  NAND2X1 U227 ( .A(n284), .B(n122), .Y(n125) );
  AOI211X1 U228 ( .A0(n285), .A1(n55), .B0(n286), .C0(n287), .Y(n263) );
  AOI31X1 U229 ( .A0(n132), .A1(n288), .A2(n289), .B0(n52), .Y(n287) );
  AOI22X1 U230 ( .A0(n102), .A1(n69), .B0(n184), .B1(n33), .Y(n289) );
  NOR2X1 U231 ( .A(n290), .B(n163), .Y(n184) );
  NAND2X1 U232 ( .A(n200), .B(n284), .Y(n102) );
  INVX1 U233 ( .A(n225), .Y(n288) );
  OAI22X1 U234 ( .A0(n291), .A1(n114), .B0(n292), .B1(n10), .Y(n286) );
  INVX1 U235 ( .A(n89), .Y(n10) );
  AOI211X1 U236 ( .A0(n5), .A1(n79), .B0(n293), .C0(n294), .Y(n292) );
  AOI21X1 U237 ( .A0(n101), .A1(n150), .B0(n20), .Y(n294) );
  OAI2BB2X1 U238 ( .B0(n27), .B1(n295), .A0N(n34), .A1N(n24), .Y(n293) );
  OAI221XL U239 ( .A0(n298), .A1(n27), .B0(n20), .B1(n122), .C0(n132), .Y(n297) );
  NOR2X1 U240 ( .A(n159), .B(n217), .Y(n198) );
  NAND2X1 U241 ( .A(a[1]), .B(n47), .Y(n122) );
  NOR2X1 U242 ( .A(n299), .B(n242), .Y(n298) );
  INVX1 U243 ( .A(n99), .Y(n296) );
  NAND2X1 U244 ( .A(n200), .B(n300), .Y(n99) );
  MXI2X1 U245 ( .A(n301), .B(n147), .S0(n302), .Y(n285) );
  MXI2X1 U246 ( .A(n303), .B(n61), .S0(n69), .Y(n301) );
  INVX1 U247 ( .A(n187), .Y(n61) );
  MX2X1 U248 ( .A(n304), .B(n305), .S0(a[6]), .Y(d[1]) );
  OAI221XL U249 ( .A0(n306), .A1(n52), .B0(n307), .B1(n114), .C0(n308), .Y(
        n305) );
  AOI22X1 U250 ( .A0(n89), .A1(n309), .B0(n55), .B1(n310), .Y(n308) );
  OAI221XL U251 ( .A0(n27), .A1(n44), .B0(n4), .B1(n48), .C0(n311), .Y(n310)
         );
  AND2X1 U252 ( .A(n223), .B(n240), .Y(n28) );
  INVX1 U253 ( .A(n185), .Y(n48) );
  AOI21X1 U254 ( .A0(n226), .A1(n188), .B0(n242), .Y(n185) );
  OAI221XL U255 ( .A0(n149), .A1(n20), .B0(n4), .B1(n227), .C0(n312), .Y(n309)
         );
  AOI21X1 U256 ( .A0(n313), .A1(n33), .B0(n269), .Y(n312) );
  NAND2X1 U257 ( .A(n284), .B(n105), .Y(n227) );
  INVX1 U258 ( .A(n41), .Y(n105) );
  NOR2X1 U259 ( .A(n149), .B(n226), .Y(n41) );
  OAI22X1 U260 ( .A0(n92), .A1(n18), .B0(n316), .B1(n27), .Y(n315) );
  AOI21X1 U261 ( .A0(a[1]), .A1(n58), .B0(n98), .Y(n316) );
  INVX1 U262 ( .A(n295), .Y(n92) );
  NOR2X1 U263 ( .A(n45), .B(n163), .Y(n160) );
  INVX1 U264 ( .A(n151), .Y(n314) );
  NAND2X1 U265 ( .A(n100), .B(n199), .Y(n151) );
  AOI211X1 U266 ( .A0(n33), .A1(n120), .B0(n317), .C0(n318), .Y(n306) );
  INVX1 U267 ( .A(n258), .Y(n182) );
  OAI221XL U268 ( .A0(n20), .A1(n100), .B0(a[3]), .B1(n4), .C0(n262), .Y(n317)
         );
  INVX1 U269 ( .A(n210), .Y(n100) );
  NAND2X1 U270 ( .A(n34), .B(n200), .Y(n120) );
  INVX1 U271 ( .A(n290), .Y(n200) );
  NOR2X1 U272 ( .A(n226), .B(n58), .Y(n290) );
  OAI221XL U273 ( .A0(n319), .A1(n52), .B0(n320), .B1(n114), .C0(n321), .Y(
        n304) );
  AOI22X1 U274 ( .A0(n55), .A1(n322), .B0(n89), .B1(n323), .Y(n321) );
  OAI221XL U275 ( .A0(n47), .A1(n27), .B0(n65), .B1(n20), .C0(n324), .Y(n323)
         );
  AOI21X1 U276 ( .A0(n40), .A1(a[4]), .B0(n135), .Y(n324) );
  NOR2X1 U277 ( .A(n71), .B(n18), .Y(n135) );
  NAND2X1 U278 ( .A(n19), .B(n189), .Y(n71) );
  OAI21XL U279 ( .A0(n325), .A1(n18), .B0(n326), .Y(n322) );
  AOI31X1 U280 ( .A0(n111), .A1(n149), .A2(n327), .B0(n225), .Y(n326) );
  OAI21XL U281 ( .A0(n69), .A1(n284), .B0(n27), .Y(n327) );
  INVX1 U282 ( .A(n98), .Y(n284) );
  NOR2X1 U283 ( .A(n47), .B(a[1]), .Y(n98) );
  INVX1 U284 ( .A(n145), .Y(n149) );
  INVX1 U285 ( .A(n16), .Y(n114) );
  NOR2X1 U286 ( .A(a[0]), .B(a[5]), .Y(n16) );
  OAI32X1 U287 ( .A0(n4), .A1(n145), .A2(n210), .B0(n137), .B1(n27), .Y(n328)
         );
  AND2X1 U288 ( .A(n300), .B(n240), .Y(n23) );
  NAND2X1 U289 ( .A(n44), .B(n226), .Y(n300) );
  NOR2X1 U290 ( .A(n25), .B(n299), .Y(n313) );
  NOR2X1 U291 ( .A(n234), .B(a[5]), .Y(n14) );
  AOI221X1 U292 ( .A0(n325), .A1(n33), .B0(n24), .B1(n303), .C0(n329), .Y(n319) );
  OAI221XL U293 ( .A0(n18), .A1(n330), .B0(n20), .B1(n80), .C0(n75), .Y(n329)
         );
  INVX1 U294 ( .A(n269), .Y(n75) );
  NOR2X1 U295 ( .A(n111), .B(n18), .Y(n269) );
  INVX1 U296 ( .A(n299), .Y(n80) );
  MX4X1 U297 ( .A(n331), .B(n332), .C(n333), .D(n334), .S0(a[6]), .S1(n234), 
        .Y(d[0]) );
  NOR2X1 U298 ( .A(n258), .B(n335), .Y(n334) );
  MXI2X1 U299 ( .A(n336), .B(n337), .S0(n252), .Y(n335) );
  OAI21XL U300 ( .A0(n4), .A1(n121), .B0(n339), .Y(n338) );
  NOR2X1 U301 ( .A(n18), .B(n136), .Y(n280) );
  NAND2X1 U302 ( .A(n126), .B(n101), .Y(n178) );
  INVX1 U303 ( .A(n45), .Y(n126) );
  OAI32X1 U304 ( .A0(n27), .A1(n278), .A2(n95), .B0(n341), .B1(n4), .Y(n340)
         );
  NOR2X1 U305 ( .A(n299), .B(n210), .Y(n341) );
  NOR2X1 U306 ( .A(n136), .B(a[1]), .Y(n299) );
  NAND2X1 U307 ( .A(n204), .B(n330), .Y(n239) );
  INVX1 U308 ( .A(n179), .Y(n330) );
  NOR2X1 U309 ( .A(n188), .B(a[1]), .Y(n179) );
  NAND2X1 U310 ( .A(n278), .B(a[1]), .Y(n204) );
  NOR2X1 U311 ( .A(n18), .B(n226), .Y(n258) );
  AOI211X1 U312 ( .A0(n5), .A1(n68), .B0(n342), .C0(n343), .Y(n333) );
  AOI21X1 U313 ( .A0(n240), .A1(n37), .B0(n344), .Y(n343) );
  INVX1 U314 ( .A(n173), .Y(n344) );
  INVX1 U315 ( .A(n163), .Y(n37) );
  NOR2X1 U316 ( .A(a[1]), .B(a[3]), .Y(n163) );
  MXI2X1 U317 ( .A(n345), .B(n346), .S0(n252), .Y(n342) );
  NOR2X1 U318 ( .A(n27), .B(n210), .Y(n173) );
  NOR2X1 U319 ( .A(n226), .B(n259), .Y(n210) );
  NAND2X1 U320 ( .A(n19), .B(n199), .Y(n295) );
  NAND2X1 U321 ( .A(n199), .B(n205), .Y(n82) );
  NAND2X1 U322 ( .A(n94), .B(n226), .Y(n199) );
  INVX1 U323 ( .A(n278), .Y(n94) );
  NOR2X1 U324 ( .A(n225), .B(n40), .Y(n345) );
  NOR2X1 U325 ( .A(n20), .B(n159), .Y(n225) );
  NAND2X1 U326 ( .A(n240), .B(n189), .Y(n68) );
  INVX1 U327 ( .A(n157), .Y(n240) );
  NOR2X1 U328 ( .A(n44), .B(n226), .Y(n157) );
  MXI2X1 U329 ( .A(n347), .B(n348), .S0(n252), .Y(n332) );
  OAI211X1 U330 ( .A0(n349), .A1(n74), .B0(n350), .C0(n351), .Y(n348) );
  NAND2X1 U331 ( .A(n278), .B(n6), .Y(n74) );
  INVX1 U332 ( .A(n352), .Y(n349) );
  OAI221XL U333 ( .A0(n20), .A1(n34), .B0(n325), .B1(n4), .C0(n353), .Y(n347)
         );
  AOI31X1 U334 ( .A0(n6), .A1(n352), .A2(n259), .B0(n354), .Y(n353) );
  AOI21X1 U335 ( .A0(n19), .A1(n223), .B0(n27), .Y(n354) );
  NAND2X1 U336 ( .A(n145), .B(n226), .Y(n223) );
  INVX1 U337 ( .A(n281), .Y(n19) );
  NOR2X1 U338 ( .A(n226), .B(n136), .Y(n281) );
  XNOR2X1 U339 ( .A(a[5]), .B(n226), .Y(n352) );
  AND2X1 U340 ( .A(n101), .B(n79), .Y(n325) );
  INVX1 U341 ( .A(n59), .Y(n79) );
  MXI2X1 U342 ( .A(n355), .B(n356), .S0(n252), .Y(n331) );
  OAI221XL U343 ( .A0(n18), .A1(n121), .B0(n271), .B1(n20), .C0(n357), .Y(n356) );
  AOI22X1 U344 ( .A0(n33), .A1(n147), .B0(n24), .B1(n107), .Y(n357) );
  INVX1 U345 ( .A(n172), .Y(n107) );
  NOR2X1 U346 ( .A(n188), .B(n226), .Y(n25) );
  INVX1 U347 ( .A(n159), .Y(n188) );
  NAND2X1 U348 ( .A(a[4]), .B(n226), .Y(n101) );
  NAND2X1 U349 ( .A(n44), .B(n150), .Y(n147) );
  INVX1 U350 ( .A(n217), .Y(n150) );
  NOR2X1 U351 ( .A(n226), .B(n278), .Y(n217) );
  NOR2X1 U352 ( .A(n96), .B(n59), .Y(n271) );
  NOR2X1 U353 ( .A(n226), .B(n145), .Y(n59) );
  OAI211X1 U354 ( .A0(n65), .A1(n27), .B0(n158), .C0(n358), .Y(n355) );
  INVX1 U355 ( .A(n47), .Y(n96) );
  INVX1 U356 ( .A(n42), .Y(n121) );
  NOR2X1 U357 ( .A(n145), .B(a[1]), .Y(n42) );
  INVX1 U358 ( .A(n95), .Y(n111) );
  NOR2X1 U359 ( .A(n226), .B(n159), .Y(n95) );
  NAND2BX1 U360 ( .AN(n73), .B(n6), .Y(n158) );
  NOR2X1 U361 ( .A(n259), .B(n45), .Y(n73) );
  NOR2X1 U362 ( .A(n226), .B(n47), .Y(n45) );
  AND2X1 U363 ( .A(n189), .B(n205), .Y(n65) );
  INVX1 U364 ( .A(n242), .Y(n205) );
  NOR2X1 U365 ( .A(n226), .B(a[3]), .Y(n242) );
  NAND2X1 U366 ( .A(n47), .B(n226), .Y(n189) );
endmodule


module aes_sbox_3 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358;

  AOI31XL U1 ( .A0(n79), .A1(n44), .A2(n2), .B0(n280), .Y(n339) );
  AOI31X1 U2 ( .A0(n44), .A1(n129), .A2(n130), .B0(n131), .Y(n128) );
  AOI221X1 U3 ( .A0(n40), .A1(n136), .B0(n33), .B1(n47), .C0(n156), .Y(n141)
         );
  OAI32X1 U4 ( .A0(n210), .A1(n145), .A2(n18), .B0(n27), .B1(n211), .Y(n209)
         );
  AOI222XL U5 ( .A0(n59), .A1(n43), .B0(n6), .B1(n221), .C0(n222), .C1(n187), 
        .Y(n218) );
  AOI221X1 U6 ( .A0(n278), .A1(n40), .B0(n185), .B1(n2), .C0(n279), .Y(n273)
         );
  AOI221X1 U7 ( .A0(n225), .A1(n226), .B0(n296), .B1(n6), .C0(n297), .Y(n291)
         );
  OAI32X1 U8 ( .A0(n18), .A1(a[1]), .A2(n159), .B0(a[4]), .B1(n182), .Y(n318)
         );
  AOI221XL U9 ( .A0(n314), .A1(n43), .B0(n160), .B1(n24), .C0(n315), .Y(n307)
         );
  AOI221X1 U10 ( .A0(n313), .A1(n5), .B0(n23), .B1(n2), .C0(n328), .Y(n320) );
  AOI31X1 U11 ( .A0(a[2]), .A1(n58), .A2(a[1]), .B0(n40), .Y(n350) );
  AOI222XL U12 ( .A0(n278), .A1(n24), .B0(n42), .B1(n33), .C0(n43), .C1(n136), 
        .Y(n351) );
  AOI221XL U13 ( .A0(n5), .A1(n96), .B0(n43), .B1(n239), .C0(n340), .Y(n336)
         );
  AOI221X1 U14 ( .A0(n40), .A1(n136), .B0(n33), .B1(n178), .C0(n338), .Y(n337)
         );
  OR2X2 U15 ( .A(a[2]), .B(a[7]), .Y(n1) );
  AOI221X1 U16 ( .A0(n5), .A1(n19), .B0(n33), .B1(n34), .C0(n35), .Y(n11) );
  OAI222X1 U17 ( .A0(n4), .A1(n37), .B0(n38), .B1(n20), .C0(a[4]), .C1(n39), 
        .Y(n35) );
  OAI222X1 U18 ( .A0(n20), .A1(n99), .B0(n27), .B1(n101), .C0(n184), .C1(n4), 
        .Y(n250) );
  OAI222X1 U19 ( .A0(n27), .A1(n34), .B0(n69), .B1(n205), .C0(n20), .C1(n79), 
        .Y(n260) );
  NAND2X2 U20 ( .A(n58), .B(n226), .Y(n34) );
  NOR2BXL U21 ( .AN(n101), .B(n25), .Y(n172) );
  AOI221XL U22 ( .A0(n43), .A1(n151), .B0(n25), .B1(n69), .C0(n275), .Y(n274)
         );
  NAND2XL U23 ( .A(n111), .B(n121), .Y(n303) );
  NAND2XL U24 ( .A(n111), .B(n300), .Y(n187) );
  NAND2XL U25 ( .A(n111), .B(n101), .Y(n21) );
  OAI2BB2XL U26 ( .B0(n20), .B1(n111), .A0N(n125), .A1N(n24), .Y(n220) );
  NAND2XL U27 ( .A(n198), .B(n24), .Y(n132) );
  AOI22XL U28 ( .A0(n33), .A1(a[3]), .B0(n24), .B1(n58), .Y(n277) );
  AOI22XL U29 ( .A0(n23), .A1(n24), .B0(n25), .B1(a[2]), .Y(n22) );
  AOI21XL U30 ( .A0(n44), .A1(n111), .B0(n4), .Y(n177) );
  NOR2X2 U31 ( .A(n44), .B(a[1]), .Y(n137) );
  CLKINVX3 U32 ( .A(n259), .Y(n44) );
  NOR2X2 U33 ( .A(n259), .B(n278), .Y(n47) );
  NOR2X2 U34 ( .A(a[4]), .B(a[3]), .Y(n278) );
  NOR2X2 U35 ( .A(n136), .B(n58), .Y(n259) );
  NOR2X2 U36 ( .A(n58), .B(a[3]), .Y(n159) );
  CLKINVX3 U37 ( .A(a[4]), .Y(n58) );
  NOR2X2 U38 ( .A(n136), .B(a[4]), .Y(n145) );
  CLKINVX3 U39 ( .A(a[3]), .Y(n136) );
  NOR2X4 U40 ( .A(n226), .B(n4), .Y(n40) );
  INVX4 U41 ( .A(a[2]), .Y(n69) );
  AOI21XL U42 ( .A0(n18), .A1(n162), .B0(n25), .Y(n161) );
  INVX4 U43 ( .A(n6), .Y(n18) );
  INVXL U44 ( .A(n20), .Y(n2) );
  MXI2XL U45 ( .A(n2), .B(n6), .S0(n28), .Y(n311) );
  NOR2XL U46 ( .A(n33), .B(n2), .Y(n302) );
  AOI22XL U47 ( .A0(n184), .A1(n5), .B0(n198), .B1(n43), .Y(n197) );
  AOI22XL U48 ( .A0(n40), .A1(n94), .B0(n43), .B1(n187), .Y(n244) );
  AOI21XL U49 ( .A0(n159), .A1(n43), .B0(n40), .Y(n262) );
  AOI22XL U50 ( .A0(n43), .A1(n100), .B0(n24), .B1(n125), .Y(n124) );
  AOI22XL U51 ( .A0(n43), .A1(n303), .B0(n24), .B1(n96), .Y(n358) );
  AOI222X4 U52 ( .A0(n125), .A1(n33), .B0(n145), .B1(n40), .C0(n43), .C1(n184), 
        .Y(n183) );
  AOI2BB2XL U53 ( .B0(n43), .B1(n94), .A0N(n120), .A1N(n4), .Y(n119) );
  AOI22XL U54 ( .A0(n82), .A1(n43), .B0(n83), .B1(n24), .Y(n81) );
  AOI22XL U55 ( .A0(n98), .A1(n43), .B0(n6), .B1(n99), .Y(n97) );
  AOI22XL U56 ( .A0(n217), .A1(n43), .B0(n33), .B1(n47), .Y(n216) );
  AOI221X4 U57 ( .A0(n43), .A1(n44), .B0(n45), .B1(n24), .C0(n46), .Y(n9) );
  AOI221X4 U58 ( .A0(n43), .A1(n205), .B0(n32), .B1(n6), .C0(n206), .Y(n201)
         );
  AOI221X4 U59 ( .A0(n43), .A1(n208), .B0(n76), .B1(n24), .C0(n209), .Y(n207)
         );
  AOI221X4 U60 ( .A0(n70), .A1(n43), .B0(n24), .B1(n71), .C0(n72), .Y(n53) );
  AOI222X4 U61 ( .A0(n185), .A1(n43), .B0(n186), .B1(n187), .C0(n6), .C1(n188), 
        .Y(n164) );
  AOI222X4 U62 ( .A0(n123), .A1(n43), .B0(a[2]), .B1(n203), .C0(n6), .C1(n71), 
        .Y(n202) );
  AOI221X4 U63 ( .A0(n59), .A1(n33), .B0(n43), .B1(n126), .C0(n127), .Y(n113)
         );
  AOI221X4 U64 ( .A0(n24), .A1(n82), .B0(n43), .B1(n295), .C0(n173), .Y(n346)
         );
  INVX4 U65 ( .A(n43), .Y(n20) );
  INVXL U66 ( .A(n36), .Y(n3) );
  INVX4 U67 ( .A(n3), .Y(n4) );
  INVXL U68 ( .A(n24), .Y(n36) );
  CLKINVX3 U69 ( .A(n1), .Y(n5) );
  CLKINVX3 U70 ( .A(n1), .Y(n6) );
  INVX12 U71 ( .A(n33), .Y(n27) );
  NOR2X4 U72 ( .A(n69), .B(a[7]), .Y(n33) );
  CLKINVX3 U73 ( .A(a[0]), .Y(n234) );
  NOR2X2 U74 ( .A(n252), .B(a[0]), .Y(n89) );
  AOI22XL U75 ( .A0(n70), .A1(n24), .B0(n96), .B1(n129), .Y(n241) );
  NOR2X4 U76 ( .A(n129), .B(n69), .Y(n24) );
  CLKINVX3 U77 ( .A(a[7]), .Y(n129) );
  NOR2X2 U78 ( .A(n252), .B(n234), .Y(n55) );
  CLKINVX3 U79 ( .A(a[5]), .Y(n252) );
  AOI22XL U80 ( .A0(n225), .A1(n226), .B0(n6), .B1(n227), .Y(n224) );
  INVX4 U81 ( .A(a[1]), .Y(n226) );
  OAI22XL U82 ( .A0(n201), .A1(n52), .B0(n202), .B1(n114), .Y(n193) );
  CLKINVX3 U83 ( .A(n14), .Y(n52) );
  NOR2X4 U84 ( .A(n129), .B(a[2]), .Y(n43) );
  MX2X1 U85 ( .A(n7), .B(n8), .S0(a[6]), .Y(d[7]) );
  OAI221XL U86 ( .A0(n9), .A1(n10), .B0(n11), .B1(n12), .C0(n13), .Y(n8) );
  AOI22X1 U87 ( .A0(n14), .A1(n15), .B0(n16), .B1(n17), .Y(n13) );
  OAI221XL U88 ( .A0(n18), .A1(n19), .B0(n20), .B1(n21), .C0(n22), .Y(n17) );
  OAI221XL U89 ( .A0(n26), .A1(n27), .B0(n28), .B1(n20), .C0(n29), .Y(n15) );
  AOI21X1 U90 ( .A0(n5), .A1(n30), .B0(n31), .Y(n29) );
  INVX1 U91 ( .A(n32), .Y(n26) );
  INVX1 U92 ( .A(n40), .Y(n39) );
  NOR2X1 U93 ( .A(n41), .B(n42), .Y(n38) );
  OAI221XL U94 ( .A0(n47), .A1(n18), .B0(n27), .B1(n48), .C0(n49), .Y(n46) );
  INVX1 U95 ( .A(n50), .Y(n49) );
  OAI221XL U96 ( .A0(n51), .A1(n52), .B0(n53), .B1(n10), .C0(n54), .Y(n7) );
  AOI22X1 U97 ( .A0(n55), .A1(n56), .B0(n16), .B1(n57), .Y(n54) );
  OAI221XL U98 ( .A0(n58), .A1(n18), .B0(n59), .B1(n27), .C0(n60), .Y(n57) );
  AOI2BB2X1 U99 ( .B0(n61), .B1(n24), .A0N(n62), .A1N(n20), .Y(n60) );
  OAI221XL U100 ( .A0(n63), .A1(n64), .B0(n65), .B1(n27), .C0(n66), .Y(n56) );
  INVX1 U101 ( .A(n67), .Y(n66) );
  AOI21X1 U102 ( .A0(n68), .A1(n69), .B0(n6), .Y(n63) );
  OAI211X1 U103 ( .A0(n73), .A1(n27), .B0(n74), .C0(n75), .Y(n72) );
  AOI211X1 U104 ( .A0(n5), .A1(n76), .B0(n77), .C0(n78), .Y(n51) );
  AOI21X1 U105 ( .A0(n79), .A1(n80), .B0(n27), .Y(n78) );
  INVX1 U106 ( .A(n81), .Y(n77) );
  MX2X1 U107 ( .A(n84), .B(n85), .S0(a[6]), .Y(d[6]) );
  OAI221XL U108 ( .A0(n86), .A1(n52), .B0(n87), .B1(n12), .C0(n88), .Y(n85) );
  AOI22X1 U109 ( .A0(n89), .A1(n90), .B0(n16), .B1(n91), .Y(n88) );
  OAI221XL U110 ( .A0(n73), .A1(n27), .B0(n92), .B1(n20), .C0(n93), .Y(n91) );
  AOI31X1 U111 ( .A0(n79), .A1(n94), .A2(n6), .B0(n67), .Y(n93) );
  NOR3X1 U112 ( .A(n4), .B(n95), .C(n96), .Y(n67) );
  OAI221XL U113 ( .A0(n27), .A1(n62), .B0(n4), .B1(n21), .C0(n97), .Y(n90) );
  NAND2X1 U114 ( .A(n100), .B(n101), .Y(n62) );
  AOI211X1 U115 ( .A0(n33), .A1(n102), .B0(n103), .C0(n104), .Y(n87) );
  AOI21X1 U116 ( .A0(n105), .A1(n106), .B0(n20), .Y(n104) );
  OAI22X1 U117 ( .A0(n45), .A1(n4), .B0(a[4]), .B1(n18), .Y(n103) );
  AOI211X1 U118 ( .A0(n5), .A1(n107), .B0(n108), .C0(n109), .Y(n86) );
  AOI21X1 U119 ( .A0(a[1]), .A1(n58), .B0(n27), .Y(n109) );
  OAI22X1 U120 ( .A0(n110), .A1(n4), .B0(n20), .B1(n21), .Y(n108) );
  OAI221XL U121 ( .A0(n112), .A1(n52), .B0(n113), .B1(n114), .C0(n115), .Y(n84) );
  AOI22X1 U122 ( .A0(n89), .A1(n116), .B0(n55), .B1(n117), .Y(n115) );
  OAI221XL U123 ( .A0(n18), .A1(n118), .B0(n27), .B1(n30), .C0(n119), .Y(n117)
         );
  NAND2X1 U124 ( .A(n121), .B(n122), .Y(n30) );
  OAI221XL U125 ( .A0(n18), .A1(n105), .B0(n123), .B1(n27), .C0(n124), .Y(n116) );
  OAI21XL U126 ( .A0(n18), .A1(n37), .B0(n128), .Y(n127) );
  INVX1 U127 ( .A(n132), .Y(n131) );
  AOI211X1 U128 ( .A0(n133), .A1(n69), .B0(n134), .C0(n135), .Y(n112) );
  OAI22X1 U129 ( .A0(n4), .A1(n136), .B0(n137), .B1(n27), .Y(n134) );
  INVX1 U130 ( .A(n70), .Y(n133) );
  MX2X1 U131 ( .A(n138), .B(n139), .S0(a[6]), .Y(d[5]) );
  OAI221XL U132 ( .A0(n140), .A1(n12), .B0(n141), .B1(n114), .C0(n142), .Y(
        n139) );
  AOI22X1 U133 ( .A0(n89), .A1(n143), .B0(n14), .B1(n144), .Y(n142) );
  OAI221XL U134 ( .A0(n145), .A1(n20), .B0(n4), .B1(n34), .C0(n146), .Y(n144)
         );
  AOI2BB1X1 U135 ( .A0N(n147), .A1N(n27), .B0(n148), .Y(n146) );
  AOI21X1 U136 ( .A0(n149), .A1(n150), .B0(n18), .Y(n148) );
  OAI221XL U137 ( .A0(n110), .A1(n18), .B0(n20), .B1(n151), .C0(n152), .Y(n143) );
  MXI2X1 U138 ( .A(n153), .B(n154), .S0(n155), .Y(n152) );
  NOR2X1 U139 ( .A(n145), .B(n69), .Y(n154) );
  NOR2X1 U140 ( .A(n4), .B(n136), .Y(n153) );
  OAI21XL U141 ( .A0(n157), .A1(n20), .B0(n158), .Y(n156) );
  AOI221X1 U142 ( .A0(n159), .A1(n24), .B0(n160), .B1(n33), .C0(n161), .Y(n140) );
  OAI21XL U143 ( .A0(n41), .A1(n163), .B0(n69), .Y(n162) );
  OAI221XL U144 ( .A0(n164), .A1(n114), .B0(n165), .B1(n52), .C0(n166), .Y(
        n138) );
  AOI22X1 U145 ( .A0(n89), .A1(n167), .B0(n55), .B1(n168), .Y(n166) );
  OAI211X1 U146 ( .A0(n20), .A1(n169), .B0(n170), .C0(n171), .Y(n168) );
  AOI22X1 U147 ( .A0(n137), .A1(n24), .B0(n172), .B1(n6), .Y(n171) );
  MXI2X1 U148 ( .A(n40), .B(n173), .S0(n96), .Y(n170) );
  OAI221XL U149 ( .A0(n159), .A1(n27), .B0(n145), .B1(n20), .C0(n174), .Y(n167) );
  AOI211X1 U150 ( .A0(n175), .A1(n5), .B0(n176), .C0(n177), .Y(n174) );
  INVX1 U151 ( .A(n178), .Y(n175) );
  AOI211X1 U152 ( .A0(n179), .A1(n24), .B0(n180), .C0(n181), .Y(n165) );
  NAND2X1 U153 ( .A(n74), .B(n182), .Y(n181) );
  INVX1 U154 ( .A(n183), .Y(n180) );
  OAI21XL U155 ( .A0(n69), .A1(n189), .B0(n27), .Y(n186) );
  MXI2X1 U156 ( .A(n190), .B(n191), .S0(a[6]), .Y(d[4]) );
  AOI211X1 U157 ( .A0(n89), .A1(n192), .B0(n193), .C0(n194), .Y(n191) );
  AOI31X1 U158 ( .A0(n195), .A1(n196), .A2(n197), .B0(n12), .Y(n194) );
  INVX1 U159 ( .A(n55), .Y(n12) );
  OAI2BB1X1 U160 ( .A0N(n199), .A1N(n200), .B0(n33), .Y(n195) );
  NAND2X1 U161 ( .A(n94), .B(n79), .Y(n203) );
  INVX1 U162 ( .A(n118), .Y(n123) );
  NAND2X1 U163 ( .A(n204), .B(n80), .Y(n118) );
  OAI22X1 U164 ( .A0(n28), .A1(n4), .B0(n188), .B1(n27), .Y(n206) );
  NOR2X1 U165 ( .A(n25), .B(n98), .Y(n32) );
  INVX1 U166 ( .A(n207), .Y(n192) );
  AOI211X1 U167 ( .A0(n55), .A1(n212), .B0(n213), .C0(n214), .Y(n190) );
  AOI31X1 U168 ( .A0(n215), .A1(n196), .A2(n216), .B0(n52), .Y(n214) );
  INVX1 U169 ( .A(n31), .Y(n196) );
  NOR2X1 U170 ( .A(n4), .B(n159), .Y(n31) );
  INVX1 U171 ( .A(n135), .Y(n215) );
  OAI22X1 U172 ( .A0(n218), .A1(n10), .B0(n219), .B1(n114), .Y(n213) );
  AOI211X1 U173 ( .A0(n208), .A1(n5), .B0(n220), .C0(n173), .Y(n219) );
  NOR2X1 U174 ( .A(n217), .B(n42), .Y(n208) );
  OAI21XL U175 ( .A0(n69), .A1(n223), .B0(n27), .Y(n222) );
  NAND2X1 U176 ( .A(n34), .B(n204), .Y(n221) );
  OAI221XL U177 ( .A0(n27), .A1(n64), .B0(n4), .B1(n83), .C0(n224), .Y(n212)
         );
  INVX1 U178 ( .A(n110), .Y(n64) );
  NOR2BX1 U179 ( .AN(n204), .B(n137), .Y(n110) );
  MX2X1 U180 ( .A(n228), .B(n229), .S0(a[6]), .Y(d[3]) );
  MX4X1 U181 ( .A(n230), .B(n231), .C(n232), .D(n233), .S0(n234), .S1(a[5]), 
        .Y(n229) );
  OAI211X1 U182 ( .A0(n27), .A1(n122), .B0(n158), .C0(n235), .Y(n233) );
  AOI2BB2X1 U183 ( .B0(n24), .B1(n187), .A0N(n227), .A1N(n20), .Y(n235) );
  OAI221XL U184 ( .A0(n18), .A1(n76), .B0(n59), .B1(n27), .C0(n236), .Y(n232)
         );
  OAI21XL U185 ( .A0(n237), .A1(n43), .B0(n238), .Y(n236) );
  INVX1 U186 ( .A(n239), .Y(n238) );
  AOI21X1 U187 ( .A0(n122), .A1(n106), .B0(n129), .Y(n237) );
  NAND2X1 U188 ( .A(n101), .B(n240), .Y(n76) );
  OAI221XL U189 ( .A0(n159), .A1(n27), .B0(n20), .B1(n34), .C0(n241), .Y(n231)
         );
  NOR2X1 U190 ( .A(n242), .B(n137), .Y(n70) );
  OAI211X1 U191 ( .A0(n4), .A1(n149), .B0(n243), .C0(n244), .Y(n230) );
  MXI2X1 U192 ( .A(n245), .B(n246), .S0(n130), .Y(n243) );
  XNOR2X1 U193 ( .A(n69), .B(a[1]), .Y(n130) );
  NOR2X1 U194 ( .A(a[7]), .B(n145), .Y(n246) );
  OAI21XL U195 ( .A0(n58), .A1(n27), .B0(n247), .Y(n245) );
  MXI2X1 U196 ( .A(n248), .B(n249), .S0(n234), .Y(n228) );
  MXI2X1 U197 ( .A(n250), .B(n251), .S0(n252), .Y(n249) );
  OAI221XL U198 ( .A0(n172), .A1(n18), .B0(n27), .B1(n83), .C0(n253), .Y(n251)
         );
  AOI2BB2X1 U199 ( .B0(n65), .B1(n24), .A0N(n169), .A1N(n20), .Y(n253) );
  NAND2X1 U200 ( .A(n199), .B(n204), .Y(n169) );
  NAND2X1 U201 ( .A(n200), .B(n106), .Y(n83) );
  INVX1 U202 ( .A(n211), .Y(n106) );
  AOI221X1 U203 ( .A0(n211), .A1(n5), .B0(n40), .B1(a[4]), .C0(n254), .Y(n248)
         );
  MXI2X1 U204 ( .A(n255), .B(n256), .S0(n252), .Y(n254) );
  NOR3X1 U205 ( .A(n257), .B(n258), .C(n50), .Y(n256) );
  OAI22X1 U206 ( .A0(n20), .A1(n68), .B0(n27), .B1(n37), .Y(n257) );
  AOI211X1 U207 ( .A0(n259), .A1(n24), .B0(n260), .C0(n261), .Y(n255) );
  INVX1 U208 ( .A(n262), .Y(n261) );
  NOR2X1 U209 ( .A(n94), .B(a[1]), .Y(n211) );
  MXI2X1 U210 ( .A(n263), .B(n264), .S0(a[6]), .Y(d[2]) );
  AOI211X1 U211 ( .A0(n55), .A1(n265), .B0(n266), .C0(n267), .Y(n264) );
  INVX1 U212 ( .A(n268), .Y(n267) );
  OAI31X1 U213 ( .A0(n176), .A1(n269), .A2(n270), .B0(n16), .Y(n268) );
  OAI21XL U214 ( .A0(n4), .A1(n271), .B0(n272), .Y(n270) );
  NOR2X1 U215 ( .A(n20), .B(n226), .Y(n176) );
  OAI22X1 U216 ( .A0(n273), .A1(n10), .B0(n274), .B1(n52), .Y(n266) );
  MXI2X1 U217 ( .A(n276), .B(n277), .S0(n155), .Y(n275) );
  XNOR2X1 U218 ( .A(n129), .B(a[1]), .Y(n155) );
  NAND2X1 U219 ( .A(a[2]), .B(n149), .Y(n276) );
  OAI221XL U220 ( .A0(a[1]), .A1(n247), .B0(n4), .B1(n189), .C0(n272), .Y(n279) );
  NAND2X1 U221 ( .A(n41), .B(n33), .Y(n272) );
  INVX1 U222 ( .A(n280), .Y(n247) );
  OAI221XL U223 ( .A0(n281), .A1(n27), .B0(n4), .B1(n111), .C0(n282), .Y(n265)
         );
  AOI211X1 U224 ( .A0(n5), .A1(n125), .B0(n50), .C0(n283), .Y(n282) );
  AOI21X1 U225 ( .A0(n200), .A1(n223), .B0(n20), .Y(n283) );
  NOR2X1 U226 ( .A(n199), .B(n4), .Y(n50) );
  NAND2X1 U227 ( .A(n284), .B(n122), .Y(n125) );
  AOI211X1 U228 ( .A0(n285), .A1(n55), .B0(n286), .C0(n287), .Y(n263) );
  AOI31X1 U229 ( .A0(n132), .A1(n288), .A2(n289), .B0(n52), .Y(n287) );
  AOI22X1 U230 ( .A0(n102), .A1(n69), .B0(n184), .B1(n33), .Y(n289) );
  NOR2X1 U231 ( .A(n290), .B(n163), .Y(n184) );
  NAND2X1 U232 ( .A(n200), .B(n284), .Y(n102) );
  INVX1 U233 ( .A(n225), .Y(n288) );
  OAI22X1 U234 ( .A0(n291), .A1(n114), .B0(n292), .B1(n10), .Y(n286) );
  INVX1 U235 ( .A(n89), .Y(n10) );
  AOI211X1 U236 ( .A0(n5), .A1(n79), .B0(n293), .C0(n294), .Y(n292) );
  AOI21X1 U237 ( .A0(n101), .A1(n150), .B0(n20), .Y(n294) );
  OAI2BB2X1 U238 ( .B0(n27), .B1(n295), .A0N(n34), .A1N(n24), .Y(n293) );
  OAI221XL U239 ( .A0(n298), .A1(n27), .B0(n20), .B1(n122), .C0(n132), .Y(n297) );
  NOR2X1 U240 ( .A(n159), .B(n217), .Y(n198) );
  NAND2X1 U241 ( .A(a[1]), .B(n47), .Y(n122) );
  NOR2X1 U242 ( .A(n299), .B(n242), .Y(n298) );
  INVX1 U243 ( .A(n99), .Y(n296) );
  NAND2X1 U244 ( .A(n200), .B(n300), .Y(n99) );
  MXI2X1 U245 ( .A(n301), .B(n147), .S0(n302), .Y(n285) );
  MXI2X1 U246 ( .A(n303), .B(n61), .S0(n69), .Y(n301) );
  INVX1 U247 ( .A(n187), .Y(n61) );
  MX2X1 U248 ( .A(n304), .B(n305), .S0(a[6]), .Y(d[1]) );
  OAI221XL U249 ( .A0(n306), .A1(n52), .B0(n307), .B1(n114), .C0(n308), .Y(
        n305) );
  AOI22X1 U250 ( .A0(n89), .A1(n309), .B0(n55), .B1(n310), .Y(n308) );
  OAI221XL U251 ( .A0(n27), .A1(n44), .B0(n4), .B1(n48), .C0(n311), .Y(n310)
         );
  AND2X1 U252 ( .A(n223), .B(n240), .Y(n28) );
  INVX1 U253 ( .A(n185), .Y(n48) );
  AOI21X1 U254 ( .A0(n226), .A1(n188), .B0(n242), .Y(n185) );
  OAI221XL U255 ( .A0(n149), .A1(n20), .B0(n4), .B1(n227), .C0(n312), .Y(n309)
         );
  AOI21X1 U256 ( .A0(n313), .A1(n33), .B0(n269), .Y(n312) );
  NAND2X1 U257 ( .A(n284), .B(n105), .Y(n227) );
  INVX1 U258 ( .A(n41), .Y(n105) );
  NOR2X1 U259 ( .A(n149), .B(n226), .Y(n41) );
  OAI22X1 U260 ( .A0(n92), .A1(n18), .B0(n316), .B1(n27), .Y(n315) );
  AOI21X1 U261 ( .A0(a[1]), .A1(n58), .B0(n98), .Y(n316) );
  INVX1 U262 ( .A(n295), .Y(n92) );
  NOR2X1 U263 ( .A(n45), .B(n163), .Y(n160) );
  INVX1 U264 ( .A(n151), .Y(n314) );
  NAND2X1 U265 ( .A(n100), .B(n199), .Y(n151) );
  AOI211X1 U266 ( .A0(n33), .A1(n120), .B0(n317), .C0(n318), .Y(n306) );
  INVX1 U267 ( .A(n258), .Y(n182) );
  OAI221XL U268 ( .A0(n20), .A1(n100), .B0(a[3]), .B1(n4), .C0(n262), .Y(n317)
         );
  INVX1 U269 ( .A(n210), .Y(n100) );
  NAND2X1 U270 ( .A(n34), .B(n200), .Y(n120) );
  INVX1 U271 ( .A(n290), .Y(n200) );
  NOR2X1 U272 ( .A(n226), .B(n58), .Y(n290) );
  OAI221XL U273 ( .A0(n319), .A1(n52), .B0(n320), .B1(n114), .C0(n321), .Y(
        n304) );
  AOI22X1 U274 ( .A0(n55), .A1(n322), .B0(n89), .B1(n323), .Y(n321) );
  OAI221XL U275 ( .A0(n47), .A1(n27), .B0(n65), .B1(n20), .C0(n324), .Y(n323)
         );
  AOI21X1 U276 ( .A0(n40), .A1(a[4]), .B0(n135), .Y(n324) );
  NOR2X1 U277 ( .A(n71), .B(n18), .Y(n135) );
  NAND2X1 U278 ( .A(n19), .B(n189), .Y(n71) );
  OAI21XL U279 ( .A0(n325), .A1(n18), .B0(n326), .Y(n322) );
  AOI31X1 U280 ( .A0(n111), .A1(n149), .A2(n327), .B0(n225), .Y(n326) );
  OAI21XL U281 ( .A0(n69), .A1(n284), .B0(n27), .Y(n327) );
  INVX1 U282 ( .A(n98), .Y(n284) );
  NOR2X1 U283 ( .A(n47), .B(a[1]), .Y(n98) );
  INVX1 U284 ( .A(n145), .Y(n149) );
  INVX1 U285 ( .A(n16), .Y(n114) );
  NOR2X1 U286 ( .A(a[0]), .B(a[5]), .Y(n16) );
  OAI32X1 U287 ( .A0(n4), .A1(n145), .A2(n210), .B0(n137), .B1(n27), .Y(n328)
         );
  AND2X1 U288 ( .A(n300), .B(n240), .Y(n23) );
  NAND2X1 U289 ( .A(n44), .B(n226), .Y(n300) );
  NOR2X1 U290 ( .A(n25), .B(n299), .Y(n313) );
  NOR2X1 U291 ( .A(n234), .B(a[5]), .Y(n14) );
  AOI221X1 U292 ( .A0(n325), .A1(n33), .B0(n24), .B1(n303), .C0(n329), .Y(n319) );
  OAI221XL U293 ( .A0(n18), .A1(n330), .B0(n20), .B1(n80), .C0(n75), .Y(n329)
         );
  INVX1 U294 ( .A(n269), .Y(n75) );
  NOR2X1 U295 ( .A(n111), .B(n18), .Y(n269) );
  INVX1 U296 ( .A(n299), .Y(n80) );
  MX4X1 U297 ( .A(n331), .B(n332), .C(n333), .D(n334), .S0(a[6]), .S1(n234), 
        .Y(d[0]) );
  NOR2X1 U298 ( .A(n258), .B(n335), .Y(n334) );
  MXI2X1 U299 ( .A(n336), .B(n337), .S0(n252), .Y(n335) );
  OAI21XL U300 ( .A0(n4), .A1(n121), .B0(n339), .Y(n338) );
  NOR2X1 U301 ( .A(n18), .B(n136), .Y(n280) );
  NAND2X1 U302 ( .A(n126), .B(n101), .Y(n178) );
  INVX1 U303 ( .A(n45), .Y(n126) );
  OAI32X1 U304 ( .A0(n27), .A1(n278), .A2(n95), .B0(n341), .B1(n4), .Y(n340)
         );
  NOR2X1 U305 ( .A(n299), .B(n210), .Y(n341) );
  NOR2X1 U306 ( .A(n136), .B(a[1]), .Y(n299) );
  NAND2X1 U307 ( .A(n204), .B(n330), .Y(n239) );
  INVX1 U308 ( .A(n179), .Y(n330) );
  NOR2X1 U309 ( .A(n188), .B(a[1]), .Y(n179) );
  NAND2X1 U310 ( .A(n278), .B(a[1]), .Y(n204) );
  NOR2X1 U311 ( .A(n18), .B(n226), .Y(n258) );
  AOI211X1 U312 ( .A0(n5), .A1(n68), .B0(n342), .C0(n343), .Y(n333) );
  AOI21X1 U313 ( .A0(n240), .A1(n37), .B0(n344), .Y(n343) );
  INVX1 U314 ( .A(n173), .Y(n344) );
  INVX1 U315 ( .A(n163), .Y(n37) );
  NOR2X1 U316 ( .A(a[1]), .B(a[3]), .Y(n163) );
  MXI2X1 U317 ( .A(n345), .B(n346), .S0(n252), .Y(n342) );
  NOR2X1 U318 ( .A(n27), .B(n210), .Y(n173) );
  NOR2X1 U319 ( .A(n226), .B(n259), .Y(n210) );
  NAND2X1 U320 ( .A(n19), .B(n199), .Y(n295) );
  NAND2X1 U321 ( .A(n199), .B(n205), .Y(n82) );
  NAND2X1 U322 ( .A(n94), .B(n226), .Y(n199) );
  INVX1 U323 ( .A(n278), .Y(n94) );
  NOR2X1 U324 ( .A(n225), .B(n40), .Y(n345) );
  NOR2X1 U325 ( .A(n20), .B(n159), .Y(n225) );
  NAND2X1 U326 ( .A(n240), .B(n189), .Y(n68) );
  INVX1 U327 ( .A(n157), .Y(n240) );
  NOR2X1 U328 ( .A(n44), .B(n226), .Y(n157) );
  MXI2X1 U329 ( .A(n347), .B(n348), .S0(n252), .Y(n332) );
  OAI211X1 U330 ( .A0(n349), .A1(n74), .B0(n350), .C0(n351), .Y(n348) );
  NAND2X1 U331 ( .A(n278), .B(n6), .Y(n74) );
  INVX1 U332 ( .A(n352), .Y(n349) );
  OAI221XL U333 ( .A0(n20), .A1(n34), .B0(n325), .B1(n4), .C0(n353), .Y(n347)
         );
  AOI31X1 U334 ( .A0(n6), .A1(n352), .A2(n259), .B0(n354), .Y(n353) );
  AOI21X1 U335 ( .A0(n19), .A1(n223), .B0(n27), .Y(n354) );
  NAND2X1 U336 ( .A(n145), .B(n226), .Y(n223) );
  INVX1 U337 ( .A(n281), .Y(n19) );
  NOR2X1 U338 ( .A(n226), .B(n136), .Y(n281) );
  XNOR2X1 U339 ( .A(a[5]), .B(n226), .Y(n352) );
  AND2X1 U340 ( .A(n101), .B(n79), .Y(n325) );
  INVX1 U341 ( .A(n59), .Y(n79) );
  MXI2X1 U342 ( .A(n355), .B(n356), .S0(n252), .Y(n331) );
  OAI221XL U343 ( .A0(n18), .A1(n121), .B0(n271), .B1(n20), .C0(n357), .Y(n356) );
  AOI22X1 U344 ( .A0(n33), .A1(n147), .B0(n24), .B1(n107), .Y(n357) );
  INVX1 U345 ( .A(n172), .Y(n107) );
  NOR2X1 U346 ( .A(n188), .B(n226), .Y(n25) );
  INVX1 U347 ( .A(n159), .Y(n188) );
  NAND2X1 U348 ( .A(a[4]), .B(n226), .Y(n101) );
  NAND2X1 U349 ( .A(n44), .B(n150), .Y(n147) );
  INVX1 U350 ( .A(n217), .Y(n150) );
  NOR2X1 U351 ( .A(n226), .B(n278), .Y(n217) );
  NOR2X1 U352 ( .A(n96), .B(n59), .Y(n271) );
  NOR2X1 U353 ( .A(n226), .B(n145), .Y(n59) );
  OAI211X1 U354 ( .A0(n65), .A1(n27), .B0(n158), .C0(n358), .Y(n355) );
  INVX1 U355 ( .A(n47), .Y(n96) );
  INVX1 U356 ( .A(n42), .Y(n121) );
  NOR2X1 U357 ( .A(n145), .B(a[1]), .Y(n42) );
  INVX1 U358 ( .A(n95), .Y(n111) );
  NOR2X1 U359 ( .A(n226), .B(n159), .Y(n95) );
  NAND2BX1 U360 ( .AN(n73), .B(n6), .Y(n158) );
  NOR2X1 U361 ( .A(n259), .B(n45), .Y(n73) );
  NOR2X1 U362 ( .A(n226), .B(n47), .Y(n45) );
  AND2X1 U363 ( .A(n189), .B(n205), .Y(n65) );
  INVX1 U364 ( .A(n242), .Y(n205) );
  NOR2X1 U365 ( .A(n226), .B(a[3]), .Y(n242) );
  NAND2X1 U366 ( .A(n47), .B(n226), .Y(n189) );
endmodule


module aes_sbox_2 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358;

  AOI31XL U1 ( .A0(n79), .A1(n44), .A2(n2), .B0(n280), .Y(n339) );
  AOI31X1 U2 ( .A0(n44), .A1(n129), .A2(n130), .B0(n131), .Y(n128) );
  AOI221X1 U3 ( .A0(n40), .A1(n136), .B0(n33), .B1(n47), .C0(n156), .Y(n141)
         );
  OAI32X1 U4 ( .A0(n210), .A1(n145), .A2(n18), .B0(n27), .B1(n211), .Y(n209)
         );
  AOI222XL U5 ( .A0(n59), .A1(n43), .B0(n6), .B1(n221), .C0(n222), .C1(n187), 
        .Y(n218) );
  AOI221X1 U6 ( .A0(n278), .A1(n40), .B0(n185), .B1(n2), .C0(n279), .Y(n273)
         );
  AOI221X1 U7 ( .A0(n225), .A1(n226), .B0(n296), .B1(n6), .C0(n297), .Y(n291)
         );
  OAI32X1 U8 ( .A0(n18), .A1(a[1]), .A2(n159), .B0(a[4]), .B1(n182), .Y(n318)
         );
  AOI221XL U9 ( .A0(n314), .A1(n43), .B0(n160), .B1(n24), .C0(n315), .Y(n307)
         );
  AOI221X1 U10 ( .A0(n313), .A1(n5), .B0(n23), .B1(n2), .C0(n328), .Y(n320) );
  AOI31X1 U11 ( .A0(a[2]), .A1(n58), .A2(a[1]), .B0(n40), .Y(n350) );
  AOI222XL U12 ( .A0(n278), .A1(n24), .B0(n42), .B1(n33), .C0(n43), .C1(n136), 
        .Y(n351) );
  AOI221XL U13 ( .A0(n5), .A1(n96), .B0(n43), .B1(n239), .C0(n340), .Y(n336)
         );
  AOI221X1 U14 ( .A0(n40), .A1(n136), .B0(n33), .B1(n178), .C0(n338), .Y(n337)
         );
  OR2X2 U15 ( .A(a[2]), .B(a[7]), .Y(n1) );
  AOI221X1 U16 ( .A0(n5), .A1(n19), .B0(n33), .B1(n34), .C0(n35), .Y(n11) );
  OAI222X1 U17 ( .A0(n4), .A1(n37), .B0(n38), .B1(n20), .C0(a[4]), .C1(n39), 
        .Y(n35) );
  OAI222X1 U18 ( .A0(n20), .A1(n99), .B0(n27), .B1(n101), .C0(n184), .C1(n4), 
        .Y(n250) );
  OAI222X1 U19 ( .A0(n27), .A1(n34), .B0(n69), .B1(n205), .C0(n20), .C1(n79), 
        .Y(n260) );
  NAND2X2 U20 ( .A(n58), .B(n226), .Y(n34) );
  NOR2BXL U21 ( .AN(n101), .B(n25), .Y(n172) );
  AOI221XL U22 ( .A0(n43), .A1(n151), .B0(n25), .B1(n69), .C0(n275), .Y(n274)
         );
  NAND2XL U23 ( .A(n111), .B(n121), .Y(n303) );
  NAND2XL U24 ( .A(n111), .B(n300), .Y(n187) );
  NAND2XL U25 ( .A(n111), .B(n101), .Y(n21) );
  OAI2BB2XL U26 ( .B0(n20), .B1(n111), .A0N(n125), .A1N(n24), .Y(n220) );
  NAND2XL U27 ( .A(n198), .B(n24), .Y(n132) );
  AOI22XL U28 ( .A0(n33), .A1(a[3]), .B0(n24), .B1(n58), .Y(n277) );
  AOI22XL U29 ( .A0(n23), .A1(n24), .B0(n25), .B1(a[2]), .Y(n22) );
  AOI21XL U30 ( .A0(n44), .A1(n111), .B0(n4), .Y(n177) );
  NOR2X2 U31 ( .A(n44), .B(a[1]), .Y(n137) );
  CLKINVX3 U32 ( .A(n259), .Y(n44) );
  NOR2X2 U33 ( .A(n259), .B(n278), .Y(n47) );
  NOR2X2 U34 ( .A(a[4]), .B(a[3]), .Y(n278) );
  NOR2X2 U35 ( .A(n136), .B(n58), .Y(n259) );
  NOR2X2 U36 ( .A(n58), .B(a[3]), .Y(n159) );
  CLKINVX3 U37 ( .A(a[4]), .Y(n58) );
  NOR2X2 U38 ( .A(n136), .B(a[4]), .Y(n145) );
  CLKINVX3 U39 ( .A(a[3]), .Y(n136) );
  NOR2X4 U40 ( .A(n226), .B(n4), .Y(n40) );
  INVX4 U41 ( .A(a[2]), .Y(n69) );
  AOI21XL U42 ( .A0(n18), .A1(n162), .B0(n25), .Y(n161) );
  INVX4 U43 ( .A(n6), .Y(n18) );
  INVXL U44 ( .A(n20), .Y(n2) );
  MXI2XL U45 ( .A(n2), .B(n6), .S0(n28), .Y(n311) );
  NOR2XL U46 ( .A(n33), .B(n2), .Y(n302) );
  AOI22XL U47 ( .A0(n184), .A1(n5), .B0(n198), .B1(n43), .Y(n197) );
  AOI22XL U48 ( .A0(n40), .A1(n94), .B0(n43), .B1(n187), .Y(n244) );
  AOI21XL U49 ( .A0(n159), .A1(n43), .B0(n40), .Y(n262) );
  AOI22XL U50 ( .A0(n43), .A1(n100), .B0(n24), .B1(n125), .Y(n124) );
  AOI22XL U51 ( .A0(n43), .A1(n303), .B0(n24), .B1(n96), .Y(n358) );
  AOI222X4 U52 ( .A0(n125), .A1(n33), .B0(n145), .B1(n40), .C0(n43), .C1(n184), 
        .Y(n183) );
  AOI2BB2XL U53 ( .B0(n43), .B1(n94), .A0N(n120), .A1N(n4), .Y(n119) );
  AOI22XL U54 ( .A0(n82), .A1(n43), .B0(n83), .B1(n24), .Y(n81) );
  AOI22XL U55 ( .A0(n98), .A1(n43), .B0(n6), .B1(n99), .Y(n97) );
  AOI22XL U56 ( .A0(n217), .A1(n43), .B0(n33), .B1(n47), .Y(n216) );
  AOI221X4 U57 ( .A0(n43), .A1(n44), .B0(n45), .B1(n24), .C0(n46), .Y(n9) );
  AOI221X4 U58 ( .A0(n43), .A1(n205), .B0(n32), .B1(n6), .C0(n206), .Y(n201)
         );
  AOI221X4 U59 ( .A0(n43), .A1(n208), .B0(n76), .B1(n24), .C0(n209), .Y(n207)
         );
  AOI221X4 U60 ( .A0(n70), .A1(n43), .B0(n24), .B1(n71), .C0(n72), .Y(n53) );
  AOI222X4 U61 ( .A0(n185), .A1(n43), .B0(n186), .B1(n187), .C0(n6), .C1(n188), 
        .Y(n164) );
  AOI222X4 U62 ( .A0(n123), .A1(n43), .B0(a[2]), .B1(n203), .C0(n6), .C1(n71), 
        .Y(n202) );
  AOI221X4 U63 ( .A0(n59), .A1(n33), .B0(n43), .B1(n126), .C0(n127), .Y(n113)
         );
  AOI221X4 U64 ( .A0(n24), .A1(n82), .B0(n43), .B1(n295), .C0(n173), .Y(n346)
         );
  INVX4 U65 ( .A(n43), .Y(n20) );
  INVXL U66 ( .A(n36), .Y(n3) );
  INVX4 U67 ( .A(n3), .Y(n4) );
  INVXL U68 ( .A(n24), .Y(n36) );
  CLKINVX3 U69 ( .A(n1), .Y(n5) );
  CLKINVX3 U70 ( .A(n1), .Y(n6) );
  INVX12 U71 ( .A(n33), .Y(n27) );
  NOR2X4 U72 ( .A(n69), .B(a[7]), .Y(n33) );
  CLKINVX3 U73 ( .A(a[0]), .Y(n234) );
  NOR2X2 U74 ( .A(n252), .B(a[0]), .Y(n89) );
  AOI22XL U75 ( .A0(n70), .A1(n24), .B0(n96), .B1(n129), .Y(n241) );
  NOR2X4 U76 ( .A(n129), .B(n69), .Y(n24) );
  CLKINVX3 U77 ( .A(a[7]), .Y(n129) );
  NOR2X2 U78 ( .A(n252), .B(n234), .Y(n55) );
  CLKINVX3 U79 ( .A(a[5]), .Y(n252) );
  AOI22XL U80 ( .A0(n225), .A1(n226), .B0(n6), .B1(n227), .Y(n224) );
  INVX4 U81 ( .A(a[1]), .Y(n226) );
  OAI22XL U82 ( .A0(n201), .A1(n52), .B0(n202), .B1(n114), .Y(n193) );
  CLKINVX3 U83 ( .A(n14), .Y(n52) );
  NOR2X4 U84 ( .A(n129), .B(a[2]), .Y(n43) );
  MX2X1 U85 ( .A(n7), .B(n8), .S0(a[6]), .Y(d[7]) );
  OAI221XL U86 ( .A0(n9), .A1(n10), .B0(n11), .B1(n12), .C0(n13), .Y(n8) );
  AOI22X1 U87 ( .A0(n14), .A1(n15), .B0(n16), .B1(n17), .Y(n13) );
  OAI221XL U88 ( .A0(n18), .A1(n19), .B0(n20), .B1(n21), .C0(n22), .Y(n17) );
  OAI221XL U89 ( .A0(n26), .A1(n27), .B0(n28), .B1(n20), .C0(n29), .Y(n15) );
  AOI21X1 U90 ( .A0(n5), .A1(n30), .B0(n31), .Y(n29) );
  INVX1 U91 ( .A(n32), .Y(n26) );
  INVX1 U92 ( .A(n40), .Y(n39) );
  NOR2X1 U93 ( .A(n41), .B(n42), .Y(n38) );
  OAI221XL U94 ( .A0(n47), .A1(n18), .B0(n27), .B1(n48), .C0(n49), .Y(n46) );
  INVX1 U95 ( .A(n50), .Y(n49) );
  OAI221XL U96 ( .A0(n51), .A1(n52), .B0(n53), .B1(n10), .C0(n54), .Y(n7) );
  AOI22X1 U97 ( .A0(n55), .A1(n56), .B0(n16), .B1(n57), .Y(n54) );
  OAI221XL U98 ( .A0(n58), .A1(n18), .B0(n59), .B1(n27), .C0(n60), .Y(n57) );
  AOI2BB2X1 U99 ( .B0(n61), .B1(n24), .A0N(n62), .A1N(n20), .Y(n60) );
  OAI221XL U100 ( .A0(n63), .A1(n64), .B0(n65), .B1(n27), .C0(n66), .Y(n56) );
  INVX1 U101 ( .A(n67), .Y(n66) );
  AOI21X1 U102 ( .A0(n68), .A1(n69), .B0(n6), .Y(n63) );
  OAI211X1 U103 ( .A0(n73), .A1(n27), .B0(n74), .C0(n75), .Y(n72) );
  AOI211X1 U104 ( .A0(n5), .A1(n76), .B0(n77), .C0(n78), .Y(n51) );
  AOI21X1 U105 ( .A0(n79), .A1(n80), .B0(n27), .Y(n78) );
  INVX1 U106 ( .A(n81), .Y(n77) );
  MX2X1 U107 ( .A(n84), .B(n85), .S0(a[6]), .Y(d[6]) );
  OAI221XL U108 ( .A0(n86), .A1(n52), .B0(n87), .B1(n12), .C0(n88), .Y(n85) );
  AOI22X1 U109 ( .A0(n89), .A1(n90), .B0(n16), .B1(n91), .Y(n88) );
  OAI221XL U110 ( .A0(n73), .A1(n27), .B0(n92), .B1(n20), .C0(n93), .Y(n91) );
  AOI31X1 U111 ( .A0(n79), .A1(n94), .A2(n6), .B0(n67), .Y(n93) );
  NOR3X1 U112 ( .A(n4), .B(n95), .C(n96), .Y(n67) );
  OAI221XL U113 ( .A0(n27), .A1(n62), .B0(n4), .B1(n21), .C0(n97), .Y(n90) );
  NAND2X1 U114 ( .A(n100), .B(n101), .Y(n62) );
  AOI211X1 U115 ( .A0(n33), .A1(n102), .B0(n103), .C0(n104), .Y(n87) );
  AOI21X1 U116 ( .A0(n105), .A1(n106), .B0(n20), .Y(n104) );
  OAI22X1 U117 ( .A0(n45), .A1(n4), .B0(a[4]), .B1(n18), .Y(n103) );
  AOI211X1 U118 ( .A0(n5), .A1(n107), .B0(n108), .C0(n109), .Y(n86) );
  AOI21X1 U119 ( .A0(a[1]), .A1(n58), .B0(n27), .Y(n109) );
  OAI22X1 U120 ( .A0(n110), .A1(n4), .B0(n20), .B1(n21), .Y(n108) );
  OAI221XL U121 ( .A0(n112), .A1(n52), .B0(n113), .B1(n114), .C0(n115), .Y(n84) );
  AOI22X1 U122 ( .A0(n89), .A1(n116), .B0(n55), .B1(n117), .Y(n115) );
  OAI221XL U123 ( .A0(n18), .A1(n118), .B0(n27), .B1(n30), .C0(n119), .Y(n117)
         );
  NAND2X1 U124 ( .A(n121), .B(n122), .Y(n30) );
  OAI221XL U125 ( .A0(n18), .A1(n105), .B0(n123), .B1(n27), .C0(n124), .Y(n116) );
  OAI21XL U126 ( .A0(n18), .A1(n37), .B0(n128), .Y(n127) );
  INVX1 U127 ( .A(n132), .Y(n131) );
  AOI211X1 U128 ( .A0(n133), .A1(n69), .B0(n134), .C0(n135), .Y(n112) );
  OAI22X1 U129 ( .A0(n4), .A1(n136), .B0(n137), .B1(n27), .Y(n134) );
  INVX1 U130 ( .A(n70), .Y(n133) );
  MX2X1 U131 ( .A(n138), .B(n139), .S0(a[6]), .Y(d[5]) );
  OAI221XL U132 ( .A0(n140), .A1(n12), .B0(n141), .B1(n114), .C0(n142), .Y(
        n139) );
  AOI22X1 U133 ( .A0(n89), .A1(n143), .B0(n14), .B1(n144), .Y(n142) );
  OAI221XL U134 ( .A0(n145), .A1(n20), .B0(n4), .B1(n34), .C0(n146), .Y(n144)
         );
  AOI2BB1X1 U135 ( .A0N(n147), .A1N(n27), .B0(n148), .Y(n146) );
  AOI21X1 U136 ( .A0(n149), .A1(n150), .B0(n18), .Y(n148) );
  OAI221XL U137 ( .A0(n110), .A1(n18), .B0(n20), .B1(n151), .C0(n152), .Y(n143) );
  MXI2X1 U138 ( .A(n153), .B(n154), .S0(n155), .Y(n152) );
  NOR2X1 U139 ( .A(n145), .B(n69), .Y(n154) );
  NOR2X1 U140 ( .A(n4), .B(n136), .Y(n153) );
  OAI21XL U141 ( .A0(n157), .A1(n20), .B0(n158), .Y(n156) );
  AOI221X1 U142 ( .A0(n159), .A1(n24), .B0(n160), .B1(n33), .C0(n161), .Y(n140) );
  OAI21XL U143 ( .A0(n41), .A1(n163), .B0(n69), .Y(n162) );
  OAI221XL U144 ( .A0(n164), .A1(n114), .B0(n165), .B1(n52), .C0(n166), .Y(
        n138) );
  AOI22X1 U145 ( .A0(n89), .A1(n167), .B0(n55), .B1(n168), .Y(n166) );
  OAI211X1 U146 ( .A0(n20), .A1(n169), .B0(n170), .C0(n171), .Y(n168) );
  AOI22X1 U147 ( .A0(n137), .A1(n24), .B0(n172), .B1(n6), .Y(n171) );
  MXI2X1 U148 ( .A(n40), .B(n173), .S0(n96), .Y(n170) );
  OAI221XL U149 ( .A0(n159), .A1(n27), .B0(n145), .B1(n20), .C0(n174), .Y(n167) );
  AOI211X1 U150 ( .A0(n175), .A1(n5), .B0(n176), .C0(n177), .Y(n174) );
  INVX1 U151 ( .A(n178), .Y(n175) );
  AOI211X1 U152 ( .A0(n179), .A1(n24), .B0(n180), .C0(n181), .Y(n165) );
  NAND2X1 U153 ( .A(n74), .B(n182), .Y(n181) );
  INVX1 U154 ( .A(n183), .Y(n180) );
  OAI21XL U155 ( .A0(n69), .A1(n189), .B0(n27), .Y(n186) );
  MXI2X1 U156 ( .A(n190), .B(n191), .S0(a[6]), .Y(d[4]) );
  AOI211X1 U157 ( .A0(n89), .A1(n192), .B0(n193), .C0(n194), .Y(n191) );
  AOI31X1 U158 ( .A0(n195), .A1(n196), .A2(n197), .B0(n12), .Y(n194) );
  INVX1 U159 ( .A(n55), .Y(n12) );
  OAI2BB1X1 U160 ( .A0N(n199), .A1N(n200), .B0(n33), .Y(n195) );
  NAND2X1 U161 ( .A(n94), .B(n79), .Y(n203) );
  INVX1 U162 ( .A(n118), .Y(n123) );
  NAND2X1 U163 ( .A(n204), .B(n80), .Y(n118) );
  OAI22X1 U164 ( .A0(n28), .A1(n4), .B0(n188), .B1(n27), .Y(n206) );
  NOR2X1 U165 ( .A(n25), .B(n98), .Y(n32) );
  INVX1 U166 ( .A(n207), .Y(n192) );
  AOI211X1 U167 ( .A0(n55), .A1(n212), .B0(n213), .C0(n214), .Y(n190) );
  AOI31X1 U168 ( .A0(n215), .A1(n196), .A2(n216), .B0(n52), .Y(n214) );
  INVX1 U169 ( .A(n31), .Y(n196) );
  NOR2X1 U170 ( .A(n4), .B(n159), .Y(n31) );
  INVX1 U171 ( .A(n135), .Y(n215) );
  OAI22X1 U172 ( .A0(n218), .A1(n10), .B0(n219), .B1(n114), .Y(n213) );
  AOI211X1 U173 ( .A0(n208), .A1(n5), .B0(n220), .C0(n173), .Y(n219) );
  NOR2X1 U174 ( .A(n217), .B(n42), .Y(n208) );
  OAI21XL U175 ( .A0(n69), .A1(n223), .B0(n27), .Y(n222) );
  NAND2X1 U176 ( .A(n34), .B(n204), .Y(n221) );
  OAI221XL U177 ( .A0(n27), .A1(n64), .B0(n4), .B1(n83), .C0(n224), .Y(n212)
         );
  INVX1 U178 ( .A(n110), .Y(n64) );
  NOR2BX1 U179 ( .AN(n204), .B(n137), .Y(n110) );
  MX2X1 U180 ( .A(n228), .B(n229), .S0(a[6]), .Y(d[3]) );
  MX4X1 U181 ( .A(n230), .B(n231), .C(n232), .D(n233), .S0(n234), .S1(a[5]), 
        .Y(n229) );
  OAI211X1 U182 ( .A0(n27), .A1(n122), .B0(n158), .C0(n235), .Y(n233) );
  AOI2BB2X1 U183 ( .B0(n24), .B1(n187), .A0N(n227), .A1N(n20), .Y(n235) );
  OAI221XL U184 ( .A0(n18), .A1(n76), .B0(n59), .B1(n27), .C0(n236), .Y(n232)
         );
  OAI21XL U185 ( .A0(n237), .A1(n43), .B0(n238), .Y(n236) );
  INVX1 U186 ( .A(n239), .Y(n238) );
  AOI21X1 U187 ( .A0(n122), .A1(n106), .B0(n129), .Y(n237) );
  NAND2X1 U188 ( .A(n101), .B(n240), .Y(n76) );
  OAI221XL U189 ( .A0(n159), .A1(n27), .B0(n20), .B1(n34), .C0(n241), .Y(n231)
         );
  NOR2X1 U190 ( .A(n242), .B(n137), .Y(n70) );
  OAI211X1 U191 ( .A0(n4), .A1(n149), .B0(n243), .C0(n244), .Y(n230) );
  MXI2X1 U192 ( .A(n245), .B(n246), .S0(n130), .Y(n243) );
  XNOR2X1 U193 ( .A(n69), .B(a[1]), .Y(n130) );
  NOR2X1 U194 ( .A(a[7]), .B(n145), .Y(n246) );
  OAI21XL U195 ( .A0(n58), .A1(n27), .B0(n247), .Y(n245) );
  MXI2X1 U196 ( .A(n248), .B(n249), .S0(n234), .Y(n228) );
  MXI2X1 U197 ( .A(n250), .B(n251), .S0(n252), .Y(n249) );
  OAI221XL U198 ( .A0(n172), .A1(n18), .B0(n27), .B1(n83), .C0(n253), .Y(n251)
         );
  AOI2BB2X1 U199 ( .B0(n65), .B1(n24), .A0N(n169), .A1N(n20), .Y(n253) );
  NAND2X1 U200 ( .A(n199), .B(n204), .Y(n169) );
  NAND2X1 U201 ( .A(n200), .B(n106), .Y(n83) );
  INVX1 U202 ( .A(n211), .Y(n106) );
  AOI221X1 U203 ( .A0(n211), .A1(n5), .B0(n40), .B1(a[4]), .C0(n254), .Y(n248)
         );
  MXI2X1 U204 ( .A(n255), .B(n256), .S0(n252), .Y(n254) );
  NOR3X1 U205 ( .A(n257), .B(n258), .C(n50), .Y(n256) );
  OAI22X1 U206 ( .A0(n20), .A1(n68), .B0(n27), .B1(n37), .Y(n257) );
  AOI211X1 U207 ( .A0(n259), .A1(n24), .B0(n260), .C0(n261), .Y(n255) );
  INVX1 U208 ( .A(n262), .Y(n261) );
  NOR2X1 U209 ( .A(n94), .B(a[1]), .Y(n211) );
  MXI2X1 U210 ( .A(n263), .B(n264), .S0(a[6]), .Y(d[2]) );
  AOI211X1 U211 ( .A0(n55), .A1(n265), .B0(n266), .C0(n267), .Y(n264) );
  INVX1 U212 ( .A(n268), .Y(n267) );
  OAI31X1 U213 ( .A0(n176), .A1(n269), .A2(n270), .B0(n16), .Y(n268) );
  OAI21XL U214 ( .A0(n4), .A1(n271), .B0(n272), .Y(n270) );
  NOR2X1 U215 ( .A(n20), .B(n226), .Y(n176) );
  OAI22X1 U216 ( .A0(n273), .A1(n10), .B0(n274), .B1(n52), .Y(n266) );
  MXI2X1 U217 ( .A(n276), .B(n277), .S0(n155), .Y(n275) );
  XNOR2X1 U218 ( .A(n129), .B(a[1]), .Y(n155) );
  NAND2X1 U219 ( .A(a[2]), .B(n149), .Y(n276) );
  OAI221XL U220 ( .A0(a[1]), .A1(n247), .B0(n4), .B1(n189), .C0(n272), .Y(n279) );
  NAND2X1 U221 ( .A(n41), .B(n33), .Y(n272) );
  INVX1 U222 ( .A(n280), .Y(n247) );
  OAI221XL U223 ( .A0(n281), .A1(n27), .B0(n4), .B1(n111), .C0(n282), .Y(n265)
         );
  AOI211X1 U224 ( .A0(n5), .A1(n125), .B0(n50), .C0(n283), .Y(n282) );
  AOI21X1 U225 ( .A0(n200), .A1(n223), .B0(n20), .Y(n283) );
  NOR2X1 U226 ( .A(n199), .B(n4), .Y(n50) );
  NAND2X1 U227 ( .A(n284), .B(n122), .Y(n125) );
  AOI211X1 U228 ( .A0(n285), .A1(n55), .B0(n286), .C0(n287), .Y(n263) );
  AOI31X1 U229 ( .A0(n132), .A1(n288), .A2(n289), .B0(n52), .Y(n287) );
  AOI22X1 U230 ( .A0(n102), .A1(n69), .B0(n184), .B1(n33), .Y(n289) );
  NOR2X1 U231 ( .A(n290), .B(n163), .Y(n184) );
  NAND2X1 U232 ( .A(n200), .B(n284), .Y(n102) );
  INVX1 U233 ( .A(n225), .Y(n288) );
  OAI22X1 U234 ( .A0(n291), .A1(n114), .B0(n292), .B1(n10), .Y(n286) );
  INVX1 U235 ( .A(n89), .Y(n10) );
  AOI211X1 U236 ( .A0(n5), .A1(n79), .B0(n293), .C0(n294), .Y(n292) );
  AOI21X1 U237 ( .A0(n101), .A1(n150), .B0(n20), .Y(n294) );
  OAI2BB2X1 U238 ( .B0(n27), .B1(n295), .A0N(n34), .A1N(n24), .Y(n293) );
  OAI221XL U239 ( .A0(n298), .A1(n27), .B0(n20), .B1(n122), .C0(n132), .Y(n297) );
  NOR2X1 U240 ( .A(n159), .B(n217), .Y(n198) );
  NAND2X1 U241 ( .A(a[1]), .B(n47), .Y(n122) );
  NOR2X1 U242 ( .A(n299), .B(n242), .Y(n298) );
  INVX1 U243 ( .A(n99), .Y(n296) );
  NAND2X1 U244 ( .A(n200), .B(n300), .Y(n99) );
  MXI2X1 U245 ( .A(n301), .B(n147), .S0(n302), .Y(n285) );
  MXI2X1 U246 ( .A(n303), .B(n61), .S0(n69), .Y(n301) );
  INVX1 U247 ( .A(n187), .Y(n61) );
  MX2X1 U248 ( .A(n304), .B(n305), .S0(a[6]), .Y(d[1]) );
  OAI221XL U249 ( .A0(n306), .A1(n52), .B0(n307), .B1(n114), .C0(n308), .Y(
        n305) );
  AOI22X1 U250 ( .A0(n89), .A1(n309), .B0(n55), .B1(n310), .Y(n308) );
  OAI221XL U251 ( .A0(n27), .A1(n44), .B0(n4), .B1(n48), .C0(n311), .Y(n310)
         );
  AND2X1 U252 ( .A(n223), .B(n240), .Y(n28) );
  INVX1 U253 ( .A(n185), .Y(n48) );
  AOI21X1 U254 ( .A0(n226), .A1(n188), .B0(n242), .Y(n185) );
  OAI221XL U255 ( .A0(n149), .A1(n20), .B0(n4), .B1(n227), .C0(n312), .Y(n309)
         );
  AOI21X1 U256 ( .A0(n313), .A1(n33), .B0(n269), .Y(n312) );
  NAND2X1 U257 ( .A(n284), .B(n105), .Y(n227) );
  INVX1 U258 ( .A(n41), .Y(n105) );
  NOR2X1 U259 ( .A(n149), .B(n226), .Y(n41) );
  OAI22X1 U260 ( .A0(n92), .A1(n18), .B0(n316), .B1(n27), .Y(n315) );
  AOI21X1 U261 ( .A0(a[1]), .A1(n58), .B0(n98), .Y(n316) );
  INVX1 U262 ( .A(n295), .Y(n92) );
  NOR2X1 U263 ( .A(n45), .B(n163), .Y(n160) );
  INVX1 U264 ( .A(n151), .Y(n314) );
  NAND2X1 U265 ( .A(n100), .B(n199), .Y(n151) );
  AOI211X1 U266 ( .A0(n33), .A1(n120), .B0(n317), .C0(n318), .Y(n306) );
  INVX1 U267 ( .A(n258), .Y(n182) );
  OAI221XL U268 ( .A0(n20), .A1(n100), .B0(a[3]), .B1(n4), .C0(n262), .Y(n317)
         );
  INVX1 U269 ( .A(n210), .Y(n100) );
  NAND2X1 U270 ( .A(n34), .B(n200), .Y(n120) );
  INVX1 U271 ( .A(n290), .Y(n200) );
  NOR2X1 U272 ( .A(n226), .B(n58), .Y(n290) );
  OAI221XL U273 ( .A0(n319), .A1(n52), .B0(n320), .B1(n114), .C0(n321), .Y(
        n304) );
  AOI22X1 U274 ( .A0(n55), .A1(n322), .B0(n89), .B1(n323), .Y(n321) );
  OAI221XL U275 ( .A0(n47), .A1(n27), .B0(n65), .B1(n20), .C0(n324), .Y(n323)
         );
  AOI21X1 U276 ( .A0(n40), .A1(a[4]), .B0(n135), .Y(n324) );
  NOR2X1 U277 ( .A(n71), .B(n18), .Y(n135) );
  NAND2X1 U278 ( .A(n19), .B(n189), .Y(n71) );
  OAI21XL U279 ( .A0(n325), .A1(n18), .B0(n326), .Y(n322) );
  AOI31X1 U280 ( .A0(n111), .A1(n149), .A2(n327), .B0(n225), .Y(n326) );
  OAI21XL U281 ( .A0(n69), .A1(n284), .B0(n27), .Y(n327) );
  INVX1 U282 ( .A(n98), .Y(n284) );
  NOR2X1 U283 ( .A(n47), .B(a[1]), .Y(n98) );
  INVX1 U284 ( .A(n145), .Y(n149) );
  INVX1 U285 ( .A(n16), .Y(n114) );
  NOR2X1 U286 ( .A(a[0]), .B(a[5]), .Y(n16) );
  OAI32X1 U287 ( .A0(n4), .A1(n145), .A2(n210), .B0(n137), .B1(n27), .Y(n328)
         );
  AND2X1 U288 ( .A(n300), .B(n240), .Y(n23) );
  NAND2X1 U289 ( .A(n44), .B(n226), .Y(n300) );
  NOR2X1 U290 ( .A(n25), .B(n299), .Y(n313) );
  NOR2X1 U291 ( .A(n234), .B(a[5]), .Y(n14) );
  AOI221X1 U292 ( .A0(n325), .A1(n33), .B0(n24), .B1(n303), .C0(n329), .Y(n319) );
  OAI221XL U293 ( .A0(n18), .A1(n330), .B0(n20), .B1(n80), .C0(n75), .Y(n329)
         );
  INVX1 U294 ( .A(n269), .Y(n75) );
  NOR2X1 U295 ( .A(n111), .B(n18), .Y(n269) );
  INVX1 U296 ( .A(n299), .Y(n80) );
  MX4X1 U297 ( .A(n331), .B(n332), .C(n333), .D(n334), .S0(a[6]), .S1(n234), 
        .Y(d[0]) );
  NOR2X1 U298 ( .A(n258), .B(n335), .Y(n334) );
  MXI2X1 U299 ( .A(n336), .B(n337), .S0(n252), .Y(n335) );
  OAI21XL U300 ( .A0(n4), .A1(n121), .B0(n339), .Y(n338) );
  NOR2X1 U301 ( .A(n18), .B(n136), .Y(n280) );
  NAND2X1 U302 ( .A(n126), .B(n101), .Y(n178) );
  INVX1 U303 ( .A(n45), .Y(n126) );
  OAI32X1 U304 ( .A0(n27), .A1(n278), .A2(n95), .B0(n341), .B1(n4), .Y(n340)
         );
  NOR2X1 U305 ( .A(n299), .B(n210), .Y(n341) );
  NOR2X1 U306 ( .A(n136), .B(a[1]), .Y(n299) );
  NAND2X1 U307 ( .A(n204), .B(n330), .Y(n239) );
  INVX1 U308 ( .A(n179), .Y(n330) );
  NOR2X1 U309 ( .A(n188), .B(a[1]), .Y(n179) );
  NAND2X1 U310 ( .A(n278), .B(a[1]), .Y(n204) );
  NOR2X1 U311 ( .A(n18), .B(n226), .Y(n258) );
  AOI211X1 U312 ( .A0(n5), .A1(n68), .B0(n342), .C0(n343), .Y(n333) );
  AOI21X1 U313 ( .A0(n240), .A1(n37), .B0(n344), .Y(n343) );
  INVX1 U314 ( .A(n173), .Y(n344) );
  INVX1 U315 ( .A(n163), .Y(n37) );
  NOR2X1 U316 ( .A(a[1]), .B(a[3]), .Y(n163) );
  MXI2X1 U317 ( .A(n345), .B(n346), .S0(n252), .Y(n342) );
  NOR2X1 U318 ( .A(n27), .B(n210), .Y(n173) );
  NOR2X1 U319 ( .A(n226), .B(n259), .Y(n210) );
  NAND2X1 U320 ( .A(n19), .B(n199), .Y(n295) );
  NAND2X1 U321 ( .A(n199), .B(n205), .Y(n82) );
  NAND2X1 U322 ( .A(n94), .B(n226), .Y(n199) );
  INVX1 U323 ( .A(n278), .Y(n94) );
  NOR2X1 U324 ( .A(n225), .B(n40), .Y(n345) );
  NOR2X1 U325 ( .A(n20), .B(n159), .Y(n225) );
  NAND2X1 U326 ( .A(n240), .B(n189), .Y(n68) );
  INVX1 U327 ( .A(n157), .Y(n240) );
  NOR2X1 U328 ( .A(n44), .B(n226), .Y(n157) );
  MXI2X1 U329 ( .A(n347), .B(n348), .S0(n252), .Y(n332) );
  OAI211X1 U330 ( .A0(n349), .A1(n74), .B0(n350), .C0(n351), .Y(n348) );
  NAND2X1 U331 ( .A(n278), .B(n6), .Y(n74) );
  INVX1 U332 ( .A(n352), .Y(n349) );
  OAI221XL U333 ( .A0(n20), .A1(n34), .B0(n325), .B1(n4), .C0(n353), .Y(n347)
         );
  AOI31X1 U334 ( .A0(n6), .A1(n352), .A2(n259), .B0(n354), .Y(n353) );
  AOI21X1 U335 ( .A0(n19), .A1(n223), .B0(n27), .Y(n354) );
  NAND2X1 U336 ( .A(n145), .B(n226), .Y(n223) );
  INVX1 U337 ( .A(n281), .Y(n19) );
  NOR2X1 U338 ( .A(n226), .B(n136), .Y(n281) );
  XNOR2X1 U339 ( .A(a[5]), .B(n226), .Y(n352) );
  AND2X1 U340 ( .A(n101), .B(n79), .Y(n325) );
  INVX1 U341 ( .A(n59), .Y(n79) );
  MXI2X1 U342 ( .A(n355), .B(n356), .S0(n252), .Y(n331) );
  OAI221XL U343 ( .A0(n18), .A1(n121), .B0(n271), .B1(n20), .C0(n357), .Y(n356) );
  AOI22X1 U344 ( .A0(n33), .A1(n147), .B0(n24), .B1(n107), .Y(n357) );
  INVX1 U345 ( .A(n172), .Y(n107) );
  NOR2X1 U346 ( .A(n188), .B(n226), .Y(n25) );
  INVX1 U347 ( .A(n159), .Y(n188) );
  NAND2X1 U348 ( .A(a[4]), .B(n226), .Y(n101) );
  NAND2X1 U349 ( .A(n44), .B(n150), .Y(n147) );
  INVX1 U350 ( .A(n217), .Y(n150) );
  NOR2X1 U351 ( .A(n226), .B(n278), .Y(n217) );
  NOR2X1 U352 ( .A(n96), .B(n59), .Y(n271) );
  NOR2X1 U353 ( .A(n226), .B(n145), .Y(n59) );
  OAI211X1 U354 ( .A0(n65), .A1(n27), .B0(n158), .C0(n358), .Y(n355) );
  INVX1 U355 ( .A(n47), .Y(n96) );
  INVX1 U356 ( .A(n42), .Y(n121) );
  NOR2X1 U357 ( .A(n145), .B(a[1]), .Y(n42) );
  INVX1 U358 ( .A(n95), .Y(n111) );
  NOR2X1 U359 ( .A(n226), .B(n159), .Y(n95) );
  NAND2BX1 U360 ( .AN(n73), .B(n6), .Y(n158) );
  NOR2X1 U361 ( .A(n259), .B(n45), .Y(n73) );
  NOR2X1 U362 ( .A(n226), .B(n47), .Y(n45) );
  AND2X1 U363 ( .A(n189), .B(n205), .Y(n65) );
  INVX1 U364 ( .A(n242), .Y(n205) );
  NOR2X1 U365 ( .A(n226), .B(a[3]), .Y(n242) );
  NAND2X1 U366 ( .A(n47), .B(n226), .Y(n189) );
endmodule


module aes_sbox_1 ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358;

  AOI31XL U1 ( .A0(n79), .A1(n44), .A2(n2), .B0(n280), .Y(n339) );
  AOI31X1 U2 ( .A0(n44), .A1(n129), .A2(n130), .B0(n131), .Y(n128) );
  AOI221X1 U3 ( .A0(n40), .A1(n136), .B0(n33), .B1(n47), .C0(n156), .Y(n141)
         );
  OAI32X1 U4 ( .A0(n210), .A1(n145), .A2(n18), .B0(n27), .B1(n211), .Y(n209)
         );
  AOI222XL U5 ( .A0(n59), .A1(n43), .B0(n6), .B1(n221), .C0(n222), .C1(n187), 
        .Y(n218) );
  AOI221X1 U6 ( .A0(n278), .A1(n40), .B0(n185), .B1(n2), .C0(n279), .Y(n273)
         );
  AOI221X1 U7 ( .A0(n225), .A1(n226), .B0(n296), .B1(n6), .C0(n297), .Y(n291)
         );
  OAI32X1 U8 ( .A0(n18), .A1(a[1]), .A2(n159), .B0(a[4]), .B1(n182), .Y(n318)
         );
  AOI221XL U9 ( .A0(n314), .A1(n43), .B0(n160), .B1(n24), .C0(n315), .Y(n307)
         );
  AOI221X1 U10 ( .A0(n313), .A1(n5), .B0(n23), .B1(n2), .C0(n328), .Y(n320) );
  AOI31X1 U11 ( .A0(a[2]), .A1(n58), .A2(a[1]), .B0(n40), .Y(n350) );
  AOI222XL U12 ( .A0(n278), .A1(n24), .B0(n42), .B1(n33), .C0(n43), .C1(n136), 
        .Y(n351) );
  AOI221XL U13 ( .A0(n5), .A1(n96), .B0(n43), .B1(n239), .C0(n340), .Y(n336)
         );
  AOI221X1 U14 ( .A0(n40), .A1(n136), .B0(n33), .B1(n178), .C0(n338), .Y(n337)
         );
  OR2X2 U15 ( .A(a[2]), .B(a[7]), .Y(n1) );
  AOI221X1 U16 ( .A0(n5), .A1(n19), .B0(n33), .B1(n34), .C0(n35), .Y(n11) );
  OAI222X1 U17 ( .A0(n4), .A1(n37), .B0(n38), .B1(n20), .C0(a[4]), .C1(n39), 
        .Y(n35) );
  OAI222X1 U18 ( .A0(n20), .A1(n99), .B0(n27), .B1(n101), .C0(n184), .C1(n4), 
        .Y(n250) );
  OAI222X1 U19 ( .A0(n27), .A1(n34), .B0(n69), .B1(n205), .C0(n20), .C1(n79), 
        .Y(n260) );
  NAND2X2 U20 ( .A(n58), .B(n226), .Y(n34) );
  NOR2BXL U21 ( .AN(n101), .B(n25), .Y(n172) );
  AOI221XL U22 ( .A0(n43), .A1(n151), .B0(n25), .B1(n69), .C0(n275), .Y(n274)
         );
  NAND2XL U23 ( .A(n111), .B(n121), .Y(n303) );
  NAND2XL U24 ( .A(n111), .B(n300), .Y(n187) );
  NAND2XL U25 ( .A(n111), .B(n101), .Y(n21) );
  OAI2BB2XL U26 ( .B0(n20), .B1(n111), .A0N(n125), .A1N(n24), .Y(n220) );
  NAND2XL U27 ( .A(n198), .B(n24), .Y(n132) );
  AOI22XL U28 ( .A0(n33), .A1(a[3]), .B0(n24), .B1(n58), .Y(n277) );
  AOI22XL U29 ( .A0(n23), .A1(n24), .B0(n25), .B1(a[2]), .Y(n22) );
  AOI21XL U30 ( .A0(n44), .A1(n111), .B0(n4), .Y(n177) );
  NOR2X2 U31 ( .A(n44), .B(a[1]), .Y(n137) );
  CLKINVX3 U32 ( .A(n259), .Y(n44) );
  NOR2X2 U33 ( .A(n259), .B(n278), .Y(n47) );
  NOR2X2 U34 ( .A(a[4]), .B(a[3]), .Y(n278) );
  NOR2X2 U35 ( .A(n136), .B(n58), .Y(n259) );
  NOR2X2 U36 ( .A(n58), .B(a[3]), .Y(n159) );
  CLKINVX3 U37 ( .A(a[4]), .Y(n58) );
  NOR2X2 U38 ( .A(n136), .B(a[4]), .Y(n145) );
  CLKINVX3 U39 ( .A(a[3]), .Y(n136) );
  NOR2X4 U40 ( .A(n226), .B(n4), .Y(n40) );
  INVX4 U41 ( .A(a[2]), .Y(n69) );
  AOI21XL U42 ( .A0(n18), .A1(n162), .B0(n25), .Y(n161) );
  INVX4 U43 ( .A(n6), .Y(n18) );
  INVXL U44 ( .A(n20), .Y(n2) );
  MXI2XL U45 ( .A(n2), .B(n6), .S0(n28), .Y(n311) );
  NOR2XL U46 ( .A(n33), .B(n2), .Y(n302) );
  AOI22XL U47 ( .A0(n184), .A1(n5), .B0(n198), .B1(n43), .Y(n197) );
  AOI22XL U48 ( .A0(n40), .A1(n94), .B0(n43), .B1(n187), .Y(n244) );
  AOI21XL U49 ( .A0(n159), .A1(n43), .B0(n40), .Y(n262) );
  AOI22XL U50 ( .A0(n43), .A1(n100), .B0(n24), .B1(n125), .Y(n124) );
  AOI22XL U51 ( .A0(n43), .A1(n303), .B0(n24), .B1(n96), .Y(n358) );
  AOI222X4 U52 ( .A0(n125), .A1(n33), .B0(n145), .B1(n40), .C0(n43), .C1(n184), 
        .Y(n183) );
  AOI2BB2XL U53 ( .B0(n43), .B1(n94), .A0N(n120), .A1N(n4), .Y(n119) );
  AOI22XL U54 ( .A0(n82), .A1(n43), .B0(n83), .B1(n24), .Y(n81) );
  AOI22XL U55 ( .A0(n98), .A1(n43), .B0(n6), .B1(n99), .Y(n97) );
  AOI22XL U56 ( .A0(n217), .A1(n43), .B0(n33), .B1(n47), .Y(n216) );
  AOI221X4 U57 ( .A0(n43), .A1(n44), .B0(n45), .B1(n24), .C0(n46), .Y(n9) );
  AOI221X4 U58 ( .A0(n43), .A1(n205), .B0(n32), .B1(n6), .C0(n206), .Y(n201)
         );
  AOI221X4 U59 ( .A0(n43), .A1(n208), .B0(n76), .B1(n24), .C0(n209), .Y(n207)
         );
  AOI221X4 U60 ( .A0(n70), .A1(n43), .B0(n24), .B1(n71), .C0(n72), .Y(n53) );
  AOI222X4 U61 ( .A0(n185), .A1(n43), .B0(n186), .B1(n187), .C0(n6), .C1(n188), 
        .Y(n164) );
  AOI222X4 U62 ( .A0(n123), .A1(n43), .B0(a[2]), .B1(n203), .C0(n6), .C1(n71), 
        .Y(n202) );
  AOI221X4 U63 ( .A0(n59), .A1(n33), .B0(n43), .B1(n126), .C0(n127), .Y(n113)
         );
  AOI221X4 U64 ( .A0(n24), .A1(n82), .B0(n43), .B1(n295), .C0(n173), .Y(n346)
         );
  INVX4 U65 ( .A(n43), .Y(n20) );
  INVXL U66 ( .A(n36), .Y(n3) );
  INVX4 U67 ( .A(n3), .Y(n4) );
  INVXL U68 ( .A(n24), .Y(n36) );
  CLKINVX3 U69 ( .A(n1), .Y(n5) );
  CLKINVX3 U70 ( .A(n1), .Y(n6) );
  INVX12 U71 ( .A(n33), .Y(n27) );
  NOR2X4 U72 ( .A(n69), .B(a[7]), .Y(n33) );
  CLKINVX3 U73 ( .A(a[0]), .Y(n234) );
  NOR2X2 U74 ( .A(n252), .B(a[0]), .Y(n89) );
  AOI22XL U75 ( .A0(n70), .A1(n24), .B0(n96), .B1(n129), .Y(n241) );
  NOR2X4 U76 ( .A(n129), .B(n69), .Y(n24) );
  CLKINVX3 U77 ( .A(a[7]), .Y(n129) );
  NOR2X2 U78 ( .A(n252), .B(n234), .Y(n55) );
  CLKINVX3 U79 ( .A(a[5]), .Y(n252) );
  AOI22XL U80 ( .A0(n225), .A1(n226), .B0(n6), .B1(n227), .Y(n224) );
  INVX4 U81 ( .A(a[1]), .Y(n226) );
  OAI22XL U82 ( .A0(n201), .A1(n52), .B0(n202), .B1(n114), .Y(n193) );
  CLKINVX3 U83 ( .A(n14), .Y(n52) );
  NOR2X4 U84 ( .A(n129), .B(a[2]), .Y(n43) );
  MX2X1 U85 ( .A(n7), .B(n8), .S0(a[6]), .Y(d[7]) );
  OAI221XL U86 ( .A0(n9), .A1(n10), .B0(n11), .B1(n12), .C0(n13), .Y(n8) );
  AOI22X1 U87 ( .A0(n14), .A1(n15), .B0(n16), .B1(n17), .Y(n13) );
  OAI221XL U88 ( .A0(n18), .A1(n19), .B0(n20), .B1(n21), .C0(n22), .Y(n17) );
  OAI221XL U89 ( .A0(n26), .A1(n27), .B0(n28), .B1(n20), .C0(n29), .Y(n15) );
  AOI21X1 U90 ( .A0(n5), .A1(n30), .B0(n31), .Y(n29) );
  INVX1 U91 ( .A(n32), .Y(n26) );
  INVX1 U92 ( .A(n40), .Y(n39) );
  NOR2X1 U93 ( .A(n41), .B(n42), .Y(n38) );
  OAI221XL U94 ( .A0(n47), .A1(n18), .B0(n27), .B1(n48), .C0(n49), .Y(n46) );
  INVX1 U95 ( .A(n50), .Y(n49) );
  OAI221XL U96 ( .A0(n51), .A1(n52), .B0(n53), .B1(n10), .C0(n54), .Y(n7) );
  AOI22X1 U97 ( .A0(n55), .A1(n56), .B0(n16), .B1(n57), .Y(n54) );
  OAI221XL U98 ( .A0(n58), .A1(n18), .B0(n59), .B1(n27), .C0(n60), .Y(n57) );
  AOI2BB2X1 U99 ( .B0(n61), .B1(n24), .A0N(n62), .A1N(n20), .Y(n60) );
  OAI221XL U100 ( .A0(n63), .A1(n64), .B0(n65), .B1(n27), .C0(n66), .Y(n56) );
  INVX1 U101 ( .A(n67), .Y(n66) );
  AOI21X1 U102 ( .A0(n68), .A1(n69), .B0(n6), .Y(n63) );
  OAI211X1 U103 ( .A0(n73), .A1(n27), .B0(n74), .C0(n75), .Y(n72) );
  AOI211X1 U104 ( .A0(n5), .A1(n76), .B0(n77), .C0(n78), .Y(n51) );
  AOI21X1 U105 ( .A0(n79), .A1(n80), .B0(n27), .Y(n78) );
  INVX1 U106 ( .A(n81), .Y(n77) );
  MX2X1 U107 ( .A(n84), .B(n85), .S0(a[6]), .Y(d[6]) );
  OAI221XL U108 ( .A0(n86), .A1(n52), .B0(n87), .B1(n12), .C0(n88), .Y(n85) );
  AOI22X1 U109 ( .A0(n89), .A1(n90), .B0(n16), .B1(n91), .Y(n88) );
  OAI221XL U110 ( .A0(n73), .A1(n27), .B0(n92), .B1(n20), .C0(n93), .Y(n91) );
  AOI31X1 U111 ( .A0(n79), .A1(n94), .A2(n6), .B0(n67), .Y(n93) );
  NOR3X1 U112 ( .A(n4), .B(n95), .C(n96), .Y(n67) );
  OAI221XL U113 ( .A0(n27), .A1(n62), .B0(n4), .B1(n21), .C0(n97), .Y(n90) );
  NAND2X1 U114 ( .A(n100), .B(n101), .Y(n62) );
  AOI211X1 U115 ( .A0(n33), .A1(n102), .B0(n103), .C0(n104), .Y(n87) );
  AOI21X1 U116 ( .A0(n105), .A1(n106), .B0(n20), .Y(n104) );
  OAI22X1 U117 ( .A0(n45), .A1(n4), .B0(a[4]), .B1(n18), .Y(n103) );
  AOI211X1 U118 ( .A0(n5), .A1(n107), .B0(n108), .C0(n109), .Y(n86) );
  AOI21X1 U119 ( .A0(a[1]), .A1(n58), .B0(n27), .Y(n109) );
  OAI22X1 U120 ( .A0(n110), .A1(n4), .B0(n20), .B1(n21), .Y(n108) );
  OAI221XL U121 ( .A0(n112), .A1(n52), .B0(n113), .B1(n114), .C0(n115), .Y(n84) );
  AOI22X1 U122 ( .A0(n89), .A1(n116), .B0(n55), .B1(n117), .Y(n115) );
  OAI221XL U123 ( .A0(n18), .A1(n118), .B0(n27), .B1(n30), .C0(n119), .Y(n117)
         );
  NAND2X1 U124 ( .A(n121), .B(n122), .Y(n30) );
  OAI221XL U125 ( .A0(n18), .A1(n105), .B0(n123), .B1(n27), .C0(n124), .Y(n116) );
  OAI21XL U126 ( .A0(n18), .A1(n37), .B0(n128), .Y(n127) );
  INVX1 U127 ( .A(n132), .Y(n131) );
  AOI211X1 U128 ( .A0(n133), .A1(n69), .B0(n134), .C0(n135), .Y(n112) );
  OAI22X1 U129 ( .A0(n4), .A1(n136), .B0(n137), .B1(n27), .Y(n134) );
  INVX1 U130 ( .A(n70), .Y(n133) );
  MX2X1 U131 ( .A(n138), .B(n139), .S0(a[6]), .Y(d[5]) );
  OAI221XL U132 ( .A0(n140), .A1(n12), .B0(n141), .B1(n114), .C0(n142), .Y(
        n139) );
  AOI22X1 U133 ( .A0(n89), .A1(n143), .B0(n14), .B1(n144), .Y(n142) );
  OAI221XL U134 ( .A0(n145), .A1(n20), .B0(n4), .B1(n34), .C0(n146), .Y(n144)
         );
  AOI2BB1X1 U135 ( .A0N(n147), .A1N(n27), .B0(n148), .Y(n146) );
  AOI21X1 U136 ( .A0(n149), .A1(n150), .B0(n18), .Y(n148) );
  OAI221XL U137 ( .A0(n110), .A1(n18), .B0(n20), .B1(n151), .C0(n152), .Y(n143) );
  MXI2X1 U138 ( .A(n153), .B(n154), .S0(n155), .Y(n152) );
  NOR2X1 U139 ( .A(n145), .B(n69), .Y(n154) );
  NOR2X1 U140 ( .A(n4), .B(n136), .Y(n153) );
  OAI21XL U141 ( .A0(n157), .A1(n20), .B0(n158), .Y(n156) );
  AOI221X1 U142 ( .A0(n159), .A1(n24), .B0(n160), .B1(n33), .C0(n161), .Y(n140) );
  OAI21XL U143 ( .A0(n41), .A1(n163), .B0(n69), .Y(n162) );
  OAI221XL U144 ( .A0(n164), .A1(n114), .B0(n165), .B1(n52), .C0(n166), .Y(
        n138) );
  AOI22X1 U145 ( .A0(n89), .A1(n167), .B0(n55), .B1(n168), .Y(n166) );
  OAI211X1 U146 ( .A0(n20), .A1(n169), .B0(n170), .C0(n171), .Y(n168) );
  AOI22X1 U147 ( .A0(n137), .A1(n24), .B0(n172), .B1(n6), .Y(n171) );
  MXI2X1 U148 ( .A(n40), .B(n173), .S0(n96), .Y(n170) );
  OAI221XL U149 ( .A0(n159), .A1(n27), .B0(n145), .B1(n20), .C0(n174), .Y(n167) );
  AOI211X1 U150 ( .A0(n175), .A1(n5), .B0(n176), .C0(n177), .Y(n174) );
  INVX1 U151 ( .A(n178), .Y(n175) );
  AOI211X1 U152 ( .A0(n179), .A1(n24), .B0(n180), .C0(n181), .Y(n165) );
  NAND2X1 U153 ( .A(n74), .B(n182), .Y(n181) );
  INVX1 U154 ( .A(n183), .Y(n180) );
  OAI21XL U155 ( .A0(n69), .A1(n189), .B0(n27), .Y(n186) );
  MXI2X1 U156 ( .A(n190), .B(n191), .S0(a[6]), .Y(d[4]) );
  AOI211X1 U157 ( .A0(n89), .A1(n192), .B0(n193), .C0(n194), .Y(n191) );
  AOI31X1 U158 ( .A0(n195), .A1(n196), .A2(n197), .B0(n12), .Y(n194) );
  INVX1 U159 ( .A(n55), .Y(n12) );
  OAI2BB1X1 U160 ( .A0N(n199), .A1N(n200), .B0(n33), .Y(n195) );
  NAND2X1 U161 ( .A(n94), .B(n79), .Y(n203) );
  INVX1 U162 ( .A(n118), .Y(n123) );
  NAND2X1 U163 ( .A(n204), .B(n80), .Y(n118) );
  OAI22X1 U164 ( .A0(n28), .A1(n4), .B0(n188), .B1(n27), .Y(n206) );
  NOR2X1 U165 ( .A(n25), .B(n98), .Y(n32) );
  INVX1 U166 ( .A(n207), .Y(n192) );
  AOI211X1 U167 ( .A0(n55), .A1(n212), .B0(n213), .C0(n214), .Y(n190) );
  AOI31X1 U168 ( .A0(n215), .A1(n196), .A2(n216), .B0(n52), .Y(n214) );
  INVX1 U169 ( .A(n31), .Y(n196) );
  NOR2X1 U170 ( .A(n4), .B(n159), .Y(n31) );
  INVX1 U171 ( .A(n135), .Y(n215) );
  OAI22X1 U172 ( .A0(n218), .A1(n10), .B0(n219), .B1(n114), .Y(n213) );
  AOI211X1 U173 ( .A0(n208), .A1(n5), .B0(n220), .C0(n173), .Y(n219) );
  NOR2X1 U174 ( .A(n217), .B(n42), .Y(n208) );
  OAI21XL U175 ( .A0(n69), .A1(n223), .B0(n27), .Y(n222) );
  NAND2X1 U176 ( .A(n34), .B(n204), .Y(n221) );
  OAI221XL U177 ( .A0(n27), .A1(n64), .B0(n4), .B1(n83), .C0(n224), .Y(n212)
         );
  INVX1 U178 ( .A(n110), .Y(n64) );
  NOR2BX1 U179 ( .AN(n204), .B(n137), .Y(n110) );
  MX2X1 U180 ( .A(n228), .B(n229), .S0(a[6]), .Y(d[3]) );
  MX4X1 U181 ( .A(n230), .B(n231), .C(n232), .D(n233), .S0(n234), .S1(a[5]), 
        .Y(n229) );
  OAI211X1 U182 ( .A0(n27), .A1(n122), .B0(n158), .C0(n235), .Y(n233) );
  AOI2BB2X1 U183 ( .B0(n24), .B1(n187), .A0N(n227), .A1N(n20), .Y(n235) );
  OAI221XL U184 ( .A0(n18), .A1(n76), .B0(n59), .B1(n27), .C0(n236), .Y(n232)
         );
  OAI21XL U185 ( .A0(n237), .A1(n43), .B0(n238), .Y(n236) );
  INVX1 U186 ( .A(n239), .Y(n238) );
  AOI21X1 U187 ( .A0(n122), .A1(n106), .B0(n129), .Y(n237) );
  NAND2X1 U188 ( .A(n101), .B(n240), .Y(n76) );
  OAI221XL U189 ( .A0(n159), .A1(n27), .B0(n20), .B1(n34), .C0(n241), .Y(n231)
         );
  NOR2X1 U190 ( .A(n242), .B(n137), .Y(n70) );
  OAI211X1 U191 ( .A0(n4), .A1(n149), .B0(n243), .C0(n244), .Y(n230) );
  MXI2X1 U192 ( .A(n245), .B(n246), .S0(n130), .Y(n243) );
  XNOR2X1 U193 ( .A(n69), .B(a[1]), .Y(n130) );
  NOR2X1 U194 ( .A(a[7]), .B(n145), .Y(n246) );
  OAI21XL U195 ( .A0(n58), .A1(n27), .B0(n247), .Y(n245) );
  MXI2X1 U196 ( .A(n248), .B(n249), .S0(n234), .Y(n228) );
  MXI2X1 U197 ( .A(n250), .B(n251), .S0(n252), .Y(n249) );
  OAI221XL U198 ( .A0(n172), .A1(n18), .B0(n27), .B1(n83), .C0(n253), .Y(n251)
         );
  AOI2BB2X1 U199 ( .B0(n65), .B1(n24), .A0N(n169), .A1N(n20), .Y(n253) );
  NAND2X1 U200 ( .A(n199), .B(n204), .Y(n169) );
  NAND2X1 U201 ( .A(n200), .B(n106), .Y(n83) );
  INVX1 U202 ( .A(n211), .Y(n106) );
  AOI221X1 U203 ( .A0(n211), .A1(n5), .B0(n40), .B1(a[4]), .C0(n254), .Y(n248)
         );
  MXI2X1 U204 ( .A(n255), .B(n256), .S0(n252), .Y(n254) );
  NOR3X1 U205 ( .A(n257), .B(n258), .C(n50), .Y(n256) );
  OAI22X1 U206 ( .A0(n20), .A1(n68), .B0(n27), .B1(n37), .Y(n257) );
  AOI211X1 U207 ( .A0(n259), .A1(n24), .B0(n260), .C0(n261), .Y(n255) );
  INVX1 U208 ( .A(n262), .Y(n261) );
  NOR2X1 U209 ( .A(n94), .B(a[1]), .Y(n211) );
  MXI2X1 U210 ( .A(n263), .B(n264), .S0(a[6]), .Y(d[2]) );
  AOI211X1 U211 ( .A0(n55), .A1(n265), .B0(n266), .C0(n267), .Y(n264) );
  INVX1 U212 ( .A(n268), .Y(n267) );
  OAI31X1 U213 ( .A0(n176), .A1(n269), .A2(n270), .B0(n16), .Y(n268) );
  OAI21XL U214 ( .A0(n4), .A1(n271), .B0(n272), .Y(n270) );
  NOR2X1 U215 ( .A(n20), .B(n226), .Y(n176) );
  OAI22X1 U216 ( .A0(n273), .A1(n10), .B0(n274), .B1(n52), .Y(n266) );
  MXI2X1 U217 ( .A(n276), .B(n277), .S0(n155), .Y(n275) );
  XNOR2X1 U218 ( .A(n129), .B(a[1]), .Y(n155) );
  NAND2X1 U219 ( .A(a[2]), .B(n149), .Y(n276) );
  OAI221XL U220 ( .A0(a[1]), .A1(n247), .B0(n4), .B1(n189), .C0(n272), .Y(n279) );
  NAND2X1 U221 ( .A(n41), .B(n33), .Y(n272) );
  INVX1 U222 ( .A(n280), .Y(n247) );
  OAI221XL U223 ( .A0(n281), .A1(n27), .B0(n4), .B1(n111), .C0(n282), .Y(n265)
         );
  AOI211X1 U224 ( .A0(n5), .A1(n125), .B0(n50), .C0(n283), .Y(n282) );
  AOI21X1 U225 ( .A0(n200), .A1(n223), .B0(n20), .Y(n283) );
  NOR2X1 U226 ( .A(n199), .B(n4), .Y(n50) );
  NAND2X1 U227 ( .A(n284), .B(n122), .Y(n125) );
  AOI211X1 U228 ( .A0(n285), .A1(n55), .B0(n286), .C0(n287), .Y(n263) );
  AOI31X1 U229 ( .A0(n132), .A1(n288), .A2(n289), .B0(n52), .Y(n287) );
  AOI22X1 U230 ( .A0(n102), .A1(n69), .B0(n184), .B1(n33), .Y(n289) );
  NOR2X1 U231 ( .A(n290), .B(n163), .Y(n184) );
  NAND2X1 U232 ( .A(n200), .B(n284), .Y(n102) );
  INVX1 U233 ( .A(n225), .Y(n288) );
  OAI22X1 U234 ( .A0(n291), .A1(n114), .B0(n292), .B1(n10), .Y(n286) );
  INVX1 U235 ( .A(n89), .Y(n10) );
  AOI211X1 U236 ( .A0(n5), .A1(n79), .B0(n293), .C0(n294), .Y(n292) );
  AOI21X1 U237 ( .A0(n101), .A1(n150), .B0(n20), .Y(n294) );
  OAI2BB2X1 U238 ( .B0(n27), .B1(n295), .A0N(n34), .A1N(n24), .Y(n293) );
  OAI221XL U239 ( .A0(n298), .A1(n27), .B0(n20), .B1(n122), .C0(n132), .Y(n297) );
  NOR2X1 U240 ( .A(n159), .B(n217), .Y(n198) );
  NAND2X1 U241 ( .A(a[1]), .B(n47), .Y(n122) );
  NOR2X1 U242 ( .A(n299), .B(n242), .Y(n298) );
  INVX1 U243 ( .A(n99), .Y(n296) );
  NAND2X1 U244 ( .A(n200), .B(n300), .Y(n99) );
  MXI2X1 U245 ( .A(n301), .B(n147), .S0(n302), .Y(n285) );
  MXI2X1 U246 ( .A(n303), .B(n61), .S0(n69), .Y(n301) );
  INVX1 U247 ( .A(n187), .Y(n61) );
  MX2X1 U248 ( .A(n304), .B(n305), .S0(a[6]), .Y(d[1]) );
  OAI221XL U249 ( .A0(n306), .A1(n52), .B0(n307), .B1(n114), .C0(n308), .Y(
        n305) );
  AOI22X1 U250 ( .A0(n89), .A1(n309), .B0(n55), .B1(n310), .Y(n308) );
  OAI221XL U251 ( .A0(n27), .A1(n44), .B0(n4), .B1(n48), .C0(n311), .Y(n310)
         );
  AND2X1 U252 ( .A(n223), .B(n240), .Y(n28) );
  INVX1 U253 ( .A(n185), .Y(n48) );
  AOI21X1 U254 ( .A0(n226), .A1(n188), .B0(n242), .Y(n185) );
  OAI221XL U255 ( .A0(n149), .A1(n20), .B0(n4), .B1(n227), .C0(n312), .Y(n309)
         );
  AOI21X1 U256 ( .A0(n313), .A1(n33), .B0(n269), .Y(n312) );
  NAND2X1 U257 ( .A(n284), .B(n105), .Y(n227) );
  INVX1 U258 ( .A(n41), .Y(n105) );
  NOR2X1 U259 ( .A(n149), .B(n226), .Y(n41) );
  OAI22X1 U260 ( .A0(n92), .A1(n18), .B0(n316), .B1(n27), .Y(n315) );
  AOI21X1 U261 ( .A0(a[1]), .A1(n58), .B0(n98), .Y(n316) );
  INVX1 U262 ( .A(n295), .Y(n92) );
  NOR2X1 U263 ( .A(n45), .B(n163), .Y(n160) );
  INVX1 U264 ( .A(n151), .Y(n314) );
  NAND2X1 U265 ( .A(n100), .B(n199), .Y(n151) );
  AOI211X1 U266 ( .A0(n33), .A1(n120), .B0(n317), .C0(n318), .Y(n306) );
  INVX1 U267 ( .A(n258), .Y(n182) );
  OAI221XL U268 ( .A0(n20), .A1(n100), .B0(a[3]), .B1(n4), .C0(n262), .Y(n317)
         );
  INVX1 U269 ( .A(n210), .Y(n100) );
  NAND2X1 U270 ( .A(n34), .B(n200), .Y(n120) );
  INVX1 U271 ( .A(n290), .Y(n200) );
  NOR2X1 U272 ( .A(n226), .B(n58), .Y(n290) );
  OAI221XL U273 ( .A0(n319), .A1(n52), .B0(n320), .B1(n114), .C0(n321), .Y(
        n304) );
  AOI22X1 U274 ( .A0(n55), .A1(n322), .B0(n89), .B1(n323), .Y(n321) );
  OAI221XL U275 ( .A0(n47), .A1(n27), .B0(n65), .B1(n20), .C0(n324), .Y(n323)
         );
  AOI21X1 U276 ( .A0(n40), .A1(a[4]), .B0(n135), .Y(n324) );
  NOR2X1 U277 ( .A(n71), .B(n18), .Y(n135) );
  NAND2X1 U278 ( .A(n19), .B(n189), .Y(n71) );
  OAI21XL U279 ( .A0(n325), .A1(n18), .B0(n326), .Y(n322) );
  AOI31X1 U280 ( .A0(n111), .A1(n149), .A2(n327), .B0(n225), .Y(n326) );
  OAI21XL U281 ( .A0(n69), .A1(n284), .B0(n27), .Y(n327) );
  INVX1 U282 ( .A(n98), .Y(n284) );
  NOR2X1 U283 ( .A(n47), .B(a[1]), .Y(n98) );
  INVX1 U284 ( .A(n145), .Y(n149) );
  INVX1 U285 ( .A(n16), .Y(n114) );
  NOR2X1 U286 ( .A(a[0]), .B(a[5]), .Y(n16) );
  OAI32X1 U287 ( .A0(n4), .A1(n145), .A2(n210), .B0(n137), .B1(n27), .Y(n328)
         );
  AND2X1 U288 ( .A(n300), .B(n240), .Y(n23) );
  NAND2X1 U289 ( .A(n44), .B(n226), .Y(n300) );
  NOR2X1 U290 ( .A(n25), .B(n299), .Y(n313) );
  NOR2X1 U291 ( .A(n234), .B(a[5]), .Y(n14) );
  AOI221X1 U292 ( .A0(n325), .A1(n33), .B0(n24), .B1(n303), .C0(n329), .Y(n319) );
  OAI221XL U293 ( .A0(n18), .A1(n330), .B0(n20), .B1(n80), .C0(n75), .Y(n329)
         );
  INVX1 U294 ( .A(n269), .Y(n75) );
  NOR2X1 U295 ( .A(n111), .B(n18), .Y(n269) );
  INVX1 U296 ( .A(n299), .Y(n80) );
  MX4X1 U297 ( .A(n331), .B(n332), .C(n333), .D(n334), .S0(a[6]), .S1(n234), 
        .Y(d[0]) );
  NOR2X1 U298 ( .A(n258), .B(n335), .Y(n334) );
  MXI2X1 U299 ( .A(n336), .B(n337), .S0(n252), .Y(n335) );
  OAI21XL U300 ( .A0(n4), .A1(n121), .B0(n339), .Y(n338) );
  NOR2X1 U301 ( .A(n18), .B(n136), .Y(n280) );
  NAND2X1 U302 ( .A(n126), .B(n101), .Y(n178) );
  INVX1 U303 ( .A(n45), .Y(n126) );
  OAI32X1 U304 ( .A0(n27), .A1(n278), .A2(n95), .B0(n341), .B1(n4), .Y(n340)
         );
  NOR2X1 U305 ( .A(n299), .B(n210), .Y(n341) );
  NOR2X1 U306 ( .A(n136), .B(a[1]), .Y(n299) );
  NAND2X1 U307 ( .A(n204), .B(n330), .Y(n239) );
  INVX1 U308 ( .A(n179), .Y(n330) );
  NOR2X1 U309 ( .A(n188), .B(a[1]), .Y(n179) );
  NAND2X1 U310 ( .A(n278), .B(a[1]), .Y(n204) );
  NOR2X1 U311 ( .A(n18), .B(n226), .Y(n258) );
  AOI211X1 U312 ( .A0(n5), .A1(n68), .B0(n342), .C0(n343), .Y(n333) );
  AOI21X1 U313 ( .A0(n240), .A1(n37), .B0(n344), .Y(n343) );
  INVX1 U314 ( .A(n173), .Y(n344) );
  INVX1 U315 ( .A(n163), .Y(n37) );
  NOR2X1 U316 ( .A(a[1]), .B(a[3]), .Y(n163) );
  MXI2X1 U317 ( .A(n345), .B(n346), .S0(n252), .Y(n342) );
  NOR2X1 U318 ( .A(n27), .B(n210), .Y(n173) );
  NOR2X1 U319 ( .A(n226), .B(n259), .Y(n210) );
  NAND2X1 U320 ( .A(n19), .B(n199), .Y(n295) );
  NAND2X1 U321 ( .A(n199), .B(n205), .Y(n82) );
  NAND2X1 U322 ( .A(n94), .B(n226), .Y(n199) );
  INVX1 U323 ( .A(n278), .Y(n94) );
  NOR2X1 U324 ( .A(n225), .B(n40), .Y(n345) );
  NOR2X1 U325 ( .A(n20), .B(n159), .Y(n225) );
  NAND2X1 U326 ( .A(n240), .B(n189), .Y(n68) );
  INVX1 U327 ( .A(n157), .Y(n240) );
  NOR2X1 U328 ( .A(n44), .B(n226), .Y(n157) );
  MXI2X1 U329 ( .A(n347), .B(n348), .S0(n252), .Y(n332) );
  OAI211X1 U330 ( .A0(n349), .A1(n74), .B0(n350), .C0(n351), .Y(n348) );
  NAND2X1 U331 ( .A(n278), .B(n6), .Y(n74) );
  INVX1 U332 ( .A(n352), .Y(n349) );
  OAI221XL U333 ( .A0(n20), .A1(n34), .B0(n325), .B1(n4), .C0(n353), .Y(n347)
         );
  AOI31X1 U334 ( .A0(n6), .A1(n352), .A2(n259), .B0(n354), .Y(n353) );
  AOI21X1 U335 ( .A0(n19), .A1(n223), .B0(n27), .Y(n354) );
  NAND2X1 U336 ( .A(n145), .B(n226), .Y(n223) );
  INVX1 U337 ( .A(n281), .Y(n19) );
  NOR2X1 U338 ( .A(n226), .B(n136), .Y(n281) );
  XNOR2X1 U339 ( .A(a[5]), .B(n226), .Y(n352) );
  AND2X1 U340 ( .A(n101), .B(n79), .Y(n325) );
  INVX1 U341 ( .A(n59), .Y(n79) );
  MXI2X1 U342 ( .A(n355), .B(n356), .S0(n252), .Y(n331) );
  OAI221XL U343 ( .A0(n18), .A1(n121), .B0(n271), .B1(n20), .C0(n357), .Y(n356) );
  AOI22X1 U344 ( .A0(n33), .A1(n147), .B0(n24), .B1(n107), .Y(n357) );
  INVX1 U345 ( .A(n172), .Y(n107) );
  NOR2X1 U346 ( .A(n188), .B(n226), .Y(n25) );
  INVX1 U347 ( .A(n159), .Y(n188) );
  NAND2X1 U348 ( .A(a[4]), .B(n226), .Y(n101) );
  NAND2X1 U349 ( .A(n44), .B(n150), .Y(n147) );
  INVX1 U350 ( .A(n217), .Y(n150) );
  NOR2X1 U351 ( .A(n226), .B(n278), .Y(n217) );
  NOR2X1 U352 ( .A(n96), .B(n59), .Y(n271) );
  NOR2X1 U353 ( .A(n226), .B(n145), .Y(n59) );
  OAI211X1 U354 ( .A0(n65), .A1(n27), .B0(n158), .C0(n358), .Y(n355) );
  INVX1 U355 ( .A(n47), .Y(n96) );
  INVX1 U356 ( .A(n42), .Y(n121) );
  NOR2X1 U357 ( .A(n145), .B(a[1]), .Y(n42) );
  INVX1 U358 ( .A(n95), .Y(n111) );
  NOR2X1 U359 ( .A(n226), .B(n159), .Y(n95) );
  NAND2BX1 U360 ( .AN(n73), .B(n6), .Y(n158) );
  NOR2X1 U361 ( .A(n259), .B(n45), .Y(n73) );
  NOR2X1 U362 ( .A(n226), .B(n47), .Y(n45) );
  AND2X1 U363 ( .A(n189), .B(n205), .Y(n65) );
  INVX1 U364 ( .A(n242), .Y(n205) );
  NOR2X1 U365 ( .A(n226), .B(a[3]), .Y(n242) );
  NAND2X1 U366 ( .A(n47), .B(n226), .Y(n189) );
endmodule


module aes_rcon ( clk, kld, out );
  output [31:0] out;
  input clk, kld;
  wire   N44, N45, N46, N47, N48, N49, N51, N55, n1, n2, n9, n14, n4, n5, n6,
         n7, n8, n10, n11, n12, n13, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27;
  wire   [3:0] rcnt;
  assign out[23] = 1'b0;
  assign out[22] = 1'b0;
  assign out[21] = 1'b0;
  assign out[20] = 1'b0;
  assign out[19] = 1'b0;
  assign out[18] = 1'b0;
  assign out[17] = 1'b0;
  assign out[16] = 1'b0;
  assign out[15] = 1'b0;
  assign out[14] = 1'b0;
  assign out[13] = 1'b0;
  assign out[12] = 1'b0;
  assign out[11] = 1'b0;
  assign out[10] = 1'b0;
  assign out[9] = 1'b0;
  assign out[8] = 1'b0;
  assign out[7] = 1'b0;
  assign out[6] = 1'b0;
  assign out[5] = 1'b0;
  assign out[4] = 1'b0;
  assign out[3] = 1'b0;
  assign out[2] = 1'b0;
  assign out[1] = 1'b0;
  assign out[0] = 1'b0;

  DFFX1 \rcnt_reg[3]  ( .D(N55), .CK(clk), .Q(n27), .QN(n6) );
  DFFTRX1 \rcnt_reg[2]  ( .D(n2), .RN(n9), .CK(clk), .Q(rcnt[2]), .QN(n5) );
  DFFTRX1 \rcnt_reg[1]  ( .D(n14), .RN(n9), .CK(clk), .Q(rcnt[1]) );
  DFFTRX1 \out_reg[30]  ( .D(n14), .RN(n1), .CK(clk), .Q(out[30]) );
  DFFHQX1 \out_reg[24]  ( .D(N44), .CK(clk), .Q(out[24]) );
  DFFHQX1 \out_reg[31]  ( .D(N51), .CK(clk), .Q(out[31]) );
  DFFHQX1 \out_reg[27]  ( .D(N47), .CK(clk), .Q(out[27]) );
  DFFHQX1 \out_reg[26]  ( .D(N46), .CK(clk), .Q(out[26]) );
  DFFHQX1 \out_reg[25]  ( .D(N45), .CK(clk), .Q(out[25]) );
  DFFHQX1 \out_reg[29]  ( .D(N49), .CK(clk), .Q(out[29]) );
  DFFHQX1 \out_reg[28]  ( .D(N48), .CK(clk), .Q(out[28]) );
  JKFFX1 \rcnt_reg[0]  ( .J(n9), .K(1'b1), .CK(clk), .Q(rcnt[0]), .QN(n4) );
  INVX1 U3 ( .A(n7), .Y(n1) );
  OAI21XL U4 ( .A0(N44), .A1(n6), .B0(n8), .Y(N55) );
  NOR3X1 U30 ( .A(n10), .B(kld), .C(n11), .Y(N51) );
  NOR4BX1 U31 ( .AN(n12), .B(kld), .C(n13), .D(rcnt[0]), .Y(N49) );
  XNOR2X1 U32 ( .A(n2), .B(n15), .Y(n13) );
  OAI22X1 U33 ( .A0(n14), .A1(n7), .B0(n16), .B1(n17), .Y(N48) );
  INVX1 U34 ( .A(n18), .Y(n16) );
  NAND4X1 U35 ( .A(n19), .B(rcnt[0]), .C(n2), .D(n9), .Y(n7) );
  AOI21X1 U36 ( .A0(n10), .A1(n20), .B0(n17), .Y(N47) );
  NAND2X1 U37 ( .A(n18), .B(rcnt[0]), .Y(n20) );
  NAND3X1 U38 ( .A(n14), .B(n4), .C(n19), .Y(n10) );
  NOR2X1 U39 ( .A(n17), .B(n21), .Y(N46) );
  MXI2X1 U40 ( .A(n22), .B(n18), .S0(n4), .Y(n21) );
  NOR2X1 U41 ( .A(n19), .B(n14), .Y(n18) );
  INVX1 U42 ( .A(n12), .Y(n14) );
  INVX1 U43 ( .A(n15), .Y(n19) );
  NOR2X1 U44 ( .A(n12), .B(n15), .Y(n22) );
  XOR2X1 U45 ( .A(n27), .B(n23), .Y(n15) );
  NOR2X1 U46 ( .A(n5), .B(n24), .Y(n23) );
  NAND2X1 U47 ( .A(n11), .B(n9), .Y(n17) );
  INVX1 U48 ( .A(n2), .Y(n11) );
  XOR2X1 U49 ( .A(n24), .B(n5), .Y(n2) );
  OAI31X1 U50 ( .A0(n25), .A1(kld), .A2(n26), .B0(n8), .Y(N45) );
  NAND4X1 U51 ( .A(n26), .B(n25), .C(n9), .D(n6), .Y(n8) );
  OAI2BB1X1 U52 ( .A0N(n25), .A1N(n26), .B0(n9), .Y(N44) );
  INVX1 U53 ( .A(kld), .Y(n9) );
  XNOR2X1 U54 ( .A(rcnt[2]), .B(n12), .Y(n26) );
  OAI21XL U55 ( .A0(n12), .A1(n5), .B0(n24), .Y(n25) );
  NAND2X1 U56 ( .A(rcnt[1]), .B(rcnt[0]), .Y(n24) );
  XOR2X1 U57 ( .A(rcnt[1]), .B(n4), .Y(n12) );
endmodule


module aes_cipher_top ( clk, rst, ld, done, key, text_in, text_out );
  input [127:0] key;
  input [127:0] text_in;
  output [127:0] text_out;
  input clk, rst, ld;
  output done;
  wire   N21, N32, N33, N34, N35, N36, N37, N38, N39, N48, N49, N50, N51, N52,
         N53, N54, N55, N64, N65, N66, N67, N68, N69, N70, N71, N80, N81, N82,
         N83, N84, N85, N86, N87, N96, N97, N98, N99, N100, N101, N102, N103,
         N112, N113, N114, N115, N116, N117, N118, N119, N128, N129, N130,
         N131, N132, N133, N134, N135, N144, N145, N146, N147, N148, N149,
         N150, N151, N160, N161, N162, N163, N164, N165, N166, N167, N176,
         N177, N178, N179, N180, N181, N182, N183, N192, N193, N194, N195,
         N196, N197, N198, N199, N208, N209, N210, N211, N212, N213, N214,
         N215, N224, N225, N226, N227, N228, N229, N230, N231, N240, N241,
         N242, N243, N244, N245, N246, N247, N256, N257, N258, N259, N260,
         N261, N262, N263, N272, N273, N274, N275, N276, N277, N278, N279,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463,
         N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474,
         N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485,
         N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496,
         N497, N498, N499, N500, N501, N502, N503, n1, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         \u0/n265 , \u0/n264 , \u0/n263 , \u0/n262 , \u0/n261 , \u0/n260 ,
         \u0/n259 , \u0/n258 , \u0/n128 , \u0/n127 , \u0/n126 , \u0/n125 ,
         \u0/n124 , \u0/n123 , \u0/n122 , \u0/n121 , \u0/n120 , \u0/n119 ,
         \u0/n118 , \u0/n117 , \u0/n116 , \u0/n115 , \u0/n114 , \u0/n113 ,
         \u0/n112 , \u0/n111 , \u0/n110 , \u0/n109 , \u0/n108 , \u0/n107 ,
         \u0/n106 , \u0/n105 , \u0/n104 , \u0/n103 , \u0/n102 , \u0/n101 ,
         \u0/n100 , \u0/n99 , \u0/n98 , \u0/n97 , \u0/n96 , \u0/n95 , \u0/n94 ,
         \u0/n93 , \u0/n92 , \u0/n91 , \u0/n90 , \u0/n89 , \u0/n88 , \u0/n87 ,
         \u0/n86 , \u0/n85 , \u0/n84 , \u0/n83 , \u0/n82 , \u0/n81 , \u0/n80 ,
         \u0/n79 , \u0/n78 , \u0/n77 , \u0/n76 , \u0/n75 , \u0/n74 , \u0/n73 ,
         \u0/n72 , \u0/n71 , \u0/n70 , \u0/n69 , \u0/n68 , \u0/n67 , \u0/n66 ,
         \u0/n65 , \u0/n64 , \u0/n63 , \u0/n62 , \u0/n61 , \u0/n60 , \u0/n59 ,
         \u0/n58 , \u0/n57 , \u0/n56 , \u0/n55 , \u0/n54 , \u0/n53 , \u0/n52 ,
         \u0/n51 , \u0/n50 , \u0/n49 , \u0/n48 , \u0/n47 , \u0/n46 , \u0/n45 ,
         \u0/n44 , \u0/n43 , \u0/n42 , \u0/n41 , \u0/n40 , \u0/n39 , \u0/n38 ,
         \u0/n37 , \u0/n36 , \u0/n35 , \u0/n34 , \u0/n33 , \u0/n32 , \u0/n31 ,
         \u0/n30 , \u0/n29 , \u0/n28 , \u0/n27 , \u0/n26 , \u0/n25 , \u0/n24 ,
         \u0/n23 , \u0/n22 , \u0/n21 , \u0/n20 , \u0/n19 , \u0/n18 , \u0/n17 ,
         \u0/n16 , \u0/n15 , \u0/n14 , \u0/n13 , \u0/n12 , \u0/n11 , \u0/n10 ,
         \u0/n9 , \u0/n8 , \u0/n7 , \u0/n6 , \u0/n5 , \u0/n4 , \u0/n3 ,
         \u0/n2 , \u0/n1 , \u0/N239 , \u0/N238 , \u0/N237 , \u0/N236 ,
         \u0/N235 , \u0/N234 , \u0/N233 , \u0/N232 , \u0/N231 , \u0/N230 ,
         \u0/N229 , \u0/N228 , \u0/N227 , \u0/N226 , \u0/N225 , \u0/N224 ,
         \u0/N223 , \u0/N222 , \u0/N221 , \u0/N220 , \u0/N219 , \u0/N218 ,
         \u0/N217 , \u0/N216 , \u0/N215 , \u0/N214 , \u0/N213 , \u0/N212 ,
         \u0/N211 , \u0/N210 , \u0/N209 , \u0/N208 , \u0/N173 , \u0/N172 ,
         \u0/N171 , \u0/N170 , \u0/N169 , \u0/N168 , \u0/N167 , \u0/N166 ,
         \u0/N165 , \u0/N164 , \u0/N163 , \u0/N162 , \u0/N161 , \u0/N160 ,
         \u0/N159 , \u0/N158 , \u0/N157 , \u0/N156 , \u0/N155 , \u0/N154 ,
         \u0/N153 , \u0/N152 , \u0/N151 , \u0/N150 , \u0/N149 , \u0/N148 ,
         \u0/N147 , \u0/N146 , \u0/N145 , \u0/N144 , \u0/N143 , \u0/N142 ,
         \u0/N107 , \u0/N106 , \u0/N105 , \u0/N104 , \u0/N103 , \u0/N102 ,
         \u0/N101 , \u0/N100 , \u0/N99 , \u0/N98 , \u0/N97 , \u0/N96 ,
         \u0/N95 , \u0/N94 , \u0/N93 , \u0/N92 , \u0/N91 , \u0/N90 , \u0/N89 ,
         \u0/N88 , \u0/N87 , \u0/N86 , \u0/N85 , \u0/N84 , \u0/N83 , \u0/N82 ,
         \u0/N81 , \u0/N80 , \u0/N79 , \u0/N78 , \u0/N77 , \u0/N76 , \u0/N41 ,
         \u0/N40 , \u0/N39 , \u0/N38 , \u0/N37 , \u0/N36 , \u0/N35 , \u0/N34 ,
         \u0/N33 , \u0/N32 , \u0/N31 , \u0/N30 , \u0/N29 , \u0/N28 , \u0/N27 ,
         \u0/N26 , \u0/N25 , \u0/N24 , \u0/N23 , \u0/N22 , \u0/N21 , \u0/N20 ,
         \u0/N19 , \u0/N18 , \u0/N17 , \u0/N16 , \u0/N15 , \u0/N14 , \u0/N13 ,
         \u0/N12 , \u0/N11 , \u0/N10 , \us00/n358 , \us00/n357 , \us00/n356 ,
         \us00/n355 , \us00/n354 , \us00/n353 , \us00/n352 , \us00/n351 ,
         \us00/n350 , \us00/n349 , \us00/n348 , \us00/n347 , \us00/n346 ,
         \us00/n345 , \us00/n344 , \us00/n343 , \us00/n342 , \us00/n341 ,
         \us00/n340 , \us00/n339 , \us00/n338 , \us00/n337 , \us00/n336 ,
         \us00/n335 , \us00/n334 , \us00/n333 , \us00/n332 , \us00/n331 ,
         \us00/n330 , \us00/n329 , \us00/n328 , \us00/n327 , \us00/n326 ,
         \us00/n325 , \us00/n324 , \us00/n323 , \us00/n322 , \us00/n321 ,
         \us00/n320 , \us00/n319 , \us00/n318 , \us00/n317 , \us00/n316 ,
         \us00/n315 , \us00/n314 , \us00/n313 , \us00/n312 , \us00/n311 ,
         \us00/n310 , \us00/n309 , \us00/n308 , \us00/n307 , \us00/n306 ,
         \us00/n305 , \us00/n304 , \us00/n303 , \us00/n302 , \us00/n301 ,
         \us00/n300 , \us00/n299 , \us00/n298 , \us00/n297 , \us00/n296 ,
         \us00/n295 , \us00/n294 , \us00/n293 , \us00/n292 , \us00/n291 ,
         \us00/n290 , \us00/n289 , \us00/n288 , \us00/n287 , \us00/n286 ,
         \us00/n285 , \us00/n284 , \us00/n283 , \us00/n282 , \us00/n281 ,
         \us00/n280 , \us00/n279 , \us00/n278 , \us00/n277 , \us00/n276 ,
         \us00/n275 , \us00/n274 , \us00/n273 , \us00/n272 , \us00/n271 ,
         \us00/n270 , \us00/n269 , \us00/n268 , \us00/n267 , \us00/n266 ,
         \us00/n265 , \us00/n264 , \us00/n263 , \us00/n262 , \us00/n261 ,
         \us00/n260 , \us00/n259 , \us00/n258 , \us00/n257 , \us00/n256 ,
         \us00/n255 , \us00/n254 , \us00/n253 , \us00/n252 , \us00/n251 ,
         \us00/n250 , \us00/n249 , \us00/n248 , \us00/n247 , \us00/n246 ,
         \us00/n245 , \us00/n244 , \us00/n243 , \us00/n242 , \us00/n241 ,
         \us00/n240 , \us00/n239 , \us00/n238 , \us00/n237 , \us00/n236 ,
         \us00/n235 , \us00/n234 , \us00/n233 , \us00/n232 , \us00/n231 ,
         \us00/n230 , \us00/n229 , \us00/n228 , \us00/n227 , \us00/n226 ,
         \us00/n225 , \us00/n224 , \us00/n223 , \us00/n222 , \us00/n221 ,
         \us00/n220 , \us00/n219 , \us00/n218 , \us00/n217 , \us00/n216 ,
         \us00/n215 , \us00/n214 , \us00/n213 , \us00/n212 , \us00/n211 ,
         \us00/n210 , \us00/n209 , \us00/n208 , \us00/n207 , \us00/n206 ,
         \us00/n205 , \us00/n204 , \us00/n203 , \us00/n202 , \us00/n201 ,
         \us00/n200 , \us00/n199 , \us00/n198 , \us00/n197 , \us00/n196 ,
         \us00/n195 , \us00/n194 , \us00/n193 , \us00/n192 , \us00/n191 ,
         \us00/n190 , \us00/n189 , \us00/n188 , \us00/n187 , \us00/n186 ,
         \us00/n185 , \us00/n184 , \us00/n183 , \us00/n182 , \us00/n181 ,
         \us00/n180 , \us00/n179 , \us00/n178 , \us00/n177 , \us00/n176 ,
         \us00/n175 , \us00/n174 , \us00/n173 , \us00/n172 , \us00/n171 ,
         \us00/n170 , \us00/n169 , \us00/n168 , \us00/n167 , \us00/n166 ,
         \us00/n165 , \us00/n164 , \us00/n163 , \us00/n162 , \us00/n161 ,
         \us00/n160 , \us00/n159 , \us00/n158 , \us00/n157 , \us00/n156 ,
         \us00/n155 , \us00/n154 , \us00/n153 , \us00/n152 , \us00/n151 ,
         \us00/n150 , \us00/n149 , \us00/n148 , \us00/n147 , \us00/n146 ,
         \us00/n145 , \us00/n144 , \us00/n143 , \us00/n142 , \us00/n141 ,
         \us00/n140 , \us00/n139 , \us00/n138 , \us00/n137 , \us00/n136 ,
         \us00/n135 , \us00/n134 , \us00/n133 , \us00/n132 , \us00/n131 ,
         \us00/n130 , \us00/n129 , \us00/n128 , \us00/n127 , \us00/n126 ,
         \us00/n125 , \us00/n124 , \us00/n123 , \us00/n122 , \us00/n121 ,
         \us00/n120 , \us00/n119 , \us00/n118 , \us00/n117 , \us00/n116 ,
         \us00/n115 , \us00/n114 , \us00/n113 , \us00/n112 , \us00/n111 ,
         \us00/n110 , \us00/n109 , \us00/n108 , \us00/n107 , \us00/n106 ,
         \us00/n105 , \us00/n104 , \us00/n103 , \us00/n102 , \us00/n101 ,
         \us00/n100 , \us00/n99 , \us00/n98 , \us00/n97 , \us00/n96 ,
         \us00/n95 , \us00/n94 , \us00/n93 , \us00/n92 , \us00/n91 ,
         \us00/n90 , \us00/n89 , \us00/n88 , \us00/n87 , \us00/n86 ,
         \us00/n85 , \us00/n84 , \us00/n83 , \us00/n82 , \us00/n81 ,
         \us00/n80 , \us00/n79 , \us00/n78 , \us00/n77 , \us00/n76 ,
         \us00/n75 , \us00/n74 , \us00/n73 , \us00/n72 , \us00/n71 ,
         \us00/n70 , \us00/n69 , \us00/n68 , \us00/n67 , \us00/n66 ,
         \us00/n65 , \us00/n64 , \us00/n63 , \us00/n62 , \us00/n61 ,
         \us00/n60 , \us00/n59 , \us00/n58 , \us00/n57 , \us00/n56 ,
         \us00/n55 , \us00/n54 , \us00/n53 , \us00/n52 , \us00/n51 ,
         \us00/n50 , \us00/n49 , \us00/n48 , \us00/n47 , \us00/n46 ,
         \us00/n45 , \us00/n44 , \us00/n43 , \us00/n42 , \us00/n41 ,
         \us00/n40 , \us00/n39 , \us00/n38 , \us00/n37 , \us00/n36 ,
         \us00/n35 , \us00/n34 , \us00/n33 , \us00/n32 , \us00/n31 ,
         \us00/n30 , \us00/n29 , \us00/n28 , \us00/n27 , \us00/n26 ,
         \us00/n25 , \us00/n24 , \us00/n23 , \us00/n22 , \us00/n21 ,
         \us00/n20 , \us00/n19 , \us00/n18 , \us00/n17 , \us00/n16 ,
         \us00/n15 , \us00/n14 , \us00/n13 , \us00/n12 , \us00/n11 ,
         \us00/n10 , \us00/n9 , \us00/n8 , \us00/n7 , \us00/n6 , \us00/n5 ,
         \us00/n4 , \us00/n3 , \us00/n2 , \us00/n1 , \us01/n358 , \us01/n357 ,
         \us01/n356 , \us01/n355 , \us01/n354 , \us01/n353 , \us01/n352 ,
         \us01/n351 , \us01/n350 , \us01/n349 , \us01/n348 , \us01/n347 ,
         \us01/n346 , \us01/n345 , \us01/n344 , \us01/n343 , \us01/n342 ,
         \us01/n341 , \us01/n340 , \us01/n339 , \us01/n338 , \us01/n337 ,
         \us01/n336 , \us01/n335 , \us01/n334 , \us01/n333 , \us01/n332 ,
         \us01/n331 , \us01/n330 , \us01/n329 , \us01/n328 , \us01/n327 ,
         \us01/n326 , \us01/n325 , \us01/n324 , \us01/n323 , \us01/n322 ,
         \us01/n321 , \us01/n320 , \us01/n319 , \us01/n318 , \us01/n317 ,
         \us01/n316 , \us01/n315 , \us01/n314 , \us01/n313 , \us01/n312 ,
         \us01/n311 , \us01/n310 , \us01/n309 , \us01/n308 , \us01/n307 ,
         \us01/n306 , \us01/n305 , \us01/n304 , \us01/n303 , \us01/n302 ,
         \us01/n301 , \us01/n300 , \us01/n299 , \us01/n298 , \us01/n297 ,
         \us01/n296 , \us01/n295 , \us01/n294 , \us01/n293 , \us01/n292 ,
         \us01/n291 , \us01/n290 , \us01/n289 , \us01/n288 , \us01/n287 ,
         \us01/n286 , \us01/n285 , \us01/n284 , \us01/n283 , \us01/n282 ,
         \us01/n281 , \us01/n280 , \us01/n279 , \us01/n278 , \us01/n277 ,
         \us01/n276 , \us01/n275 , \us01/n274 , \us01/n273 , \us01/n272 ,
         \us01/n271 , \us01/n270 , \us01/n269 , \us01/n268 , \us01/n267 ,
         \us01/n266 , \us01/n265 , \us01/n264 , \us01/n263 , \us01/n262 ,
         \us01/n261 , \us01/n260 , \us01/n259 , \us01/n258 , \us01/n257 ,
         \us01/n256 , \us01/n255 , \us01/n254 , \us01/n253 , \us01/n252 ,
         \us01/n251 , \us01/n250 , \us01/n249 , \us01/n248 , \us01/n247 ,
         \us01/n246 , \us01/n245 , \us01/n244 , \us01/n243 , \us01/n242 ,
         \us01/n241 , \us01/n240 , \us01/n239 , \us01/n238 , \us01/n237 ,
         \us01/n236 , \us01/n235 , \us01/n234 , \us01/n233 , \us01/n232 ,
         \us01/n231 , \us01/n230 , \us01/n229 , \us01/n228 , \us01/n227 ,
         \us01/n226 , \us01/n225 , \us01/n224 , \us01/n223 , \us01/n222 ,
         \us01/n221 , \us01/n220 , \us01/n219 , \us01/n218 , \us01/n217 ,
         \us01/n216 , \us01/n215 , \us01/n214 , \us01/n213 , \us01/n212 ,
         \us01/n211 , \us01/n210 , \us01/n209 , \us01/n208 , \us01/n207 ,
         \us01/n206 , \us01/n205 , \us01/n204 , \us01/n203 , \us01/n202 ,
         \us01/n201 , \us01/n200 , \us01/n199 , \us01/n198 , \us01/n197 ,
         \us01/n196 , \us01/n195 , \us01/n194 , \us01/n193 , \us01/n192 ,
         \us01/n191 , \us01/n190 , \us01/n189 , \us01/n188 , \us01/n187 ,
         \us01/n186 , \us01/n185 , \us01/n184 , \us01/n183 , \us01/n182 ,
         \us01/n181 , \us01/n180 , \us01/n179 , \us01/n178 , \us01/n177 ,
         \us01/n176 , \us01/n175 , \us01/n174 , \us01/n173 , \us01/n172 ,
         \us01/n171 , \us01/n170 , \us01/n169 , \us01/n168 , \us01/n167 ,
         \us01/n166 , \us01/n165 , \us01/n164 , \us01/n163 , \us01/n162 ,
         \us01/n161 , \us01/n160 , \us01/n159 , \us01/n158 , \us01/n157 ,
         \us01/n156 , \us01/n155 , \us01/n154 , \us01/n153 , \us01/n152 ,
         \us01/n151 , \us01/n150 , \us01/n149 , \us01/n148 , \us01/n147 ,
         \us01/n146 , \us01/n145 , \us01/n144 , \us01/n143 , \us01/n142 ,
         \us01/n141 , \us01/n140 , \us01/n139 , \us01/n138 , \us01/n137 ,
         \us01/n136 , \us01/n135 , \us01/n134 , \us01/n133 , \us01/n132 ,
         \us01/n131 , \us01/n130 , \us01/n129 , \us01/n128 , \us01/n127 ,
         \us01/n126 , \us01/n125 , \us01/n124 , \us01/n123 , \us01/n122 ,
         \us01/n121 , \us01/n120 , \us01/n119 , \us01/n118 , \us01/n117 ,
         \us01/n116 , \us01/n115 , \us01/n114 , \us01/n113 , \us01/n112 ,
         \us01/n111 , \us01/n110 , \us01/n109 , \us01/n108 , \us01/n107 ,
         \us01/n106 , \us01/n105 , \us01/n104 , \us01/n103 , \us01/n102 ,
         \us01/n101 , \us01/n100 , \us01/n99 , \us01/n98 , \us01/n97 ,
         \us01/n96 , \us01/n95 , \us01/n94 , \us01/n93 , \us01/n92 ,
         \us01/n91 , \us01/n90 , \us01/n89 , \us01/n88 , \us01/n87 ,
         \us01/n86 , \us01/n85 , \us01/n84 , \us01/n83 , \us01/n82 ,
         \us01/n81 , \us01/n80 , \us01/n79 , \us01/n78 , \us01/n77 ,
         \us01/n76 , \us01/n75 , \us01/n74 , \us01/n73 , \us01/n72 ,
         \us01/n71 , \us01/n70 , \us01/n69 , \us01/n68 , \us01/n67 ,
         \us01/n66 , \us01/n65 , \us01/n64 , \us01/n63 , \us01/n62 ,
         \us01/n61 , \us01/n60 , \us01/n59 , \us01/n58 , \us01/n57 ,
         \us01/n56 , \us01/n55 , \us01/n54 , \us01/n53 , \us01/n52 ,
         \us01/n51 , \us01/n50 , \us01/n49 , \us01/n48 , \us01/n47 ,
         \us01/n46 , \us01/n45 , \us01/n44 , \us01/n43 , \us01/n42 ,
         \us01/n41 , \us01/n40 , \us01/n39 , \us01/n38 , \us01/n37 ,
         \us01/n36 , \us01/n35 , \us01/n34 , \us01/n33 , \us01/n32 ,
         \us01/n31 , \us01/n30 , \us01/n29 , \us01/n28 , \us01/n27 ,
         \us01/n26 , \us01/n25 , \us01/n24 , \us01/n23 , \us01/n22 ,
         \us01/n21 , \us01/n20 , \us01/n19 , \us01/n18 , \us01/n17 ,
         \us01/n16 , \us01/n15 , \us01/n14 , \us01/n13 , \us01/n12 ,
         \us01/n11 , \us01/n10 , \us01/n9 , \us01/n8 , \us01/n7 , \us01/n6 ,
         \us01/n5 , \us01/n4 , \us01/n3 , \us01/n2 , \us01/n1 , \us02/n358 ,
         \us02/n357 , \us02/n356 , \us02/n355 , \us02/n354 , \us02/n353 ,
         \us02/n352 , \us02/n351 , \us02/n350 , \us02/n349 , \us02/n348 ,
         \us02/n347 , \us02/n346 , \us02/n345 , \us02/n344 , \us02/n343 ,
         \us02/n342 , \us02/n341 , \us02/n340 , \us02/n339 , \us02/n338 ,
         \us02/n337 , \us02/n336 , \us02/n335 , \us02/n334 , \us02/n333 ,
         \us02/n332 , \us02/n331 , \us02/n330 , \us02/n329 , \us02/n328 ,
         \us02/n327 , \us02/n326 , \us02/n325 , \us02/n324 , \us02/n323 ,
         \us02/n322 , \us02/n321 , \us02/n320 , \us02/n319 , \us02/n318 ,
         \us02/n317 , \us02/n316 , \us02/n315 , \us02/n314 , \us02/n313 ,
         \us02/n312 , \us02/n311 , \us02/n310 , \us02/n309 , \us02/n308 ,
         \us02/n307 , \us02/n306 , \us02/n305 , \us02/n304 , \us02/n303 ,
         \us02/n302 , \us02/n301 , \us02/n300 , \us02/n299 , \us02/n298 ,
         \us02/n297 , \us02/n296 , \us02/n295 , \us02/n294 , \us02/n293 ,
         \us02/n292 , \us02/n291 , \us02/n290 , \us02/n289 , \us02/n288 ,
         \us02/n287 , \us02/n286 , \us02/n285 , \us02/n284 , \us02/n283 ,
         \us02/n282 , \us02/n281 , \us02/n280 , \us02/n279 , \us02/n278 ,
         \us02/n277 , \us02/n276 , \us02/n275 , \us02/n274 , \us02/n273 ,
         \us02/n272 , \us02/n271 , \us02/n270 , \us02/n269 , \us02/n268 ,
         \us02/n267 , \us02/n266 , \us02/n265 , \us02/n264 , \us02/n263 ,
         \us02/n262 , \us02/n261 , \us02/n260 , \us02/n259 , \us02/n258 ,
         \us02/n257 , \us02/n256 , \us02/n255 , \us02/n254 , \us02/n253 ,
         \us02/n252 , \us02/n251 , \us02/n250 , \us02/n249 , \us02/n248 ,
         \us02/n247 , \us02/n246 , \us02/n245 , \us02/n244 , \us02/n243 ,
         \us02/n242 , \us02/n241 , \us02/n240 , \us02/n239 , \us02/n238 ,
         \us02/n237 , \us02/n236 , \us02/n235 , \us02/n234 , \us02/n233 ,
         \us02/n232 , \us02/n231 , \us02/n230 , \us02/n229 , \us02/n228 ,
         \us02/n227 , \us02/n226 , \us02/n225 , \us02/n224 , \us02/n223 ,
         \us02/n222 , \us02/n221 , \us02/n220 , \us02/n219 , \us02/n218 ,
         \us02/n217 , \us02/n216 , \us02/n215 , \us02/n214 , \us02/n213 ,
         \us02/n212 , \us02/n211 , \us02/n210 , \us02/n209 , \us02/n208 ,
         \us02/n207 , \us02/n206 , \us02/n205 , \us02/n204 , \us02/n203 ,
         \us02/n202 , \us02/n201 , \us02/n200 , \us02/n199 , \us02/n198 ,
         \us02/n197 , \us02/n196 , \us02/n195 , \us02/n194 , \us02/n193 ,
         \us02/n192 , \us02/n191 , \us02/n190 , \us02/n189 , \us02/n188 ,
         \us02/n187 , \us02/n186 , \us02/n185 , \us02/n184 , \us02/n183 ,
         \us02/n182 , \us02/n181 , \us02/n180 , \us02/n179 , \us02/n178 ,
         \us02/n177 , \us02/n176 , \us02/n175 , \us02/n174 , \us02/n173 ,
         \us02/n172 , \us02/n171 , \us02/n170 , \us02/n169 , \us02/n168 ,
         \us02/n167 , \us02/n166 , \us02/n165 , \us02/n164 , \us02/n163 ,
         \us02/n162 , \us02/n161 , \us02/n160 , \us02/n159 , \us02/n158 ,
         \us02/n157 , \us02/n156 , \us02/n155 , \us02/n154 , \us02/n153 ,
         \us02/n152 , \us02/n151 , \us02/n150 , \us02/n149 , \us02/n148 ,
         \us02/n147 , \us02/n146 , \us02/n145 , \us02/n144 , \us02/n143 ,
         \us02/n142 , \us02/n141 , \us02/n140 , \us02/n139 , \us02/n138 ,
         \us02/n137 , \us02/n136 , \us02/n135 , \us02/n134 , \us02/n133 ,
         \us02/n132 , \us02/n131 , \us02/n130 , \us02/n129 , \us02/n128 ,
         \us02/n127 , \us02/n126 , \us02/n125 , \us02/n124 , \us02/n123 ,
         \us02/n122 , \us02/n121 , \us02/n120 , \us02/n119 , \us02/n118 ,
         \us02/n117 , \us02/n116 , \us02/n115 , \us02/n114 , \us02/n113 ,
         \us02/n112 , \us02/n111 , \us02/n110 , \us02/n109 , \us02/n108 ,
         \us02/n107 , \us02/n106 , \us02/n105 , \us02/n104 , \us02/n103 ,
         \us02/n102 , \us02/n101 , \us02/n100 , \us02/n99 , \us02/n98 ,
         \us02/n97 , \us02/n96 , \us02/n95 , \us02/n94 , \us02/n93 ,
         \us02/n92 , \us02/n91 , \us02/n90 , \us02/n89 , \us02/n88 ,
         \us02/n87 , \us02/n86 , \us02/n85 , \us02/n84 , \us02/n83 ,
         \us02/n82 , \us02/n81 , \us02/n80 , \us02/n79 , \us02/n78 ,
         \us02/n77 , \us02/n76 , \us02/n75 , \us02/n74 , \us02/n73 ,
         \us02/n72 , \us02/n71 , \us02/n70 , \us02/n69 , \us02/n68 ,
         \us02/n67 , \us02/n66 , \us02/n65 , \us02/n64 , \us02/n63 ,
         \us02/n62 , \us02/n61 , \us02/n60 , \us02/n59 , \us02/n58 ,
         \us02/n57 , \us02/n56 , \us02/n55 , \us02/n54 , \us02/n53 ,
         \us02/n52 , \us02/n51 , \us02/n50 , \us02/n49 , \us02/n48 ,
         \us02/n47 , \us02/n46 , \us02/n45 , \us02/n44 , \us02/n43 ,
         \us02/n42 , \us02/n41 , \us02/n40 , \us02/n39 , \us02/n38 ,
         \us02/n37 , \us02/n36 , \us02/n35 , \us02/n34 , \us02/n33 ,
         \us02/n32 , \us02/n31 , \us02/n30 , \us02/n29 , \us02/n28 ,
         \us02/n27 , \us02/n26 , \us02/n25 , \us02/n24 , \us02/n23 ,
         \us02/n22 , \us02/n21 , \us02/n20 , \us02/n19 , \us02/n18 ,
         \us02/n17 , \us02/n16 , \us02/n15 , \us02/n14 , \us02/n13 ,
         \us02/n12 , \us02/n11 , \us02/n10 , \us02/n9 , \us02/n8 , \us02/n7 ,
         \us02/n6 , \us02/n5 , \us02/n4 , \us02/n3 , \us02/n2 , \us02/n1 ,
         \us03/n358 , \us03/n357 , \us03/n356 , \us03/n355 , \us03/n354 ,
         \us03/n353 , \us03/n352 , \us03/n351 , \us03/n350 , \us03/n349 ,
         \us03/n348 , \us03/n347 , \us03/n346 , \us03/n345 , \us03/n344 ,
         \us03/n343 , \us03/n342 , \us03/n341 , \us03/n340 , \us03/n339 ,
         \us03/n338 , \us03/n337 , \us03/n336 , \us03/n335 , \us03/n334 ,
         \us03/n333 , \us03/n332 , \us03/n331 , \us03/n330 , \us03/n329 ,
         \us03/n328 , \us03/n327 , \us03/n326 , \us03/n325 , \us03/n324 ,
         \us03/n323 , \us03/n322 , \us03/n321 , \us03/n320 , \us03/n319 ,
         \us03/n318 , \us03/n317 , \us03/n316 , \us03/n315 , \us03/n314 ,
         \us03/n313 , \us03/n312 , \us03/n311 , \us03/n310 , \us03/n309 ,
         \us03/n308 , \us03/n307 , \us03/n306 , \us03/n305 , \us03/n304 ,
         \us03/n303 , \us03/n302 , \us03/n301 , \us03/n300 , \us03/n299 ,
         \us03/n298 , \us03/n297 , \us03/n296 , \us03/n295 , \us03/n294 ,
         \us03/n293 , \us03/n292 , \us03/n291 , \us03/n290 , \us03/n289 ,
         \us03/n288 , \us03/n287 , \us03/n286 , \us03/n285 , \us03/n284 ,
         \us03/n283 , \us03/n282 , \us03/n281 , \us03/n280 , \us03/n279 ,
         \us03/n278 , \us03/n277 , \us03/n276 , \us03/n275 , \us03/n274 ,
         \us03/n273 , \us03/n272 , \us03/n271 , \us03/n270 , \us03/n269 ,
         \us03/n268 , \us03/n267 , \us03/n266 , \us03/n265 , \us03/n264 ,
         \us03/n263 , \us03/n262 , \us03/n261 , \us03/n260 , \us03/n259 ,
         \us03/n258 , \us03/n257 , \us03/n256 , \us03/n255 , \us03/n254 ,
         \us03/n253 , \us03/n252 , \us03/n251 , \us03/n250 , \us03/n249 ,
         \us03/n248 , \us03/n247 , \us03/n246 , \us03/n245 , \us03/n244 ,
         \us03/n243 , \us03/n242 , \us03/n241 , \us03/n240 , \us03/n239 ,
         \us03/n238 , \us03/n237 , \us03/n236 , \us03/n235 , \us03/n234 ,
         \us03/n233 , \us03/n232 , \us03/n231 , \us03/n230 , \us03/n229 ,
         \us03/n228 , \us03/n227 , \us03/n226 , \us03/n225 , \us03/n224 ,
         \us03/n223 , \us03/n222 , \us03/n221 , \us03/n220 , \us03/n219 ,
         \us03/n218 , \us03/n217 , \us03/n216 , \us03/n215 , \us03/n214 ,
         \us03/n213 , \us03/n212 , \us03/n211 , \us03/n210 , \us03/n209 ,
         \us03/n208 , \us03/n207 , \us03/n206 , \us03/n205 , \us03/n204 ,
         \us03/n203 , \us03/n202 , \us03/n201 , \us03/n200 , \us03/n199 ,
         \us03/n198 , \us03/n197 , \us03/n196 , \us03/n195 , \us03/n194 ,
         \us03/n193 , \us03/n192 , \us03/n191 , \us03/n190 , \us03/n189 ,
         \us03/n188 , \us03/n187 , \us03/n186 , \us03/n185 , \us03/n184 ,
         \us03/n183 , \us03/n182 , \us03/n181 , \us03/n180 , \us03/n179 ,
         \us03/n178 , \us03/n177 , \us03/n176 , \us03/n175 , \us03/n174 ,
         \us03/n173 , \us03/n172 , \us03/n171 , \us03/n170 , \us03/n169 ,
         \us03/n168 , \us03/n167 , \us03/n166 , \us03/n165 , \us03/n164 ,
         \us03/n163 , \us03/n162 , \us03/n161 , \us03/n160 , \us03/n159 ,
         \us03/n158 , \us03/n157 , \us03/n156 , \us03/n155 , \us03/n154 ,
         \us03/n153 , \us03/n152 , \us03/n151 , \us03/n150 , \us03/n149 ,
         \us03/n148 , \us03/n147 , \us03/n146 , \us03/n145 , \us03/n144 ,
         \us03/n143 , \us03/n142 , \us03/n141 , \us03/n140 , \us03/n139 ,
         \us03/n138 , \us03/n137 , \us03/n136 , \us03/n135 , \us03/n134 ,
         \us03/n133 , \us03/n132 , \us03/n131 , \us03/n130 , \us03/n129 ,
         \us03/n128 , \us03/n127 , \us03/n126 , \us03/n125 , \us03/n124 ,
         \us03/n123 , \us03/n122 , \us03/n121 , \us03/n120 , \us03/n119 ,
         \us03/n118 , \us03/n117 , \us03/n116 , \us03/n115 , \us03/n114 ,
         \us03/n113 , \us03/n112 , \us03/n111 , \us03/n110 , \us03/n109 ,
         \us03/n108 , \us03/n107 , \us03/n106 , \us03/n105 , \us03/n104 ,
         \us03/n103 , \us03/n102 , \us03/n101 , \us03/n100 , \us03/n99 ,
         \us03/n98 , \us03/n97 , \us03/n96 , \us03/n95 , \us03/n94 ,
         \us03/n93 , \us03/n92 , \us03/n91 , \us03/n90 , \us03/n89 ,
         \us03/n88 , \us03/n87 , \us03/n86 , \us03/n85 , \us03/n84 ,
         \us03/n83 , \us03/n82 , \us03/n81 , \us03/n80 , \us03/n79 ,
         \us03/n78 , \us03/n77 , \us03/n76 , \us03/n75 , \us03/n74 ,
         \us03/n73 , \us03/n72 , \us03/n71 , \us03/n70 , \us03/n69 ,
         \us03/n68 , \us03/n67 , \us03/n66 , \us03/n65 , \us03/n64 ,
         \us03/n63 , \us03/n62 , \us03/n61 , \us03/n60 , \us03/n59 ,
         \us03/n58 , \us03/n57 , \us03/n56 , \us03/n55 , \us03/n54 ,
         \us03/n53 , \us03/n52 , \us03/n51 , \us03/n50 , \us03/n49 ,
         \us03/n48 , \us03/n47 , \us03/n46 , \us03/n45 , \us03/n44 ,
         \us03/n43 , \us03/n42 , \us03/n41 , \us03/n40 , \us03/n39 ,
         \us03/n38 , \us03/n37 , \us03/n36 , \us03/n35 , \us03/n34 ,
         \us03/n33 , \us03/n32 , \us03/n31 , \us03/n30 , \us03/n29 ,
         \us03/n28 , \us03/n27 , \us03/n26 , \us03/n25 , \us03/n24 ,
         \us03/n23 , \us03/n22 , \us03/n21 , \us03/n20 , \us03/n19 ,
         \us03/n18 , \us03/n17 , \us03/n16 , \us03/n15 , \us03/n14 ,
         \us03/n13 , \us03/n12 , \us03/n11 , \us03/n10 , \us03/n9 , \us03/n8 ,
         \us03/n7 , \us03/n6 , \us03/n5 , \us03/n4 , \us03/n3 , \us03/n2 ,
         \us03/n1 , \us10/n358 , \us10/n357 , \us10/n356 , \us10/n355 ,
         \us10/n354 , \us10/n353 , \us10/n352 , \us10/n351 , \us10/n350 ,
         \us10/n349 , \us10/n348 , \us10/n347 , \us10/n346 , \us10/n345 ,
         \us10/n344 , \us10/n343 , \us10/n342 , \us10/n341 , \us10/n340 ,
         \us10/n339 , \us10/n338 , \us10/n337 , \us10/n336 , \us10/n335 ,
         \us10/n334 , \us10/n333 , \us10/n332 , \us10/n331 , \us10/n330 ,
         \us10/n329 , \us10/n328 , \us10/n327 , \us10/n326 , \us10/n325 ,
         \us10/n324 , \us10/n323 , \us10/n322 , \us10/n321 , \us10/n320 ,
         \us10/n319 , \us10/n318 , \us10/n317 , \us10/n316 , \us10/n315 ,
         \us10/n314 , \us10/n313 , \us10/n312 , \us10/n311 , \us10/n310 ,
         \us10/n309 , \us10/n308 , \us10/n307 , \us10/n306 , \us10/n305 ,
         \us10/n304 , \us10/n303 , \us10/n302 , \us10/n301 , \us10/n300 ,
         \us10/n299 , \us10/n298 , \us10/n297 , \us10/n296 , \us10/n295 ,
         \us10/n294 , \us10/n293 , \us10/n292 , \us10/n291 , \us10/n290 ,
         \us10/n289 , \us10/n288 , \us10/n287 , \us10/n286 , \us10/n285 ,
         \us10/n284 , \us10/n283 , \us10/n282 , \us10/n281 , \us10/n280 ,
         \us10/n279 , \us10/n278 , \us10/n277 , \us10/n276 , \us10/n275 ,
         \us10/n274 , \us10/n273 , \us10/n272 , \us10/n271 , \us10/n270 ,
         \us10/n269 , \us10/n268 , \us10/n267 , \us10/n266 , \us10/n265 ,
         \us10/n264 , \us10/n263 , \us10/n262 , \us10/n261 , \us10/n260 ,
         \us10/n259 , \us10/n258 , \us10/n257 , \us10/n256 , \us10/n255 ,
         \us10/n254 , \us10/n253 , \us10/n252 , \us10/n251 , \us10/n250 ,
         \us10/n249 , \us10/n248 , \us10/n247 , \us10/n246 , \us10/n245 ,
         \us10/n244 , \us10/n243 , \us10/n242 , \us10/n241 , \us10/n240 ,
         \us10/n239 , \us10/n238 , \us10/n237 , \us10/n236 , \us10/n235 ,
         \us10/n234 , \us10/n233 , \us10/n232 , \us10/n231 , \us10/n230 ,
         \us10/n229 , \us10/n228 , \us10/n227 , \us10/n226 , \us10/n225 ,
         \us10/n224 , \us10/n223 , \us10/n222 , \us10/n221 , \us10/n220 ,
         \us10/n219 , \us10/n218 , \us10/n217 , \us10/n216 , \us10/n215 ,
         \us10/n214 , \us10/n213 , \us10/n212 , \us10/n211 , \us10/n210 ,
         \us10/n209 , \us10/n208 , \us10/n207 , \us10/n206 , \us10/n205 ,
         \us10/n204 , \us10/n203 , \us10/n202 , \us10/n201 , \us10/n200 ,
         \us10/n199 , \us10/n198 , \us10/n197 , \us10/n196 , \us10/n195 ,
         \us10/n194 , \us10/n193 , \us10/n192 , \us10/n191 , \us10/n190 ,
         \us10/n189 , \us10/n188 , \us10/n187 , \us10/n186 , \us10/n185 ,
         \us10/n184 , \us10/n183 , \us10/n182 , \us10/n181 , \us10/n180 ,
         \us10/n179 , \us10/n178 , \us10/n177 , \us10/n176 , \us10/n175 ,
         \us10/n174 , \us10/n173 , \us10/n172 , \us10/n171 , \us10/n170 ,
         \us10/n169 , \us10/n168 , \us10/n167 , \us10/n166 , \us10/n165 ,
         \us10/n164 , \us10/n163 , \us10/n162 , \us10/n161 , \us10/n160 ,
         \us10/n159 , \us10/n158 , \us10/n157 , \us10/n156 , \us10/n155 ,
         \us10/n154 , \us10/n153 , \us10/n152 , \us10/n151 , \us10/n150 ,
         \us10/n149 , \us10/n148 , \us10/n147 , \us10/n146 , \us10/n145 ,
         \us10/n144 , \us10/n143 , \us10/n142 , \us10/n141 , \us10/n140 ,
         \us10/n139 , \us10/n138 , \us10/n137 , \us10/n136 , \us10/n135 ,
         \us10/n134 , \us10/n133 , \us10/n132 , \us10/n131 , \us10/n130 ,
         \us10/n129 , \us10/n128 , \us10/n127 , \us10/n126 , \us10/n125 ,
         \us10/n124 , \us10/n123 , \us10/n122 , \us10/n121 , \us10/n120 ,
         \us10/n119 , \us10/n118 , \us10/n117 , \us10/n116 , \us10/n115 ,
         \us10/n114 , \us10/n113 , \us10/n112 , \us10/n111 , \us10/n110 ,
         \us10/n109 , \us10/n108 , \us10/n107 , \us10/n106 , \us10/n105 ,
         \us10/n104 , \us10/n103 , \us10/n102 , \us10/n101 , \us10/n100 ,
         \us10/n99 , \us10/n98 , \us10/n97 , \us10/n96 , \us10/n95 ,
         \us10/n94 , \us10/n93 , \us10/n92 , \us10/n91 , \us10/n90 ,
         \us10/n89 , \us10/n88 , \us10/n87 , \us10/n86 , \us10/n85 ,
         \us10/n84 , \us10/n83 , \us10/n82 , \us10/n81 , \us10/n80 ,
         \us10/n79 , \us10/n78 , \us10/n77 , \us10/n76 , \us10/n75 ,
         \us10/n74 , \us10/n73 , \us10/n72 , \us10/n71 , \us10/n70 ,
         \us10/n69 , \us10/n68 , \us10/n67 , \us10/n66 , \us10/n65 ,
         \us10/n64 , \us10/n63 , \us10/n62 , \us10/n61 , \us10/n60 ,
         \us10/n59 , \us10/n58 , \us10/n57 , \us10/n56 , \us10/n55 ,
         \us10/n54 , \us10/n53 , \us10/n52 , \us10/n51 , \us10/n50 ,
         \us10/n49 , \us10/n48 , \us10/n47 , \us10/n46 , \us10/n45 ,
         \us10/n44 , \us10/n43 , \us10/n42 , \us10/n41 , \us10/n40 ,
         \us10/n39 , \us10/n38 , \us10/n37 , \us10/n36 , \us10/n35 ,
         \us10/n34 , \us10/n33 , \us10/n32 , \us10/n31 , \us10/n30 ,
         \us10/n29 , \us10/n28 , \us10/n27 , \us10/n26 , \us10/n25 ,
         \us10/n24 , \us10/n23 , \us10/n22 , \us10/n21 , \us10/n20 ,
         \us10/n19 , \us10/n18 , \us10/n17 , \us10/n16 , \us10/n15 ,
         \us10/n14 , \us10/n13 , \us10/n12 , \us10/n11 , \us10/n10 , \us10/n9 ,
         \us10/n8 , \us10/n7 , \us10/n6 , \us10/n5 , \us10/n4 , \us10/n3 ,
         \us10/n2 , \us10/n1 , \us11/n358 , \us11/n357 , \us11/n356 ,
         \us11/n355 , \us11/n354 , \us11/n353 , \us11/n352 , \us11/n351 ,
         \us11/n350 , \us11/n349 , \us11/n348 , \us11/n347 , \us11/n346 ,
         \us11/n345 , \us11/n344 , \us11/n343 , \us11/n342 , \us11/n341 ,
         \us11/n340 , \us11/n339 , \us11/n338 , \us11/n337 , \us11/n336 ,
         \us11/n335 , \us11/n334 , \us11/n333 , \us11/n332 , \us11/n331 ,
         \us11/n330 , \us11/n329 , \us11/n328 , \us11/n327 , \us11/n326 ,
         \us11/n325 , \us11/n324 , \us11/n323 , \us11/n322 , \us11/n321 ,
         \us11/n320 , \us11/n319 , \us11/n318 , \us11/n317 , \us11/n316 ,
         \us11/n315 , \us11/n314 , \us11/n313 , \us11/n312 , \us11/n311 ,
         \us11/n310 , \us11/n309 , \us11/n308 , \us11/n307 , \us11/n306 ,
         \us11/n305 , \us11/n304 , \us11/n303 , \us11/n302 , \us11/n301 ,
         \us11/n300 , \us11/n299 , \us11/n298 , \us11/n297 , \us11/n296 ,
         \us11/n295 , \us11/n294 , \us11/n293 , \us11/n292 , \us11/n291 ,
         \us11/n290 , \us11/n289 , \us11/n288 , \us11/n287 , \us11/n286 ,
         \us11/n285 , \us11/n284 , \us11/n283 , \us11/n282 , \us11/n281 ,
         \us11/n280 , \us11/n279 , \us11/n278 , \us11/n277 , \us11/n276 ,
         \us11/n275 , \us11/n274 , \us11/n273 , \us11/n272 , \us11/n271 ,
         \us11/n270 , \us11/n269 , \us11/n268 , \us11/n267 , \us11/n266 ,
         \us11/n265 , \us11/n264 , \us11/n263 , \us11/n262 , \us11/n261 ,
         \us11/n260 , \us11/n259 , \us11/n258 , \us11/n257 , \us11/n256 ,
         \us11/n255 , \us11/n254 , \us11/n253 , \us11/n252 , \us11/n251 ,
         \us11/n250 , \us11/n249 , \us11/n248 , \us11/n247 , \us11/n246 ,
         \us11/n245 , \us11/n244 , \us11/n243 , \us11/n242 , \us11/n241 ,
         \us11/n240 , \us11/n239 , \us11/n238 , \us11/n237 , \us11/n236 ,
         \us11/n235 , \us11/n234 , \us11/n233 , \us11/n232 , \us11/n231 ,
         \us11/n230 , \us11/n229 , \us11/n228 , \us11/n227 , \us11/n226 ,
         \us11/n225 , \us11/n224 , \us11/n223 , \us11/n222 , \us11/n221 ,
         \us11/n220 , \us11/n219 , \us11/n218 , \us11/n217 , \us11/n216 ,
         \us11/n215 , \us11/n214 , \us11/n213 , \us11/n212 , \us11/n211 ,
         \us11/n210 , \us11/n209 , \us11/n208 , \us11/n207 , \us11/n206 ,
         \us11/n205 , \us11/n204 , \us11/n203 , \us11/n202 , \us11/n201 ,
         \us11/n200 , \us11/n199 , \us11/n198 , \us11/n197 , \us11/n196 ,
         \us11/n195 , \us11/n194 , \us11/n193 , \us11/n192 , \us11/n191 ,
         \us11/n190 , \us11/n189 , \us11/n188 , \us11/n187 , \us11/n186 ,
         \us11/n185 , \us11/n184 , \us11/n183 , \us11/n182 , \us11/n181 ,
         \us11/n180 , \us11/n179 , \us11/n178 , \us11/n177 , \us11/n176 ,
         \us11/n175 , \us11/n174 , \us11/n173 , \us11/n172 , \us11/n171 ,
         \us11/n170 , \us11/n169 , \us11/n168 , \us11/n167 , \us11/n166 ,
         \us11/n165 , \us11/n164 , \us11/n163 , \us11/n162 , \us11/n161 ,
         \us11/n160 , \us11/n159 , \us11/n158 , \us11/n157 , \us11/n156 ,
         \us11/n155 , \us11/n154 , \us11/n153 , \us11/n152 , \us11/n151 ,
         \us11/n150 , \us11/n149 , \us11/n148 , \us11/n147 , \us11/n146 ,
         \us11/n145 , \us11/n144 , \us11/n143 , \us11/n142 , \us11/n141 ,
         \us11/n140 , \us11/n139 , \us11/n138 , \us11/n137 , \us11/n136 ,
         \us11/n135 , \us11/n134 , \us11/n133 , \us11/n132 , \us11/n131 ,
         \us11/n130 , \us11/n129 , \us11/n128 , \us11/n127 , \us11/n126 ,
         \us11/n125 , \us11/n124 , \us11/n123 , \us11/n122 , \us11/n121 ,
         \us11/n120 , \us11/n119 , \us11/n118 , \us11/n117 , \us11/n116 ,
         \us11/n115 , \us11/n114 , \us11/n113 , \us11/n112 , \us11/n111 ,
         \us11/n110 , \us11/n109 , \us11/n108 , \us11/n107 , \us11/n106 ,
         \us11/n105 , \us11/n104 , \us11/n103 , \us11/n102 , \us11/n101 ,
         \us11/n100 , \us11/n99 , \us11/n98 , \us11/n97 , \us11/n96 ,
         \us11/n95 , \us11/n94 , \us11/n93 , \us11/n92 , \us11/n91 ,
         \us11/n90 , \us11/n89 , \us11/n88 , \us11/n87 , \us11/n86 ,
         \us11/n85 , \us11/n84 , \us11/n83 , \us11/n82 , \us11/n81 ,
         \us11/n80 , \us11/n79 , \us11/n78 , \us11/n77 , \us11/n76 ,
         \us11/n75 , \us11/n74 , \us11/n73 , \us11/n72 , \us11/n71 ,
         \us11/n70 , \us11/n69 , \us11/n68 , \us11/n67 , \us11/n66 ,
         \us11/n65 , \us11/n64 , \us11/n63 , \us11/n62 , \us11/n61 ,
         \us11/n60 , \us11/n59 , \us11/n58 , \us11/n57 , \us11/n56 ,
         \us11/n55 , \us11/n54 , \us11/n53 , \us11/n52 , \us11/n51 ,
         \us11/n50 , \us11/n49 , \us11/n48 , \us11/n47 , \us11/n46 ,
         \us11/n45 , \us11/n44 , \us11/n43 , \us11/n42 , \us11/n41 ,
         \us11/n40 , \us11/n39 , \us11/n38 , \us11/n37 , \us11/n36 ,
         \us11/n35 , \us11/n34 , \us11/n33 , \us11/n32 , \us11/n31 ,
         \us11/n30 , \us11/n29 , \us11/n28 , \us11/n27 , \us11/n26 ,
         \us11/n25 , \us11/n24 , \us11/n23 , \us11/n22 , \us11/n21 ,
         \us11/n20 , \us11/n19 , \us11/n18 , \us11/n17 , \us11/n16 ,
         \us11/n15 , \us11/n14 , \us11/n13 , \us11/n12 , \us11/n11 ,
         \us11/n10 , \us11/n9 , \us11/n8 , \us11/n7 , \us11/n6 , \us11/n5 ,
         \us11/n4 , \us11/n3 , \us11/n2 , \us11/n1 , \us12/n358 , \us12/n357 ,
         \us12/n356 , \us12/n355 , \us12/n354 , \us12/n353 , \us12/n352 ,
         \us12/n351 , \us12/n350 , \us12/n349 , \us12/n348 , \us12/n347 ,
         \us12/n346 , \us12/n345 , \us12/n344 , \us12/n343 , \us12/n342 ,
         \us12/n341 , \us12/n340 , \us12/n339 , \us12/n338 , \us12/n337 ,
         \us12/n336 , \us12/n335 , \us12/n334 , \us12/n333 , \us12/n332 ,
         \us12/n331 , \us12/n330 , \us12/n329 , \us12/n328 , \us12/n327 ,
         \us12/n326 , \us12/n325 , \us12/n324 , \us12/n323 , \us12/n322 ,
         \us12/n321 , \us12/n320 , \us12/n319 , \us12/n318 , \us12/n317 ,
         \us12/n316 , \us12/n315 , \us12/n314 , \us12/n313 , \us12/n312 ,
         \us12/n311 , \us12/n310 , \us12/n309 , \us12/n308 , \us12/n307 ,
         \us12/n306 , \us12/n305 , \us12/n304 , \us12/n303 , \us12/n302 ,
         \us12/n301 , \us12/n300 , \us12/n299 , \us12/n298 , \us12/n297 ,
         \us12/n296 , \us12/n295 , \us12/n294 , \us12/n293 , \us12/n292 ,
         \us12/n291 , \us12/n290 , \us12/n289 , \us12/n288 , \us12/n287 ,
         \us12/n286 , \us12/n285 , \us12/n284 , \us12/n283 , \us12/n282 ,
         \us12/n281 , \us12/n280 , \us12/n279 , \us12/n278 , \us12/n277 ,
         \us12/n276 , \us12/n275 , \us12/n274 , \us12/n273 , \us12/n272 ,
         \us12/n271 , \us12/n270 , \us12/n269 , \us12/n268 , \us12/n267 ,
         \us12/n266 , \us12/n265 , \us12/n264 , \us12/n263 , \us12/n262 ,
         \us12/n261 , \us12/n260 , \us12/n259 , \us12/n258 , \us12/n257 ,
         \us12/n256 , \us12/n255 , \us12/n254 , \us12/n253 , \us12/n252 ,
         \us12/n251 , \us12/n250 , \us12/n249 , \us12/n248 , \us12/n247 ,
         \us12/n246 , \us12/n245 , \us12/n244 , \us12/n243 , \us12/n242 ,
         \us12/n241 , \us12/n240 , \us12/n239 , \us12/n238 , \us12/n237 ,
         \us12/n236 , \us12/n235 , \us12/n234 , \us12/n233 , \us12/n232 ,
         \us12/n231 , \us12/n230 , \us12/n229 , \us12/n228 , \us12/n227 ,
         \us12/n226 , \us12/n225 , \us12/n224 , \us12/n223 , \us12/n222 ,
         \us12/n221 , \us12/n220 , \us12/n219 , \us12/n218 , \us12/n217 ,
         \us12/n216 , \us12/n215 , \us12/n214 , \us12/n213 , \us12/n212 ,
         \us12/n211 , \us12/n210 , \us12/n209 , \us12/n208 , \us12/n207 ,
         \us12/n206 , \us12/n205 , \us12/n204 , \us12/n203 , \us12/n202 ,
         \us12/n201 , \us12/n200 , \us12/n199 , \us12/n198 , \us12/n197 ,
         \us12/n196 , \us12/n195 , \us12/n194 , \us12/n193 , \us12/n192 ,
         \us12/n191 , \us12/n190 , \us12/n189 , \us12/n188 , \us12/n187 ,
         \us12/n186 , \us12/n185 , \us12/n184 , \us12/n183 , \us12/n182 ,
         \us12/n181 , \us12/n180 , \us12/n179 , \us12/n178 , \us12/n177 ,
         \us12/n176 , \us12/n175 , \us12/n174 , \us12/n173 , \us12/n172 ,
         \us12/n171 , \us12/n170 , \us12/n169 , \us12/n168 , \us12/n167 ,
         \us12/n166 , \us12/n165 , \us12/n164 , \us12/n163 , \us12/n162 ,
         \us12/n161 , \us12/n160 , \us12/n159 , \us12/n158 , \us12/n157 ,
         \us12/n156 , \us12/n155 , \us12/n154 , \us12/n153 , \us12/n152 ,
         \us12/n151 , \us12/n150 , \us12/n149 , \us12/n148 , \us12/n147 ,
         \us12/n146 , \us12/n145 , \us12/n144 , \us12/n143 , \us12/n142 ,
         \us12/n141 , \us12/n140 , \us12/n139 , \us12/n138 , \us12/n137 ,
         \us12/n136 , \us12/n135 , \us12/n134 , \us12/n133 , \us12/n132 ,
         \us12/n131 , \us12/n130 , \us12/n129 , \us12/n128 , \us12/n127 ,
         \us12/n126 , \us12/n125 , \us12/n124 , \us12/n123 , \us12/n122 ,
         \us12/n121 , \us12/n120 , \us12/n119 , \us12/n118 , \us12/n117 ,
         \us12/n116 , \us12/n115 , \us12/n114 , \us12/n113 , \us12/n112 ,
         \us12/n111 , \us12/n110 , \us12/n109 , \us12/n108 , \us12/n107 ,
         \us12/n106 , \us12/n105 , \us12/n104 , \us12/n103 , \us12/n102 ,
         \us12/n101 , \us12/n100 , \us12/n99 , \us12/n98 , \us12/n97 ,
         \us12/n96 , \us12/n95 , \us12/n94 , \us12/n93 , \us12/n92 ,
         \us12/n91 , \us12/n90 , \us12/n89 , \us12/n88 , \us12/n87 ,
         \us12/n86 , \us12/n85 , \us12/n84 , \us12/n83 , \us12/n82 ,
         \us12/n81 , \us12/n80 , \us12/n79 , \us12/n78 , \us12/n77 ,
         \us12/n76 , \us12/n75 , \us12/n74 , \us12/n73 , \us12/n72 ,
         \us12/n71 , \us12/n70 , \us12/n69 , \us12/n68 , \us12/n67 ,
         \us12/n66 , \us12/n65 , \us12/n64 , \us12/n63 , \us12/n62 ,
         \us12/n61 , \us12/n60 , \us12/n59 , \us12/n58 , \us12/n57 ,
         \us12/n56 , \us12/n55 , \us12/n54 , \us12/n53 , \us12/n52 ,
         \us12/n51 , \us12/n50 , \us12/n49 , \us12/n48 , \us12/n47 ,
         \us12/n46 , \us12/n45 , \us12/n44 , \us12/n43 , \us12/n42 ,
         \us12/n41 , \us12/n40 , \us12/n39 , \us12/n38 , \us12/n37 ,
         \us12/n36 , \us12/n35 , \us12/n34 , \us12/n33 , \us12/n32 ,
         \us12/n31 , \us12/n30 , \us12/n29 , \us12/n28 , \us12/n27 ,
         \us12/n26 , \us12/n25 , \us12/n24 , \us12/n23 , \us12/n22 ,
         \us12/n21 , \us12/n20 , \us12/n19 , \us12/n18 , \us12/n17 ,
         \us12/n16 , \us12/n15 , \us12/n14 , \us12/n13 , \us12/n12 ,
         \us12/n11 , \us12/n10 , \us12/n9 , \us12/n8 , \us12/n7 , \us12/n6 ,
         \us12/n5 , \us12/n4 , \us12/n3 , \us12/n2 , \us12/n1 , \us13/n358 ,
         \us13/n357 , \us13/n356 , \us13/n355 , \us13/n354 , \us13/n353 ,
         \us13/n352 , \us13/n351 , \us13/n350 , \us13/n349 , \us13/n348 ,
         \us13/n347 , \us13/n346 , \us13/n345 , \us13/n344 , \us13/n343 ,
         \us13/n342 , \us13/n341 , \us13/n340 , \us13/n339 , \us13/n338 ,
         \us13/n337 , \us13/n336 , \us13/n335 , \us13/n334 , \us13/n333 ,
         \us13/n332 , \us13/n331 , \us13/n330 , \us13/n329 , \us13/n328 ,
         \us13/n327 , \us13/n326 , \us13/n325 , \us13/n324 , \us13/n323 ,
         \us13/n322 , \us13/n321 , \us13/n320 , \us13/n319 , \us13/n318 ,
         \us13/n317 , \us13/n316 , \us13/n315 , \us13/n314 , \us13/n313 ,
         \us13/n312 , \us13/n311 , \us13/n310 , \us13/n309 , \us13/n308 ,
         \us13/n307 , \us13/n306 , \us13/n305 , \us13/n304 , \us13/n303 ,
         \us13/n302 , \us13/n301 , \us13/n300 , \us13/n299 , \us13/n298 ,
         \us13/n297 , \us13/n296 , \us13/n295 , \us13/n294 , \us13/n293 ,
         \us13/n292 , \us13/n291 , \us13/n290 , \us13/n289 , \us13/n288 ,
         \us13/n287 , \us13/n286 , \us13/n285 , \us13/n284 , \us13/n283 ,
         \us13/n282 , \us13/n281 , \us13/n280 , \us13/n279 , \us13/n278 ,
         \us13/n277 , \us13/n276 , \us13/n275 , \us13/n274 , \us13/n273 ,
         \us13/n272 , \us13/n271 , \us13/n270 , \us13/n269 , \us13/n268 ,
         \us13/n267 , \us13/n266 , \us13/n265 , \us13/n264 , \us13/n263 ,
         \us13/n262 , \us13/n261 , \us13/n260 , \us13/n259 , \us13/n258 ,
         \us13/n257 , \us13/n256 , \us13/n255 , \us13/n254 , \us13/n253 ,
         \us13/n252 , \us13/n251 , \us13/n250 , \us13/n249 , \us13/n248 ,
         \us13/n247 , \us13/n246 , \us13/n245 , \us13/n244 , \us13/n243 ,
         \us13/n242 , \us13/n241 , \us13/n240 , \us13/n239 , \us13/n238 ,
         \us13/n237 , \us13/n236 , \us13/n235 , \us13/n234 , \us13/n233 ,
         \us13/n232 , \us13/n231 , \us13/n230 , \us13/n229 , \us13/n228 ,
         \us13/n227 , \us13/n226 , \us13/n225 , \us13/n224 , \us13/n223 ,
         \us13/n222 , \us13/n221 , \us13/n220 , \us13/n219 , \us13/n218 ,
         \us13/n217 , \us13/n216 , \us13/n215 , \us13/n214 , \us13/n213 ,
         \us13/n212 , \us13/n211 , \us13/n210 , \us13/n209 , \us13/n208 ,
         \us13/n207 , \us13/n206 , \us13/n205 , \us13/n204 , \us13/n203 ,
         \us13/n202 , \us13/n201 , \us13/n200 , \us13/n199 , \us13/n198 ,
         \us13/n197 , \us13/n196 , \us13/n195 , \us13/n194 , \us13/n193 ,
         \us13/n192 , \us13/n191 , \us13/n190 , \us13/n189 , \us13/n188 ,
         \us13/n187 , \us13/n186 , \us13/n185 , \us13/n184 , \us13/n183 ,
         \us13/n182 , \us13/n181 , \us13/n180 , \us13/n179 , \us13/n178 ,
         \us13/n177 , \us13/n176 , \us13/n175 , \us13/n174 , \us13/n173 ,
         \us13/n172 , \us13/n171 , \us13/n170 , \us13/n169 , \us13/n168 ,
         \us13/n167 , \us13/n166 , \us13/n165 , \us13/n164 , \us13/n163 ,
         \us13/n162 , \us13/n161 , \us13/n160 , \us13/n159 , \us13/n158 ,
         \us13/n157 , \us13/n156 , \us13/n155 , \us13/n154 , \us13/n153 ,
         \us13/n152 , \us13/n151 , \us13/n150 , \us13/n149 , \us13/n148 ,
         \us13/n147 , \us13/n146 , \us13/n145 , \us13/n144 , \us13/n143 ,
         \us13/n142 , \us13/n141 , \us13/n140 , \us13/n139 , \us13/n138 ,
         \us13/n137 , \us13/n136 , \us13/n135 , \us13/n134 , \us13/n133 ,
         \us13/n132 , \us13/n131 , \us13/n130 , \us13/n129 , \us13/n128 ,
         \us13/n127 , \us13/n126 , \us13/n125 , \us13/n124 , \us13/n123 ,
         \us13/n122 , \us13/n121 , \us13/n120 , \us13/n119 , \us13/n118 ,
         \us13/n117 , \us13/n116 , \us13/n115 , \us13/n114 , \us13/n113 ,
         \us13/n112 , \us13/n111 , \us13/n110 , \us13/n109 , \us13/n108 ,
         \us13/n107 , \us13/n106 , \us13/n105 , \us13/n104 , \us13/n103 ,
         \us13/n102 , \us13/n101 , \us13/n100 , \us13/n99 , \us13/n98 ,
         \us13/n97 , \us13/n96 , \us13/n95 , \us13/n94 , \us13/n93 ,
         \us13/n92 , \us13/n91 , \us13/n90 , \us13/n89 , \us13/n88 ,
         \us13/n87 , \us13/n86 , \us13/n85 , \us13/n84 , \us13/n83 ,
         \us13/n82 , \us13/n81 , \us13/n80 , \us13/n79 , \us13/n78 ,
         \us13/n77 , \us13/n76 , \us13/n75 , \us13/n74 , \us13/n73 ,
         \us13/n72 , \us13/n71 , \us13/n70 , \us13/n69 , \us13/n68 ,
         \us13/n67 , \us13/n66 , \us13/n65 , \us13/n64 , \us13/n63 ,
         \us13/n62 , \us13/n61 , \us13/n60 , \us13/n59 , \us13/n58 ,
         \us13/n57 , \us13/n56 , \us13/n55 , \us13/n54 , \us13/n53 ,
         \us13/n52 , \us13/n51 , \us13/n50 , \us13/n49 , \us13/n48 ,
         \us13/n47 , \us13/n46 , \us13/n45 , \us13/n44 , \us13/n43 ,
         \us13/n42 , \us13/n41 , \us13/n40 , \us13/n39 , \us13/n38 ,
         \us13/n37 , \us13/n36 , \us13/n35 , \us13/n34 , \us13/n33 ,
         \us13/n32 , \us13/n31 , \us13/n30 , \us13/n29 , \us13/n28 ,
         \us13/n27 , \us13/n26 , \us13/n25 , \us13/n24 , \us13/n23 ,
         \us13/n22 , \us13/n21 , \us13/n20 , \us13/n19 , \us13/n18 ,
         \us13/n17 , \us13/n16 , \us13/n15 , \us13/n14 , \us13/n13 ,
         \us13/n12 , \us13/n11 , \us13/n10 , \us13/n9 , \us13/n8 , \us13/n7 ,
         \us13/n6 , \us13/n5 , \us13/n4 , \us13/n3 , \us13/n2 , \us13/n1 ,
         \us20/n358 , \us20/n357 , \us20/n356 , \us20/n355 , \us20/n354 ,
         \us20/n353 , \us20/n352 , \us20/n351 , \us20/n350 , \us20/n349 ,
         \us20/n348 , \us20/n347 , \us20/n346 , \us20/n345 , \us20/n344 ,
         \us20/n343 , \us20/n342 , \us20/n341 , \us20/n340 , \us20/n339 ,
         \us20/n338 , \us20/n337 , \us20/n336 , \us20/n335 , \us20/n334 ,
         \us20/n333 , \us20/n332 , \us20/n331 , \us20/n330 , \us20/n329 ,
         \us20/n328 , \us20/n327 , \us20/n326 , \us20/n325 , \us20/n324 ,
         \us20/n323 , \us20/n322 , \us20/n321 , \us20/n320 , \us20/n319 ,
         \us20/n318 , \us20/n317 , \us20/n316 , \us20/n315 , \us20/n314 ,
         \us20/n313 , \us20/n312 , \us20/n311 , \us20/n310 , \us20/n309 ,
         \us20/n308 , \us20/n307 , \us20/n306 , \us20/n305 , \us20/n304 ,
         \us20/n303 , \us20/n302 , \us20/n301 , \us20/n300 , \us20/n299 ,
         \us20/n298 , \us20/n297 , \us20/n296 , \us20/n295 , \us20/n294 ,
         \us20/n293 , \us20/n292 , \us20/n291 , \us20/n290 , \us20/n289 ,
         \us20/n288 , \us20/n287 , \us20/n286 , \us20/n285 , \us20/n284 ,
         \us20/n283 , \us20/n282 , \us20/n281 , \us20/n280 , \us20/n279 ,
         \us20/n278 , \us20/n277 , \us20/n276 , \us20/n275 , \us20/n274 ,
         \us20/n273 , \us20/n272 , \us20/n271 , \us20/n270 , \us20/n269 ,
         \us20/n268 , \us20/n267 , \us20/n266 , \us20/n265 , \us20/n264 ,
         \us20/n263 , \us20/n262 , \us20/n261 , \us20/n260 , \us20/n259 ,
         \us20/n258 , \us20/n257 , \us20/n256 , \us20/n255 , \us20/n254 ,
         \us20/n253 , \us20/n252 , \us20/n251 , \us20/n250 , \us20/n249 ,
         \us20/n248 , \us20/n247 , \us20/n246 , \us20/n245 , \us20/n244 ,
         \us20/n243 , \us20/n242 , \us20/n241 , \us20/n240 , \us20/n239 ,
         \us20/n238 , \us20/n237 , \us20/n236 , \us20/n235 , \us20/n234 ,
         \us20/n233 , \us20/n232 , \us20/n231 , \us20/n230 , \us20/n229 ,
         \us20/n228 , \us20/n227 , \us20/n226 , \us20/n225 , \us20/n224 ,
         \us20/n223 , \us20/n222 , \us20/n221 , \us20/n220 , \us20/n219 ,
         \us20/n218 , \us20/n217 , \us20/n216 , \us20/n215 , \us20/n214 ,
         \us20/n213 , \us20/n212 , \us20/n211 , \us20/n210 , \us20/n209 ,
         \us20/n208 , \us20/n207 , \us20/n206 , \us20/n205 , \us20/n204 ,
         \us20/n203 , \us20/n202 , \us20/n201 , \us20/n200 , \us20/n199 ,
         \us20/n198 , \us20/n197 , \us20/n196 , \us20/n195 , \us20/n194 ,
         \us20/n193 , \us20/n192 , \us20/n191 , \us20/n190 , \us20/n189 ,
         \us20/n188 , \us20/n187 , \us20/n186 , \us20/n185 , \us20/n184 ,
         \us20/n183 , \us20/n182 , \us20/n181 , \us20/n180 , \us20/n179 ,
         \us20/n178 , \us20/n177 , \us20/n176 , \us20/n175 , \us20/n174 ,
         \us20/n173 , \us20/n172 , \us20/n171 , \us20/n170 , \us20/n169 ,
         \us20/n168 , \us20/n167 , \us20/n166 , \us20/n165 , \us20/n164 ,
         \us20/n163 , \us20/n162 , \us20/n161 , \us20/n160 , \us20/n159 ,
         \us20/n158 , \us20/n157 , \us20/n156 , \us20/n155 , \us20/n154 ,
         \us20/n153 , \us20/n152 , \us20/n151 , \us20/n150 , \us20/n149 ,
         \us20/n148 , \us20/n147 , \us20/n146 , \us20/n145 , \us20/n144 ,
         \us20/n143 , \us20/n142 , \us20/n141 , \us20/n140 , \us20/n139 ,
         \us20/n138 , \us20/n137 , \us20/n136 , \us20/n135 , \us20/n134 ,
         \us20/n133 , \us20/n132 , \us20/n131 , \us20/n130 , \us20/n129 ,
         \us20/n128 , \us20/n127 , \us20/n126 , \us20/n125 , \us20/n124 ,
         \us20/n123 , \us20/n122 , \us20/n121 , \us20/n120 , \us20/n119 ,
         \us20/n118 , \us20/n117 , \us20/n116 , \us20/n115 , \us20/n114 ,
         \us20/n113 , \us20/n112 , \us20/n111 , \us20/n110 , \us20/n109 ,
         \us20/n108 , \us20/n107 , \us20/n106 , \us20/n105 , \us20/n104 ,
         \us20/n103 , \us20/n102 , \us20/n101 , \us20/n100 , \us20/n99 ,
         \us20/n98 , \us20/n97 , \us20/n96 , \us20/n95 , \us20/n94 ,
         \us20/n93 , \us20/n92 , \us20/n91 , \us20/n90 , \us20/n89 ,
         \us20/n88 , \us20/n87 , \us20/n86 , \us20/n85 , \us20/n84 ,
         \us20/n83 , \us20/n82 , \us20/n81 , \us20/n80 , \us20/n79 ,
         \us20/n78 , \us20/n77 , \us20/n76 , \us20/n75 , \us20/n74 ,
         \us20/n73 , \us20/n72 , \us20/n71 , \us20/n70 , \us20/n69 ,
         \us20/n68 , \us20/n67 , \us20/n66 , \us20/n65 , \us20/n64 ,
         \us20/n63 , \us20/n62 , \us20/n61 , \us20/n60 , \us20/n59 ,
         \us20/n58 , \us20/n57 , \us20/n56 , \us20/n55 , \us20/n54 ,
         \us20/n53 , \us20/n52 , \us20/n51 , \us20/n50 , \us20/n49 ,
         \us20/n48 , \us20/n47 , \us20/n46 , \us20/n45 , \us20/n44 ,
         \us20/n43 , \us20/n42 , \us20/n41 , \us20/n40 , \us20/n39 ,
         \us20/n38 , \us20/n37 , \us20/n36 , \us20/n35 , \us20/n34 ,
         \us20/n33 , \us20/n32 , \us20/n31 , \us20/n30 , \us20/n29 ,
         \us20/n28 , \us20/n27 , \us20/n26 , \us20/n25 , \us20/n24 ,
         \us20/n23 , \us20/n22 , \us20/n21 , \us20/n20 , \us20/n19 ,
         \us20/n18 , \us20/n17 , \us20/n16 , \us20/n15 , \us20/n14 ,
         \us20/n13 , \us20/n12 , \us20/n11 , \us20/n10 , \us20/n9 , \us20/n8 ,
         \us20/n7 , \us20/n6 , \us20/n5 , \us20/n4 , \us20/n3 , \us20/n2 ,
         \us20/n1 , \us21/n358 , \us21/n357 , \us21/n356 , \us21/n355 ,
         \us21/n354 , \us21/n353 , \us21/n352 , \us21/n351 , \us21/n350 ,
         \us21/n349 , \us21/n348 , \us21/n347 , \us21/n346 , \us21/n345 ,
         \us21/n344 , \us21/n343 , \us21/n342 , \us21/n341 , \us21/n340 ,
         \us21/n339 , \us21/n338 , \us21/n337 , \us21/n336 , \us21/n335 ,
         \us21/n334 , \us21/n333 , \us21/n332 , \us21/n331 , \us21/n330 ,
         \us21/n329 , \us21/n328 , \us21/n327 , \us21/n326 , \us21/n325 ,
         \us21/n324 , \us21/n323 , \us21/n322 , \us21/n321 , \us21/n320 ,
         \us21/n319 , \us21/n318 , \us21/n317 , \us21/n316 , \us21/n315 ,
         \us21/n314 , \us21/n313 , \us21/n312 , \us21/n311 , \us21/n310 ,
         \us21/n309 , \us21/n308 , \us21/n307 , \us21/n306 , \us21/n305 ,
         \us21/n304 , \us21/n303 , \us21/n302 , \us21/n301 , \us21/n300 ,
         \us21/n299 , \us21/n298 , \us21/n297 , \us21/n296 , \us21/n295 ,
         \us21/n294 , \us21/n293 , \us21/n292 , \us21/n291 , \us21/n290 ,
         \us21/n289 , \us21/n288 , \us21/n287 , \us21/n286 , \us21/n285 ,
         \us21/n284 , \us21/n283 , \us21/n282 , \us21/n281 , \us21/n280 ,
         \us21/n279 , \us21/n278 , \us21/n277 , \us21/n276 , \us21/n275 ,
         \us21/n274 , \us21/n273 , \us21/n272 , \us21/n271 , \us21/n270 ,
         \us21/n269 , \us21/n268 , \us21/n267 , \us21/n266 , \us21/n265 ,
         \us21/n264 , \us21/n263 , \us21/n262 , \us21/n261 , \us21/n260 ,
         \us21/n259 , \us21/n258 , \us21/n257 , \us21/n256 , \us21/n255 ,
         \us21/n254 , \us21/n253 , \us21/n252 , \us21/n251 , \us21/n250 ,
         \us21/n249 , \us21/n248 , \us21/n247 , \us21/n246 , \us21/n245 ,
         \us21/n244 , \us21/n243 , \us21/n242 , \us21/n241 , \us21/n240 ,
         \us21/n239 , \us21/n238 , \us21/n237 , \us21/n236 , \us21/n235 ,
         \us21/n234 , \us21/n233 , \us21/n232 , \us21/n231 , \us21/n230 ,
         \us21/n229 , \us21/n228 , \us21/n227 , \us21/n226 , \us21/n225 ,
         \us21/n224 , \us21/n223 , \us21/n222 , \us21/n221 , \us21/n220 ,
         \us21/n219 , \us21/n218 , \us21/n217 , \us21/n216 , \us21/n215 ,
         \us21/n214 , \us21/n213 , \us21/n212 , \us21/n211 , \us21/n210 ,
         \us21/n209 , \us21/n208 , \us21/n207 , \us21/n206 , \us21/n205 ,
         \us21/n204 , \us21/n203 , \us21/n202 , \us21/n201 , \us21/n200 ,
         \us21/n199 , \us21/n198 , \us21/n197 , \us21/n196 , \us21/n195 ,
         \us21/n194 , \us21/n193 , \us21/n192 , \us21/n191 , \us21/n190 ,
         \us21/n189 , \us21/n188 , \us21/n187 , \us21/n186 , \us21/n185 ,
         \us21/n184 , \us21/n183 , \us21/n182 , \us21/n181 , \us21/n180 ,
         \us21/n179 , \us21/n178 , \us21/n177 , \us21/n176 , \us21/n175 ,
         \us21/n174 , \us21/n173 , \us21/n172 , \us21/n171 , \us21/n170 ,
         \us21/n169 , \us21/n168 , \us21/n167 , \us21/n166 , \us21/n165 ,
         \us21/n164 , \us21/n163 , \us21/n162 , \us21/n161 , \us21/n160 ,
         \us21/n159 , \us21/n158 , \us21/n157 , \us21/n156 , \us21/n155 ,
         \us21/n154 , \us21/n153 , \us21/n152 , \us21/n151 , \us21/n150 ,
         \us21/n149 , \us21/n148 , \us21/n147 , \us21/n146 , \us21/n145 ,
         \us21/n144 , \us21/n143 , \us21/n142 , \us21/n141 , \us21/n140 ,
         \us21/n139 , \us21/n138 , \us21/n137 , \us21/n136 , \us21/n135 ,
         \us21/n134 , \us21/n133 , \us21/n132 , \us21/n131 , \us21/n130 ,
         \us21/n129 , \us21/n128 , \us21/n127 , \us21/n126 , \us21/n125 ,
         \us21/n124 , \us21/n123 , \us21/n122 , \us21/n121 , \us21/n120 ,
         \us21/n119 , \us21/n118 , \us21/n117 , \us21/n116 , \us21/n115 ,
         \us21/n114 , \us21/n113 , \us21/n112 , \us21/n111 , \us21/n110 ,
         \us21/n109 , \us21/n108 , \us21/n107 , \us21/n106 , \us21/n105 ,
         \us21/n104 , \us21/n103 , \us21/n102 , \us21/n101 , \us21/n100 ,
         \us21/n99 , \us21/n98 , \us21/n97 , \us21/n96 , \us21/n95 ,
         \us21/n94 , \us21/n93 , \us21/n92 , \us21/n91 , \us21/n90 ,
         \us21/n89 , \us21/n88 , \us21/n87 , \us21/n86 , \us21/n85 ,
         \us21/n84 , \us21/n83 , \us21/n82 , \us21/n81 , \us21/n80 ,
         \us21/n79 , \us21/n78 , \us21/n77 , \us21/n76 , \us21/n75 ,
         \us21/n74 , \us21/n73 , \us21/n72 , \us21/n71 , \us21/n70 ,
         \us21/n69 , \us21/n68 , \us21/n67 , \us21/n66 , \us21/n65 ,
         \us21/n64 , \us21/n63 , \us21/n62 , \us21/n61 , \us21/n60 ,
         \us21/n59 , \us21/n58 , \us21/n57 , \us21/n56 , \us21/n55 ,
         \us21/n54 , \us21/n53 , \us21/n52 , \us21/n51 , \us21/n50 ,
         \us21/n49 , \us21/n48 , \us21/n47 , \us21/n46 , \us21/n45 ,
         \us21/n44 , \us21/n43 , \us21/n42 , \us21/n41 , \us21/n40 ,
         \us21/n39 , \us21/n38 , \us21/n37 , \us21/n36 , \us21/n35 ,
         \us21/n34 , \us21/n33 , \us21/n32 , \us21/n31 , \us21/n30 ,
         \us21/n29 , \us21/n28 , \us21/n27 , \us21/n26 , \us21/n25 ,
         \us21/n24 , \us21/n23 , \us21/n22 , \us21/n21 , \us21/n20 ,
         \us21/n19 , \us21/n18 , \us21/n17 , \us21/n16 , \us21/n15 ,
         \us21/n14 , \us21/n13 , \us21/n12 , \us21/n11 , \us21/n10 , \us21/n9 ,
         \us21/n8 , \us21/n7 , \us21/n6 , \us21/n5 , \us21/n4 , \us21/n3 ,
         \us21/n2 , \us21/n1 , \us22/n358 , \us22/n357 , \us22/n356 ,
         \us22/n355 , \us22/n354 , \us22/n353 , \us22/n352 , \us22/n351 ,
         \us22/n350 , \us22/n349 , \us22/n348 , \us22/n347 , \us22/n346 ,
         \us22/n345 , \us22/n344 , \us22/n343 , \us22/n342 , \us22/n341 ,
         \us22/n340 , \us22/n339 , \us22/n338 , \us22/n337 , \us22/n336 ,
         \us22/n335 , \us22/n334 , \us22/n333 , \us22/n332 , \us22/n331 ,
         \us22/n330 , \us22/n329 , \us22/n328 , \us22/n327 , \us22/n326 ,
         \us22/n325 , \us22/n324 , \us22/n323 , \us22/n322 , \us22/n321 ,
         \us22/n320 , \us22/n319 , \us22/n318 , \us22/n317 , \us22/n316 ,
         \us22/n315 , \us22/n314 , \us22/n313 , \us22/n312 , \us22/n311 ,
         \us22/n310 , \us22/n309 , \us22/n308 , \us22/n307 , \us22/n306 ,
         \us22/n305 , \us22/n304 , \us22/n303 , \us22/n302 , \us22/n301 ,
         \us22/n300 , \us22/n299 , \us22/n298 , \us22/n297 , \us22/n296 ,
         \us22/n295 , \us22/n294 , \us22/n293 , \us22/n292 , \us22/n291 ,
         \us22/n290 , \us22/n289 , \us22/n288 , \us22/n287 , \us22/n286 ,
         \us22/n285 , \us22/n284 , \us22/n283 , \us22/n282 , \us22/n281 ,
         \us22/n280 , \us22/n279 , \us22/n278 , \us22/n277 , \us22/n276 ,
         \us22/n275 , \us22/n274 , \us22/n273 , \us22/n272 , \us22/n271 ,
         \us22/n270 , \us22/n269 , \us22/n268 , \us22/n267 , \us22/n266 ,
         \us22/n265 , \us22/n264 , \us22/n263 , \us22/n262 , \us22/n261 ,
         \us22/n260 , \us22/n259 , \us22/n258 , \us22/n257 , \us22/n256 ,
         \us22/n255 , \us22/n254 , \us22/n253 , \us22/n252 , \us22/n251 ,
         \us22/n250 , \us22/n249 , \us22/n248 , \us22/n247 , \us22/n246 ,
         \us22/n245 , \us22/n244 , \us22/n243 , \us22/n242 , \us22/n241 ,
         \us22/n240 , \us22/n239 , \us22/n238 , \us22/n237 , \us22/n236 ,
         \us22/n235 , \us22/n234 , \us22/n233 , \us22/n232 , \us22/n231 ,
         \us22/n230 , \us22/n229 , \us22/n228 , \us22/n227 , \us22/n226 ,
         \us22/n225 , \us22/n224 , \us22/n223 , \us22/n222 , \us22/n221 ,
         \us22/n220 , \us22/n219 , \us22/n218 , \us22/n217 , \us22/n216 ,
         \us22/n215 , \us22/n214 , \us22/n213 , \us22/n212 , \us22/n211 ,
         \us22/n210 , \us22/n209 , \us22/n208 , \us22/n207 , \us22/n206 ,
         \us22/n205 , \us22/n204 , \us22/n203 , \us22/n202 , \us22/n201 ,
         \us22/n200 , \us22/n199 , \us22/n198 , \us22/n197 , \us22/n196 ,
         \us22/n195 , \us22/n194 , \us22/n193 , \us22/n192 , \us22/n191 ,
         \us22/n190 , \us22/n189 , \us22/n188 , \us22/n187 , \us22/n186 ,
         \us22/n185 , \us22/n184 , \us22/n183 , \us22/n182 , \us22/n181 ,
         \us22/n180 , \us22/n179 , \us22/n178 , \us22/n177 , \us22/n176 ,
         \us22/n175 , \us22/n174 , \us22/n173 , \us22/n172 , \us22/n171 ,
         \us22/n170 , \us22/n169 , \us22/n168 , \us22/n167 , \us22/n166 ,
         \us22/n165 , \us22/n164 , \us22/n163 , \us22/n162 , \us22/n161 ,
         \us22/n160 , \us22/n159 , \us22/n158 , \us22/n157 , \us22/n156 ,
         \us22/n155 , \us22/n154 , \us22/n153 , \us22/n152 , \us22/n151 ,
         \us22/n150 , \us22/n149 , \us22/n148 , \us22/n147 , \us22/n146 ,
         \us22/n145 , \us22/n144 , \us22/n143 , \us22/n142 , \us22/n141 ,
         \us22/n140 , \us22/n139 , \us22/n138 , \us22/n137 , \us22/n136 ,
         \us22/n135 , \us22/n134 , \us22/n133 , \us22/n132 , \us22/n131 ,
         \us22/n130 , \us22/n129 , \us22/n128 , \us22/n127 , \us22/n126 ,
         \us22/n125 , \us22/n124 , \us22/n123 , \us22/n122 , \us22/n121 ,
         \us22/n120 , \us22/n119 , \us22/n118 , \us22/n117 , \us22/n116 ,
         \us22/n115 , \us22/n114 , \us22/n113 , \us22/n112 , \us22/n111 ,
         \us22/n110 , \us22/n109 , \us22/n108 , \us22/n107 , \us22/n106 ,
         \us22/n105 , \us22/n104 , \us22/n103 , \us22/n102 , \us22/n101 ,
         \us22/n100 , \us22/n99 , \us22/n98 , \us22/n97 , \us22/n96 ,
         \us22/n95 , \us22/n94 , \us22/n93 , \us22/n92 , \us22/n91 ,
         \us22/n90 , \us22/n89 , \us22/n88 , \us22/n87 , \us22/n86 ,
         \us22/n85 , \us22/n84 , \us22/n83 , \us22/n82 , \us22/n81 ,
         \us22/n80 , \us22/n79 , \us22/n78 , \us22/n77 , \us22/n76 ,
         \us22/n75 , \us22/n74 , \us22/n73 , \us22/n72 , \us22/n71 ,
         \us22/n70 , \us22/n69 , \us22/n68 , \us22/n67 , \us22/n66 ,
         \us22/n65 , \us22/n64 , \us22/n63 , \us22/n62 , \us22/n61 ,
         \us22/n60 , \us22/n59 , \us22/n58 , \us22/n57 , \us22/n56 ,
         \us22/n55 , \us22/n54 , \us22/n53 , \us22/n52 , \us22/n51 ,
         \us22/n50 , \us22/n49 , \us22/n48 , \us22/n47 , \us22/n46 ,
         \us22/n45 , \us22/n44 , \us22/n43 , \us22/n42 , \us22/n41 ,
         \us22/n40 , \us22/n39 , \us22/n38 , \us22/n37 , \us22/n36 ,
         \us22/n35 , \us22/n34 , \us22/n33 , \us22/n32 , \us22/n31 ,
         \us22/n30 , \us22/n29 , \us22/n28 , \us22/n27 , \us22/n26 ,
         \us22/n25 , \us22/n24 , \us22/n23 , \us22/n22 , \us22/n21 ,
         \us22/n20 , \us22/n19 , \us22/n18 , \us22/n17 , \us22/n16 ,
         \us22/n15 , \us22/n14 , \us22/n13 , \us22/n12 , \us22/n11 ,
         \us22/n10 , \us22/n9 , \us22/n8 , \us22/n7 , \us22/n6 , \us22/n5 ,
         \us22/n4 , \us22/n3 , \us22/n2 , \us22/n1 , \us23/n358 , \us23/n357 ,
         \us23/n356 , \us23/n355 , \us23/n354 , \us23/n353 , \us23/n352 ,
         \us23/n351 , \us23/n350 , \us23/n349 , \us23/n348 , \us23/n347 ,
         \us23/n346 , \us23/n345 , \us23/n344 , \us23/n343 , \us23/n342 ,
         \us23/n341 , \us23/n340 , \us23/n339 , \us23/n338 , \us23/n337 ,
         \us23/n336 , \us23/n335 , \us23/n334 , \us23/n333 , \us23/n332 ,
         \us23/n331 , \us23/n330 , \us23/n329 , \us23/n328 , \us23/n327 ,
         \us23/n326 , \us23/n325 , \us23/n324 , \us23/n323 , \us23/n322 ,
         \us23/n321 , \us23/n320 , \us23/n319 , \us23/n318 , \us23/n317 ,
         \us23/n316 , \us23/n315 , \us23/n314 , \us23/n313 , \us23/n312 ,
         \us23/n311 , \us23/n310 , \us23/n309 , \us23/n308 , \us23/n307 ,
         \us23/n306 , \us23/n305 , \us23/n304 , \us23/n303 , \us23/n302 ,
         \us23/n301 , \us23/n300 , \us23/n299 , \us23/n298 , \us23/n297 ,
         \us23/n296 , \us23/n295 , \us23/n294 , \us23/n293 , \us23/n292 ,
         \us23/n291 , \us23/n290 , \us23/n289 , \us23/n288 , \us23/n287 ,
         \us23/n286 , \us23/n285 , \us23/n284 , \us23/n283 , \us23/n282 ,
         \us23/n281 , \us23/n280 , \us23/n279 , \us23/n278 , \us23/n277 ,
         \us23/n276 , \us23/n275 , \us23/n274 , \us23/n273 , \us23/n272 ,
         \us23/n271 , \us23/n270 , \us23/n269 , \us23/n268 , \us23/n267 ,
         \us23/n266 , \us23/n265 , \us23/n264 , \us23/n263 , \us23/n262 ,
         \us23/n261 , \us23/n260 , \us23/n259 , \us23/n258 , \us23/n257 ,
         \us23/n256 , \us23/n255 , \us23/n254 , \us23/n253 , \us23/n252 ,
         \us23/n251 , \us23/n250 , \us23/n249 , \us23/n248 , \us23/n247 ,
         \us23/n246 , \us23/n245 , \us23/n244 , \us23/n243 , \us23/n242 ,
         \us23/n241 , \us23/n240 , \us23/n239 , \us23/n238 , \us23/n237 ,
         \us23/n236 , \us23/n235 , \us23/n234 , \us23/n233 , \us23/n232 ,
         \us23/n231 , \us23/n230 , \us23/n229 , \us23/n228 , \us23/n227 ,
         \us23/n226 , \us23/n225 , \us23/n224 , \us23/n223 , \us23/n222 ,
         \us23/n221 , \us23/n220 , \us23/n219 , \us23/n218 , \us23/n217 ,
         \us23/n216 , \us23/n215 , \us23/n214 , \us23/n213 , \us23/n212 ,
         \us23/n211 , \us23/n210 , \us23/n209 , \us23/n208 , \us23/n207 ,
         \us23/n206 , \us23/n205 , \us23/n204 , \us23/n203 , \us23/n202 ,
         \us23/n201 , \us23/n200 , \us23/n199 , \us23/n198 , \us23/n197 ,
         \us23/n196 , \us23/n195 , \us23/n194 , \us23/n193 , \us23/n192 ,
         \us23/n191 , \us23/n190 , \us23/n189 , \us23/n188 , \us23/n187 ,
         \us23/n186 , \us23/n185 , \us23/n184 , \us23/n183 , \us23/n182 ,
         \us23/n181 , \us23/n180 , \us23/n179 , \us23/n178 , \us23/n177 ,
         \us23/n176 , \us23/n175 , \us23/n174 , \us23/n173 , \us23/n172 ,
         \us23/n171 , \us23/n170 , \us23/n169 , \us23/n168 , \us23/n167 ,
         \us23/n166 , \us23/n165 , \us23/n164 , \us23/n163 , \us23/n162 ,
         \us23/n161 , \us23/n160 , \us23/n159 , \us23/n158 , \us23/n157 ,
         \us23/n156 , \us23/n155 , \us23/n154 , \us23/n153 , \us23/n152 ,
         \us23/n151 , \us23/n150 , \us23/n149 , \us23/n148 , \us23/n147 ,
         \us23/n146 , \us23/n145 , \us23/n144 , \us23/n143 , \us23/n142 ,
         \us23/n141 , \us23/n140 , \us23/n139 , \us23/n138 , \us23/n137 ,
         \us23/n136 , \us23/n135 , \us23/n134 , \us23/n133 , \us23/n132 ,
         \us23/n131 , \us23/n130 , \us23/n129 , \us23/n128 , \us23/n127 ,
         \us23/n126 , \us23/n125 , \us23/n124 , \us23/n123 , \us23/n122 ,
         \us23/n121 , \us23/n120 , \us23/n119 , \us23/n118 , \us23/n117 ,
         \us23/n116 , \us23/n115 , \us23/n114 , \us23/n113 , \us23/n112 ,
         \us23/n111 , \us23/n110 , \us23/n109 , \us23/n108 , \us23/n107 ,
         \us23/n106 , \us23/n105 , \us23/n104 , \us23/n103 , \us23/n102 ,
         \us23/n101 , \us23/n100 , \us23/n99 , \us23/n98 , \us23/n97 ,
         \us23/n96 , \us23/n95 , \us23/n94 , \us23/n93 , \us23/n92 ,
         \us23/n91 , \us23/n90 , \us23/n89 , \us23/n88 , \us23/n87 ,
         \us23/n86 , \us23/n85 , \us23/n84 , \us23/n83 , \us23/n82 ,
         \us23/n81 , \us23/n80 , \us23/n79 , \us23/n78 , \us23/n77 ,
         \us23/n76 , \us23/n75 , \us23/n74 , \us23/n73 , \us23/n72 ,
         \us23/n71 , \us23/n70 , \us23/n69 , \us23/n68 , \us23/n67 ,
         \us23/n66 , \us23/n65 , \us23/n64 , \us23/n63 , \us23/n62 ,
         \us23/n61 , \us23/n60 , \us23/n59 , \us23/n58 , \us23/n57 ,
         \us23/n56 , \us23/n55 , \us23/n54 , \us23/n53 , \us23/n52 ,
         \us23/n51 , \us23/n50 , \us23/n49 , \us23/n48 , \us23/n47 ,
         \us23/n46 , \us23/n45 , \us23/n44 , \us23/n43 , \us23/n42 ,
         \us23/n41 , \us23/n40 , \us23/n39 , \us23/n38 , \us23/n37 ,
         \us23/n36 , \us23/n35 , \us23/n34 , \us23/n33 , \us23/n32 ,
         \us23/n31 , \us23/n30 , \us23/n29 , \us23/n28 , \us23/n27 ,
         \us23/n26 , \us23/n25 , \us23/n24 , \us23/n23 , \us23/n22 ,
         \us23/n21 , \us23/n20 , \us23/n19 , \us23/n18 , \us23/n17 ,
         \us23/n16 , \us23/n15 , \us23/n14 , \us23/n13 , \us23/n12 ,
         \us23/n11 , \us23/n10 , \us23/n9 , \us23/n8 , \us23/n7 , \us23/n6 ,
         \us23/n5 , \us23/n4 , \us23/n3 , \us23/n2 , \us23/n1 , \us30/n358 ,
         \us30/n357 , \us30/n356 , \us30/n355 , \us30/n354 , \us30/n353 ,
         \us30/n352 , \us30/n351 , \us30/n350 , \us30/n349 , \us30/n348 ,
         \us30/n347 , \us30/n346 , \us30/n345 , \us30/n344 , \us30/n343 ,
         \us30/n342 , \us30/n341 , \us30/n340 , \us30/n339 , \us30/n338 ,
         \us30/n337 , \us30/n336 , \us30/n335 , \us30/n334 , \us30/n333 ,
         \us30/n332 , \us30/n331 , \us30/n330 , \us30/n329 , \us30/n328 ,
         \us30/n327 , \us30/n326 , \us30/n325 , \us30/n324 , \us30/n323 ,
         \us30/n322 , \us30/n321 , \us30/n320 , \us30/n319 , \us30/n318 ,
         \us30/n317 , \us30/n316 , \us30/n315 , \us30/n314 , \us30/n313 ,
         \us30/n312 , \us30/n311 , \us30/n310 , \us30/n309 , \us30/n308 ,
         \us30/n307 , \us30/n306 , \us30/n305 , \us30/n304 , \us30/n303 ,
         \us30/n302 , \us30/n301 , \us30/n300 , \us30/n299 , \us30/n298 ,
         \us30/n297 , \us30/n296 , \us30/n295 , \us30/n294 , \us30/n293 ,
         \us30/n292 , \us30/n291 , \us30/n290 , \us30/n289 , \us30/n288 ,
         \us30/n287 , \us30/n286 , \us30/n285 , \us30/n284 , \us30/n283 ,
         \us30/n282 , \us30/n281 , \us30/n280 , \us30/n279 , \us30/n278 ,
         \us30/n277 , \us30/n276 , \us30/n275 , \us30/n274 , \us30/n273 ,
         \us30/n272 , \us30/n271 , \us30/n270 , \us30/n269 , \us30/n268 ,
         \us30/n267 , \us30/n266 , \us30/n265 , \us30/n264 , \us30/n263 ,
         \us30/n262 , \us30/n261 , \us30/n260 , \us30/n259 , \us30/n258 ,
         \us30/n257 , \us30/n256 , \us30/n255 , \us30/n254 , \us30/n253 ,
         \us30/n252 , \us30/n251 , \us30/n250 , \us30/n249 , \us30/n248 ,
         \us30/n247 , \us30/n246 , \us30/n245 , \us30/n244 , \us30/n243 ,
         \us30/n242 , \us30/n241 , \us30/n240 , \us30/n239 , \us30/n238 ,
         \us30/n237 , \us30/n236 , \us30/n235 , \us30/n234 , \us30/n233 ,
         \us30/n232 , \us30/n231 , \us30/n230 , \us30/n229 , \us30/n228 ,
         \us30/n227 , \us30/n226 , \us30/n225 , \us30/n224 , \us30/n223 ,
         \us30/n222 , \us30/n221 , \us30/n220 , \us30/n219 , \us30/n218 ,
         \us30/n217 , \us30/n216 , \us30/n215 , \us30/n214 , \us30/n213 ,
         \us30/n212 , \us30/n211 , \us30/n210 , \us30/n209 , \us30/n208 ,
         \us30/n207 , \us30/n206 , \us30/n205 , \us30/n204 , \us30/n203 ,
         \us30/n202 , \us30/n201 , \us30/n200 , \us30/n199 , \us30/n198 ,
         \us30/n197 , \us30/n196 , \us30/n195 , \us30/n194 , \us30/n193 ,
         \us30/n192 , \us30/n191 , \us30/n190 , \us30/n189 , \us30/n188 ,
         \us30/n187 , \us30/n186 , \us30/n185 , \us30/n184 , \us30/n183 ,
         \us30/n182 , \us30/n181 , \us30/n180 , \us30/n179 , \us30/n178 ,
         \us30/n177 , \us30/n176 , \us30/n175 , \us30/n174 , \us30/n173 ,
         \us30/n172 , \us30/n171 , \us30/n170 , \us30/n169 , \us30/n168 ,
         \us30/n167 , \us30/n166 , \us30/n165 , \us30/n164 , \us30/n163 ,
         \us30/n162 , \us30/n161 , \us30/n160 , \us30/n159 , \us30/n158 ,
         \us30/n157 , \us30/n156 , \us30/n155 , \us30/n154 , \us30/n153 ,
         \us30/n152 , \us30/n151 , \us30/n150 , \us30/n149 , \us30/n148 ,
         \us30/n147 , \us30/n146 , \us30/n145 , \us30/n144 , \us30/n143 ,
         \us30/n142 , \us30/n141 , \us30/n140 , \us30/n139 , \us30/n138 ,
         \us30/n137 , \us30/n136 , \us30/n135 , \us30/n134 , \us30/n133 ,
         \us30/n132 , \us30/n131 , \us30/n130 , \us30/n129 , \us30/n128 ,
         \us30/n127 , \us30/n126 , \us30/n125 , \us30/n124 , \us30/n123 ,
         \us30/n122 , \us30/n121 , \us30/n120 , \us30/n119 , \us30/n118 ,
         \us30/n117 , \us30/n116 , \us30/n115 , \us30/n114 , \us30/n113 ,
         \us30/n112 , \us30/n111 , \us30/n110 , \us30/n109 , \us30/n108 ,
         \us30/n107 , \us30/n106 , \us30/n105 , \us30/n104 , \us30/n103 ,
         \us30/n102 , \us30/n101 , \us30/n100 , \us30/n99 , \us30/n98 ,
         \us30/n97 , \us30/n96 , \us30/n95 , \us30/n94 , \us30/n93 ,
         \us30/n92 , \us30/n91 , \us30/n90 , \us30/n89 , \us30/n88 ,
         \us30/n87 , \us30/n86 , \us30/n85 , \us30/n84 , \us30/n83 ,
         \us30/n82 , \us30/n81 , \us30/n80 , \us30/n79 , \us30/n78 ,
         \us30/n77 , \us30/n76 , \us30/n75 , \us30/n74 , \us30/n73 ,
         \us30/n72 , \us30/n71 , \us30/n70 , \us30/n69 , \us30/n68 ,
         \us30/n67 , \us30/n66 , \us30/n65 , \us30/n64 , \us30/n63 ,
         \us30/n62 , \us30/n61 , \us30/n60 , \us30/n59 , \us30/n58 ,
         \us30/n57 , \us30/n56 , \us30/n55 , \us30/n54 , \us30/n53 ,
         \us30/n52 , \us30/n51 , \us30/n50 , \us30/n49 , \us30/n48 ,
         \us30/n47 , \us30/n46 , \us30/n45 , \us30/n44 , \us30/n43 ,
         \us30/n42 , \us30/n41 , \us30/n40 , \us30/n39 , \us30/n38 ,
         \us30/n37 , \us30/n36 , \us30/n35 , \us30/n34 , \us30/n33 ,
         \us30/n32 , \us30/n31 , \us30/n30 , \us30/n29 , \us30/n28 ,
         \us30/n27 , \us30/n26 , \us30/n25 , \us30/n24 , \us30/n23 ,
         \us30/n22 , \us30/n21 , \us30/n20 , \us30/n19 , \us30/n18 ,
         \us30/n17 , \us30/n16 , \us30/n15 , \us30/n14 , \us30/n13 ,
         \us30/n12 , \us30/n11 , \us30/n10 , \us30/n9 , \us30/n8 , \us30/n7 ,
         \us30/n6 , \us30/n5 , \us30/n4 , \us30/n3 , \us30/n2 , \us30/n1 ,
         \us31/n358 , \us31/n357 , \us31/n356 , \us31/n355 , \us31/n354 ,
         \us31/n353 , \us31/n352 , \us31/n351 , \us31/n350 , \us31/n349 ,
         \us31/n348 , \us31/n347 , \us31/n346 , \us31/n345 , \us31/n344 ,
         \us31/n343 , \us31/n342 , \us31/n341 , \us31/n340 , \us31/n339 ,
         \us31/n338 , \us31/n337 , \us31/n336 , \us31/n335 , \us31/n334 ,
         \us31/n333 , \us31/n332 , \us31/n331 , \us31/n330 , \us31/n329 ,
         \us31/n328 , \us31/n327 , \us31/n326 , \us31/n325 , \us31/n324 ,
         \us31/n323 , \us31/n322 , \us31/n321 , \us31/n320 , \us31/n319 ,
         \us31/n318 , \us31/n317 , \us31/n316 , \us31/n315 , \us31/n314 ,
         \us31/n313 , \us31/n312 , \us31/n311 , \us31/n310 , \us31/n309 ,
         \us31/n308 , \us31/n307 , \us31/n306 , \us31/n305 , \us31/n304 ,
         \us31/n303 , \us31/n302 , \us31/n301 , \us31/n300 , \us31/n299 ,
         \us31/n298 , \us31/n297 , \us31/n296 , \us31/n295 , \us31/n294 ,
         \us31/n293 , \us31/n292 , \us31/n291 , \us31/n290 , \us31/n289 ,
         \us31/n288 , \us31/n287 , \us31/n286 , \us31/n285 , \us31/n284 ,
         \us31/n283 , \us31/n282 , \us31/n281 , \us31/n280 , \us31/n279 ,
         \us31/n278 , \us31/n277 , \us31/n276 , \us31/n275 , \us31/n274 ,
         \us31/n273 , \us31/n272 , \us31/n271 , \us31/n270 , \us31/n269 ,
         \us31/n268 , \us31/n267 , \us31/n266 , \us31/n265 , \us31/n264 ,
         \us31/n263 , \us31/n262 , \us31/n261 , \us31/n260 , \us31/n259 ,
         \us31/n258 , \us31/n257 , \us31/n256 , \us31/n255 , \us31/n254 ,
         \us31/n253 , \us31/n252 , \us31/n251 , \us31/n250 , \us31/n249 ,
         \us31/n248 , \us31/n247 , \us31/n246 , \us31/n245 , \us31/n244 ,
         \us31/n243 , \us31/n242 , \us31/n241 , \us31/n240 , \us31/n239 ,
         \us31/n238 , \us31/n237 , \us31/n236 , \us31/n235 , \us31/n234 ,
         \us31/n233 , \us31/n232 , \us31/n231 , \us31/n230 , \us31/n229 ,
         \us31/n228 , \us31/n227 , \us31/n226 , \us31/n225 , \us31/n224 ,
         \us31/n223 , \us31/n222 , \us31/n221 , \us31/n220 , \us31/n219 ,
         \us31/n218 , \us31/n217 , \us31/n216 , \us31/n215 , \us31/n214 ,
         \us31/n213 , \us31/n212 , \us31/n211 , \us31/n210 , \us31/n209 ,
         \us31/n208 , \us31/n207 , \us31/n206 , \us31/n205 , \us31/n204 ,
         \us31/n203 , \us31/n202 , \us31/n201 , \us31/n200 , \us31/n199 ,
         \us31/n198 , \us31/n197 , \us31/n196 , \us31/n195 , \us31/n194 ,
         \us31/n193 , \us31/n192 , \us31/n191 , \us31/n190 , \us31/n189 ,
         \us31/n188 , \us31/n187 , \us31/n186 , \us31/n185 , \us31/n184 ,
         \us31/n183 , \us31/n182 , \us31/n181 , \us31/n180 , \us31/n179 ,
         \us31/n178 , \us31/n177 , \us31/n176 , \us31/n175 , \us31/n174 ,
         \us31/n173 , \us31/n172 , \us31/n171 , \us31/n170 , \us31/n169 ,
         \us31/n168 , \us31/n167 , \us31/n166 , \us31/n165 , \us31/n164 ,
         \us31/n163 , \us31/n162 , \us31/n161 , \us31/n160 , \us31/n159 ,
         \us31/n158 , \us31/n157 , \us31/n156 , \us31/n155 , \us31/n154 ,
         \us31/n153 , \us31/n152 , \us31/n151 , \us31/n150 , \us31/n149 ,
         \us31/n148 , \us31/n147 , \us31/n146 , \us31/n145 , \us31/n144 ,
         \us31/n143 , \us31/n142 , \us31/n141 , \us31/n140 , \us31/n139 ,
         \us31/n138 , \us31/n137 , \us31/n136 , \us31/n135 , \us31/n134 ,
         \us31/n133 , \us31/n132 , \us31/n131 , \us31/n130 , \us31/n129 ,
         \us31/n128 , \us31/n127 , \us31/n126 , \us31/n125 , \us31/n124 ,
         \us31/n123 , \us31/n122 , \us31/n121 , \us31/n120 , \us31/n119 ,
         \us31/n118 , \us31/n117 , \us31/n116 , \us31/n115 , \us31/n114 ,
         \us31/n113 , \us31/n112 , \us31/n111 , \us31/n110 , \us31/n109 ,
         \us31/n108 , \us31/n107 , \us31/n106 , \us31/n105 , \us31/n104 ,
         \us31/n103 , \us31/n102 , \us31/n101 , \us31/n100 , \us31/n99 ,
         \us31/n98 , \us31/n97 , \us31/n96 , \us31/n95 , \us31/n94 ,
         \us31/n93 , \us31/n92 , \us31/n91 , \us31/n90 , \us31/n89 ,
         \us31/n88 , \us31/n87 , \us31/n86 , \us31/n85 , \us31/n84 ,
         \us31/n83 , \us31/n82 , \us31/n81 , \us31/n80 , \us31/n79 ,
         \us31/n78 , \us31/n77 , \us31/n76 , \us31/n75 , \us31/n74 ,
         \us31/n73 , \us31/n72 , \us31/n71 , \us31/n70 , \us31/n69 ,
         \us31/n68 , \us31/n67 , \us31/n66 , \us31/n65 , \us31/n64 ,
         \us31/n63 , \us31/n62 , \us31/n61 , \us31/n60 , \us31/n59 ,
         \us31/n58 , \us31/n57 , \us31/n56 , \us31/n55 , \us31/n54 ,
         \us31/n53 , \us31/n52 , \us31/n51 , \us31/n50 , \us31/n49 ,
         \us31/n48 , \us31/n47 , \us31/n46 , \us31/n45 , \us31/n44 ,
         \us31/n43 , \us31/n42 , \us31/n41 , \us31/n40 , \us31/n39 ,
         \us31/n38 , \us31/n37 , \us31/n36 , \us31/n35 , \us31/n34 ,
         \us31/n33 , \us31/n32 , \us31/n31 , \us31/n30 , \us31/n29 ,
         \us31/n28 , \us31/n27 , \us31/n26 , \us31/n25 , \us31/n24 ,
         \us31/n23 , \us31/n22 , \us31/n21 , \us31/n20 , \us31/n19 ,
         \us31/n18 , \us31/n17 , \us31/n16 , \us31/n15 , \us31/n14 ,
         \us31/n13 , \us31/n12 , \us31/n11 , \us31/n10 , \us31/n9 , \us31/n8 ,
         \us31/n7 , \us31/n6 , \us31/n5 , \us31/n4 , \us31/n3 , \us31/n2 ,
         \us31/n1 , \us32/n358 , \us32/n357 , \us32/n356 , \us32/n355 ,
         \us32/n354 , \us32/n353 , \us32/n352 , \us32/n351 , \us32/n350 ,
         \us32/n349 , \us32/n348 , \us32/n347 , \us32/n346 , \us32/n345 ,
         \us32/n344 , \us32/n343 , \us32/n342 , \us32/n341 , \us32/n340 ,
         \us32/n339 , \us32/n338 , \us32/n337 , \us32/n336 , \us32/n335 ,
         \us32/n334 , \us32/n333 , \us32/n332 , \us32/n331 , \us32/n330 ,
         \us32/n329 , \us32/n328 , \us32/n327 , \us32/n326 , \us32/n325 ,
         \us32/n324 , \us32/n323 , \us32/n322 , \us32/n321 , \us32/n320 ,
         \us32/n319 , \us32/n318 , \us32/n317 , \us32/n316 , \us32/n315 ,
         \us32/n314 , \us32/n313 , \us32/n312 , \us32/n311 , \us32/n310 ,
         \us32/n309 , \us32/n308 , \us32/n307 , \us32/n306 , \us32/n305 ,
         \us32/n304 , \us32/n303 , \us32/n302 , \us32/n301 , \us32/n300 ,
         \us32/n299 , \us32/n298 , \us32/n297 , \us32/n296 , \us32/n295 ,
         \us32/n294 , \us32/n293 , \us32/n292 , \us32/n291 , \us32/n290 ,
         \us32/n289 , \us32/n288 , \us32/n287 , \us32/n286 , \us32/n285 ,
         \us32/n284 , \us32/n283 , \us32/n282 , \us32/n281 , \us32/n280 ,
         \us32/n279 , \us32/n278 , \us32/n277 , \us32/n276 , \us32/n275 ,
         \us32/n274 , \us32/n273 , \us32/n272 , \us32/n271 , \us32/n270 ,
         \us32/n269 , \us32/n268 , \us32/n267 , \us32/n266 , \us32/n265 ,
         \us32/n264 , \us32/n263 , \us32/n262 , \us32/n261 , \us32/n260 ,
         \us32/n259 , \us32/n258 , \us32/n257 , \us32/n256 , \us32/n255 ,
         \us32/n254 , \us32/n253 , \us32/n252 , \us32/n251 , \us32/n250 ,
         \us32/n249 , \us32/n248 , \us32/n247 , \us32/n246 , \us32/n245 ,
         \us32/n244 , \us32/n243 , \us32/n242 , \us32/n241 , \us32/n240 ,
         \us32/n239 , \us32/n238 , \us32/n237 , \us32/n236 , \us32/n235 ,
         \us32/n234 , \us32/n233 , \us32/n232 , \us32/n231 , \us32/n230 ,
         \us32/n229 , \us32/n228 , \us32/n227 , \us32/n226 , \us32/n225 ,
         \us32/n224 , \us32/n223 , \us32/n222 , \us32/n221 , \us32/n220 ,
         \us32/n219 , \us32/n218 , \us32/n217 , \us32/n216 , \us32/n215 ,
         \us32/n214 , \us32/n213 , \us32/n212 , \us32/n211 , \us32/n210 ,
         \us32/n209 , \us32/n208 , \us32/n207 , \us32/n206 , \us32/n205 ,
         \us32/n204 , \us32/n203 , \us32/n202 , \us32/n201 , \us32/n200 ,
         \us32/n199 , \us32/n198 , \us32/n197 , \us32/n196 , \us32/n195 ,
         \us32/n194 , \us32/n193 , \us32/n192 , \us32/n191 , \us32/n190 ,
         \us32/n189 , \us32/n188 , \us32/n187 , \us32/n186 , \us32/n185 ,
         \us32/n184 , \us32/n183 , \us32/n182 , \us32/n181 , \us32/n180 ,
         \us32/n179 , \us32/n178 , \us32/n177 , \us32/n176 , \us32/n175 ,
         \us32/n174 , \us32/n173 , \us32/n172 , \us32/n171 , \us32/n170 ,
         \us32/n169 , \us32/n168 , \us32/n167 , \us32/n166 , \us32/n165 ,
         \us32/n164 , \us32/n163 , \us32/n162 , \us32/n161 , \us32/n160 ,
         \us32/n159 , \us32/n158 , \us32/n157 , \us32/n156 , \us32/n155 ,
         \us32/n154 , \us32/n153 , \us32/n152 , \us32/n151 , \us32/n150 ,
         \us32/n149 , \us32/n148 , \us32/n147 , \us32/n146 , \us32/n145 ,
         \us32/n144 , \us32/n143 , \us32/n142 , \us32/n141 , \us32/n140 ,
         \us32/n139 , \us32/n138 , \us32/n137 , \us32/n136 , \us32/n135 ,
         \us32/n134 , \us32/n133 , \us32/n132 , \us32/n131 , \us32/n130 ,
         \us32/n129 , \us32/n128 , \us32/n127 , \us32/n126 , \us32/n125 ,
         \us32/n124 , \us32/n123 , \us32/n122 , \us32/n121 , \us32/n120 ,
         \us32/n119 , \us32/n118 , \us32/n117 , \us32/n116 , \us32/n115 ,
         \us32/n114 , \us32/n113 , \us32/n112 , \us32/n111 , \us32/n110 ,
         \us32/n109 , \us32/n108 , \us32/n107 , \us32/n106 , \us32/n105 ,
         \us32/n104 , \us32/n103 , \us32/n102 , \us32/n101 , \us32/n100 ,
         \us32/n99 , \us32/n98 , \us32/n97 , \us32/n96 , \us32/n95 ,
         \us32/n94 , \us32/n93 , \us32/n92 , \us32/n91 , \us32/n90 ,
         \us32/n89 , \us32/n88 , \us32/n87 , \us32/n86 , \us32/n85 ,
         \us32/n84 , \us32/n83 , \us32/n82 , \us32/n81 , \us32/n80 ,
         \us32/n79 , \us32/n78 , \us32/n77 , \us32/n76 , \us32/n75 ,
         \us32/n74 , \us32/n73 , \us32/n72 , \us32/n71 , \us32/n70 ,
         \us32/n69 , \us32/n68 , \us32/n67 , \us32/n66 , \us32/n65 ,
         \us32/n64 , \us32/n63 , \us32/n62 , \us32/n61 , \us32/n60 ,
         \us32/n59 , \us32/n58 , \us32/n57 , \us32/n56 , \us32/n55 ,
         \us32/n54 , \us32/n53 , \us32/n52 , \us32/n51 , \us32/n50 ,
         \us32/n49 , \us32/n48 , \us32/n47 , \us32/n46 , \us32/n45 ,
         \us32/n44 , \us32/n43 , \us32/n42 , \us32/n41 , \us32/n40 ,
         \us32/n39 , \us32/n38 , \us32/n37 , \us32/n36 , \us32/n35 ,
         \us32/n34 , \us32/n33 , \us32/n32 , \us32/n31 , \us32/n30 ,
         \us32/n29 , \us32/n28 , \us32/n27 , \us32/n26 , \us32/n25 ,
         \us32/n24 , \us32/n23 , \us32/n22 , \us32/n21 , \us32/n20 ,
         \us32/n19 , \us32/n18 , \us32/n17 , \us32/n16 , \us32/n15 ,
         \us32/n14 , \us32/n13 , \us32/n12 , \us32/n11 , \us32/n10 , \us32/n9 ,
         \us32/n8 , \us32/n7 , \us32/n6 , \us32/n5 , \us32/n4 , \us32/n3 ,
         \us32/n2 , \us32/n1 , \us33/n358 , \us33/n357 , \us33/n356 ,
         \us33/n355 , \us33/n354 , \us33/n353 , \us33/n352 , \us33/n351 ,
         \us33/n350 , \us33/n349 , \us33/n348 , \us33/n347 , \us33/n346 ,
         \us33/n345 , \us33/n344 , \us33/n343 , \us33/n342 , \us33/n341 ,
         \us33/n340 , \us33/n339 , \us33/n338 , \us33/n337 , \us33/n336 ,
         \us33/n335 , \us33/n334 , \us33/n333 , \us33/n332 , \us33/n331 ,
         \us33/n330 , \us33/n329 , \us33/n328 , \us33/n327 , \us33/n326 ,
         \us33/n325 , \us33/n324 , \us33/n323 , \us33/n322 , \us33/n321 ,
         \us33/n320 , \us33/n319 , \us33/n318 , \us33/n317 , \us33/n316 ,
         \us33/n315 , \us33/n314 , \us33/n313 , \us33/n312 , \us33/n311 ,
         \us33/n310 , \us33/n309 , \us33/n308 , \us33/n307 , \us33/n306 ,
         \us33/n305 , \us33/n304 , \us33/n303 , \us33/n302 , \us33/n301 ,
         \us33/n300 , \us33/n299 , \us33/n298 , \us33/n297 , \us33/n296 ,
         \us33/n295 , \us33/n294 , \us33/n293 , \us33/n292 , \us33/n291 ,
         \us33/n290 , \us33/n289 , \us33/n288 , \us33/n287 , \us33/n286 ,
         \us33/n285 , \us33/n284 , \us33/n283 , \us33/n282 , \us33/n281 ,
         \us33/n280 , \us33/n279 , \us33/n278 , \us33/n277 , \us33/n276 ,
         \us33/n275 , \us33/n274 , \us33/n273 , \us33/n272 , \us33/n271 ,
         \us33/n270 , \us33/n269 , \us33/n268 , \us33/n267 , \us33/n266 ,
         \us33/n265 , \us33/n264 , \us33/n263 , \us33/n262 , \us33/n261 ,
         \us33/n260 , \us33/n259 , \us33/n258 , \us33/n257 , \us33/n256 ,
         \us33/n255 , \us33/n254 , \us33/n253 , \us33/n252 , \us33/n251 ,
         \us33/n250 , \us33/n249 , \us33/n248 , \us33/n247 , \us33/n246 ,
         \us33/n245 , \us33/n244 , \us33/n243 , \us33/n242 , \us33/n241 ,
         \us33/n240 , \us33/n239 , \us33/n238 , \us33/n237 , \us33/n236 ,
         \us33/n235 , \us33/n234 , \us33/n233 , \us33/n232 , \us33/n231 ,
         \us33/n230 , \us33/n229 , \us33/n228 , \us33/n227 , \us33/n226 ,
         \us33/n225 , \us33/n224 , \us33/n223 , \us33/n222 , \us33/n221 ,
         \us33/n220 , \us33/n219 , \us33/n218 , \us33/n217 , \us33/n216 ,
         \us33/n215 , \us33/n214 , \us33/n213 , \us33/n212 , \us33/n211 ,
         \us33/n210 , \us33/n209 , \us33/n208 , \us33/n207 , \us33/n206 ,
         \us33/n205 , \us33/n204 , \us33/n203 , \us33/n202 , \us33/n201 ,
         \us33/n200 , \us33/n199 , \us33/n198 , \us33/n197 , \us33/n196 ,
         \us33/n195 , \us33/n194 , \us33/n193 , \us33/n192 , \us33/n191 ,
         \us33/n190 , \us33/n189 , \us33/n188 , \us33/n187 , \us33/n186 ,
         \us33/n185 , \us33/n184 , \us33/n183 , \us33/n182 , \us33/n181 ,
         \us33/n180 , \us33/n179 , \us33/n178 , \us33/n177 , \us33/n176 ,
         \us33/n175 , \us33/n174 , \us33/n173 , \us33/n172 , \us33/n171 ,
         \us33/n170 , \us33/n169 , \us33/n168 , \us33/n167 , \us33/n166 ,
         \us33/n165 , \us33/n164 , \us33/n163 , \us33/n162 , \us33/n161 ,
         \us33/n160 , \us33/n159 , \us33/n158 , \us33/n157 , \us33/n156 ,
         \us33/n155 , \us33/n154 , \us33/n153 , \us33/n152 , \us33/n151 ,
         \us33/n150 , \us33/n149 , \us33/n148 , \us33/n147 , \us33/n146 ,
         \us33/n145 , \us33/n144 , \us33/n143 , \us33/n142 , \us33/n141 ,
         \us33/n140 , \us33/n139 , \us33/n138 , \us33/n137 , \us33/n136 ,
         \us33/n135 , \us33/n134 , \us33/n133 , \us33/n132 , \us33/n131 ,
         \us33/n130 , \us33/n129 , \us33/n128 , \us33/n127 , \us33/n126 ,
         \us33/n125 , \us33/n124 , \us33/n123 , \us33/n122 , \us33/n121 ,
         \us33/n120 , \us33/n119 , \us33/n118 , \us33/n117 , \us33/n116 ,
         \us33/n115 , \us33/n114 , \us33/n113 , \us33/n112 , \us33/n111 ,
         \us33/n110 , \us33/n109 , \us33/n108 , \us33/n107 , \us33/n106 ,
         \us33/n105 , \us33/n104 , \us33/n103 , \us33/n102 , \us33/n101 ,
         \us33/n100 , \us33/n99 , \us33/n98 , \us33/n97 , \us33/n96 ,
         \us33/n95 , \us33/n94 , \us33/n93 , \us33/n92 , \us33/n91 ,
         \us33/n90 , \us33/n89 , \us33/n88 , \us33/n87 , \us33/n86 ,
         \us33/n85 , \us33/n84 , \us33/n83 , \us33/n82 , \us33/n81 ,
         \us33/n80 , \us33/n79 , \us33/n78 , \us33/n77 , \us33/n76 ,
         \us33/n75 , \us33/n74 , \us33/n73 , \us33/n72 , \us33/n71 ,
         \us33/n70 , \us33/n69 , \us33/n68 , \us33/n67 , \us33/n66 ,
         \us33/n65 , \us33/n64 , \us33/n63 , \us33/n62 , \us33/n61 ,
         \us33/n60 , \us33/n59 , \us33/n58 , \us33/n57 , \us33/n56 ,
         \us33/n55 , \us33/n54 , \us33/n53 , \us33/n52 , \us33/n51 ,
         \us33/n50 , \us33/n49 , \us33/n48 , \us33/n47 , \us33/n46 ,
         \us33/n45 , \us33/n44 , \us33/n43 , \us33/n42 , \us33/n41 ,
         \us33/n40 , \us33/n39 , \us33/n38 , \us33/n37 , \us33/n36 ,
         \us33/n35 , \us33/n34 , \us33/n33 , \us33/n32 , \us33/n31 ,
         \us33/n30 , \us33/n29 , \us33/n28 , \us33/n27 , \us33/n26 ,
         \us33/n25 , \us33/n24 , \us33/n23 , \us33/n22 , \us33/n21 ,
         \us33/n20 , \us33/n19 , \us33/n18 , \us33/n17 , \us33/n16 ,
         \us33/n15 , \us33/n14 , \us33/n13 , \us33/n12 , \us33/n11 ,
         \us33/n10 , \us33/n9 , \us33/n8 , \us33/n7 , \us33/n6 , \us33/n5 ,
         \us33/n4 , \us33/n3 , \us33/n2 , \us33/n1 ;
  wire   [3:0] dcnt;
  wire   [127:0] text_in_r;
  wire   [31:0] w3;
  wire   [7:0] sa33;
  wire   [7:0] sa33_next;
  wire   [7:0] sa23;
  wire   [7:0] sa23_next;
  wire   [7:0] sa13;
  wire   [7:0] sa13_next;
  wire   [7:0] sa03;
  wire   [7:0] sa03_next;
  wire   [31:0] w2;
  wire   [7:0] sa32;
  wire   [7:0] sa32_next;
  wire   [7:0] sa22;
  wire   [7:0] sa22_next;
  wire   [7:0] sa12;
  wire   [7:0] sa12_next;
  wire   [7:0] sa02;
  wire   [7:0] sa02_next;
  wire   [31:0] w1;
  wire   [7:0] sa31;
  wire   [7:0] sa31_next;
  wire   [7:0] sa21;
  wire   [7:0] sa21_next;
  wire   [7:0] sa11;
  wire   [7:0] sa11_next;
  wire   [7:0] sa01;
  wire   [7:0] sa01_next;
  wire   [31:0] w0;
  wire   [7:0] sa30;
  wire   [7:0] sa30_next;
  wire   [7:0] sa20;
  wire   [7:0] sa20_next;
  wire   [7:0] sa10;
  wire   [7:0] sa10_next;
  wire   [7:0] sa00;
  wire   [7:0] sa00_next;
  wire   [7:0] sa00_sr;
  wire   [7:0] sa01_sr;
  wire   [7:0] sa02_sr;
  wire   [7:0] sa03_sr;
  wire   [7:0] sa10_sr;
  wire   [7:0] sa11_sr;
  wire   [7:0] sa12_sr;
  wire   [7:0] sa13_sr;
  wire   [7:0] sa20_sr;
  wire   [7:0] sa21_sr;
  wire   [7:0] sa22_sr;
  wire   [7:0] sa23_sr;
  wire   [7:0] sa30_sr;
  wire   [7:0] sa31_sr;
  wire   [7:0] sa32_sr;
  wire   [7:0] sa33_sr;
  wire   [31:0] \u0/rcon ;
  wire   [31:0] \u0/subword ;

  EDFFX1 \text_in_r_reg[127]  ( .D(text_in[127]), .E(ld), .CK(clk), .Q(
        text_in_r[127]) );
  EDFFX1 \text_in_r_reg[126]  ( .D(text_in[126]), .E(ld), .CK(clk), .Q(
        text_in_r[126]) );
  EDFFX1 \text_in_r_reg[125]  ( .D(text_in[125]), .E(ld), .CK(clk), .Q(
        text_in_r[125]) );
  EDFFX1 \text_in_r_reg[124]  ( .D(text_in[124]), .E(ld), .CK(clk), .Q(
        text_in_r[124]) );
  EDFFX1 \text_in_r_reg[123]  ( .D(text_in[123]), .E(ld), .CK(clk), .Q(
        text_in_r[123]) );
  EDFFX1 \text_in_r_reg[122]  ( .D(text_in[122]), .E(ld), .CK(clk), .Q(
        text_in_r[122]) );
  EDFFX1 \text_in_r_reg[121]  ( .D(text_in[121]), .E(ld), .CK(clk), .Q(
        text_in_r[121]) );
  EDFFX1 \text_in_r_reg[120]  ( .D(text_in[120]), .E(ld), .CK(clk), .Q(
        text_in_r[120]) );
  EDFFX1 \text_in_r_reg[119]  ( .D(text_in[119]), .E(ld), .CK(clk), .Q(
        text_in_r[119]) );
  EDFFX1 \text_in_r_reg[118]  ( .D(text_in[118]), .E(ld), .CK(clk), .Q(
        text_in_r[118]) );
  EDFFX1 \text_in_r_reg[117]  ( .D(text_in[117]), .E(ld), .CK(clk), .Q(
        text_in_r[117]) );
  EDFFX1 \text_in_r_reg[116]  ( .D(text_in[116]), .E(ld), .CK(clk), .Q(
        text_in_r[116]) );
  EDFFX1 \text_in_r_reg[115]  ( .D(text_in[115]), .E(ld), .CK(clk), .Q(
        text_in_r[115]) );
  EDFFX1 \text_in_r_reg[114]  ( .D(text_in[114]), .E(ld), .CK(clk), .Q(
        text_in_r[114]) );
  EDFFX1 \text_in_r_reg[113]  ( .D(text_in[113]), .E(ld), .CK(clk), .Q(
        text_in_r[113]) );
  EDFFX1 \text_in_r_reg[112]  ( .D(text_in[112]), .E(ld), .CK(clk), .Q(
        text_in_r[112]) );
  EDFFX1 \text_in_r_reg[111]  ( .D(text_in[111]), .E(ld), .CK(clk), .Q(
        text_in_r[111]) );
  EDFFX1 \text_in_r_reg[110]  ( .D(text_in[110]), .E(ld), .CK(clk), .Q(
        text_in_r[110]) );
  EDFFX1 \text_in_r_reg[109]  ( .D(text_in[109]), .E(ld), .CK(clk), .Q(
        text_in_r[109]) );
  EDFFX1 \text_in_r_reg[108]  ( .D(text_in[108]), .E(ld), .CK(clk), .Q(
        text_in_r[108]) );
  EDFFX1 \text_in_r_reg[107]  ( .D(text_in[107]), .E(ld), .CK(clk), .Q(
        text_in_r[107]) );
  EDFFX1 \text_in_r_reg[106]  ( .D(text_in[106]), .E(ld), .CK(clk), .Q(
        text_in_r[106]) );
  EDFFX1 \text_in_r_reg[105]  ( .D(text_in[105]), .E(ld), .CK(clk), .Q(
        text_in_r[105]) );
  EDFFX1 \text_in_r_reg[104]  ( .D(text_in[104]), .E(ld), .CK(clk), .Q(
        text_in_r[104]) );
  EDFFX1 \text_in_r_reg[103]  ( .D(text_in[103]), .E(ld), .CK(clk), .Q(
        text_in_r[103]) );
  EDFFX1 \text_in_r_reg[102]  ( .D(text_in[102]), .E(ld), .CK(clk), .Q(
        text_in_r[102]) );
  EDFFX1 \text_in_r_reg[101]  ( .D(text_in[101]), .E(ld), .CK(clk), .Q(
        text_in_r[101]) );
  EDFFX1 \text_in_r_reg[100]  ( .D(text_in[100]), .E(ld), .CK(clk), .Q(
        text_in_r[100]) );
  EDFFX1 \text_in_r_reg[99]  ( .D(text_in[99]), .E(ld), .CK(clk), .Q(
        text_in_r[99]) );
  EDFFX1 \text_in_r_reg[98]  ( .D(text_in[98]), .E(ld), .CK(clk), .Q(
        text_in_r[98]) );
  EDFFX1 \text_in_r_reg[97]  ( .D(text_in[97]), .E(ld), .CK(clk), .Q(
        text_in_r[97]) );
  EDFFX1 \text_in_r_reg[96]  ( .D(text_in[96]), .E(ld), .CK(clk), .Q(
        text_in_r[96]) );
  EDFFX1 \text_in_r_reg[95]  ( .D(text_in[95]), .E(ld), .CK(clk), .Q(
        text_in_r[95]) );
  EDFFX1 \text_in_r_reg[94]  ( .D(text_in[94]), .E(ld), .CK(clk), .Q(
        text_in_r[94]) );
  EDFFX1 \text_in_r_reg[93]  ( .D(text_in[93]), .E(ld), .CK(clk), .Q(
        text_in_r[93]) );
  EDFFX1 \text_in_r_reg[92]  ( .D(text_in[92]), .E(ld), .CK(clk), .Q(
        text_in_r[92]) );
  EDFFX1 \text_in_r_reg[91]  ( .D(text_in[91]), .E(ld), .CK(clk), .Q(
        text_in_r[91]) );
  EDFFX1 \text_in_r_reg[90]  ( .D(text_in[90]), .E(ld), .CK(clk), .Q(
        text_in_r[90]) );
  EDFFX1 \text_in_r_reg[89]  ( .D(text_in[89]), .E(ld), .CK(clk), .Q(
        text_in_r[89]) );
  EDFFX1 \text_in_r_reg[88]  ( .D(text_in[88]), .E(ld), .CK(clk), .Q(
        text_in_r[88]) );
  EDFFX1 \text_in_r_reg[87]  ( .D(text_in[87]), .E(ld), .CK(clk), .Q(
        text_in_r[87]) );
  EDFFX1 \text_in_r_reg[86]  ( .D(text_in[86]), .E(ld), .CK(clk), .Q(
        text_in_r[86]) );
  EDFFX1 \text_in_r_reg[85]  ( .D(text_in[85]), .E(ld), .CK(clk), .Q(
        text_in_r[85]) );
  EDFFX1 \text_in_r_reg[84]  ( .D(text_in[84]), .E(ld), .CK(clk), .Q(
        text_in_r[84]) );
  EDFFX1 \text_in_r_reg[83]  ( .D(text_in[83]), .E(ld), .CK(clk), .Q(
        text_in_r[83]) );
  EDFFX1 \text_in_r_reg[82]  ( .D(text_in[82]), .E(ld), .CK(clk), .Q(
        text_in_r[82]) );
  EDFFX1 \text_in_r_reg[81]  ( .D(text_in[81]), .E(ld), .CK(clk), .Q(
        text_in_r[81]) );
  EDFFX1 \text_in_r_reg[80]  ( .D(text_in[80]), .E(ld), .CK(clk), .Q(
        text_in_r[80]) );
  EDFFX1 \text_in_r_reg[79]  ( .D(text_in[79]), .E(ld), .CK(clk), .Q(
        text_in_r[79]) );
  EDFFX1 \text_in_r_reg[78]  ( .D(text_in[78]), .E(ld), .CK(clk), .Q(
        text_in_r[78]) );
  EDFFX1 \text_in_r_reg[77]  ( .D(text_in[77]), .E(ld), .CK(clk), .Q(
        text_in_r[77]) );
  EDFFX1 \text_in_r_reg[76]  ( .D(text_in[76]), .E(ld), .CK(clk), .Q(
        text_in_r[76]) );
  EDFFX1 \text_in_r_reg[75]  ( .D(text_in[75]), .E(ld), .CK(clk), .Q(
        text_in_r[75]) );
  EDFFX1 \text_in_r_reg[74]  ( .D(text_in[74]), .E(ld), .CK(clk), .Q(
        text_in_r[74]) );
  EDFFX1 \text_in_r_reg[73]  ( .D(text_in[73]), .E(ld), .CK(clk), .Q(
        text_in_r[73]) );
  EDFFX1 \text_in_r_reg[72]  ( .D(text_in[72]), .E(ld), .CK(clk), .Q(
        text_in_r[72]) );
  EDFFX1 \text_in_r_reg[71]  ( .D(text_in[71]), .E(ld), .CK(clk), .Q(
        text_in_r[71]) );
  EDFFX1 \text_in_r_reg[70]  ( .D(text_in[70]), .E(ld), .CK(clk), .Q(
        text_in_r[70]) );
  EDFFX1 \text_in_r_reg[69]  ( .D(text_in[69]), .E(ld), .CK(clk), .Q(
        text_in_r[69]) );
  EDFFX1 \text_in_r_reg[68]  ( .D(text_in[68]), .E(ld), .CK(clk), .Q(
        text_in_r[68]) );
  EDFFX1 \text_in_r_reg[67]  ( .D(text_in[67]), .E(ld), .CK(clk), .Q(
        text_in_r[67]) );
  EDFFX1 \text_in_r_reg[66]  ( .D(text_in[66]), .E(ld), .CK(clk), .Q(
        text_in_r[66]) );
  EDFFX1 \text_in_r_reg[65]  ( .D(text_in[65]), .E(ld), .CK(clk), .Q(
        text_in_r[65]) );
  EDFFX1 \text_in_r_reg[64]  ( .D(text_in[64]), .E(ld), .CK(clk), .Q(
        text_in_r[64]) );
  EDFFX1 \text_in_r_reg[63]  ( .D(text_in[63]), .E(ld), .CK(clk), .Q(
        text_in_r[63]) );
  EDFFX1 \text_in_r_reg[62]  ( .D(text_in[62]), .E(ld), .CK(clk), .Q(
        text_in_r[62]) );
  EDFFX1 \text_in_r_reg[61]  ( .D(text_in[61]), .E(ld), .CK(clk), .Q(
        text_in_r[61]) );
  EDFFX1 \text_in_r_reg[60]  ( .D(text_in[60]), .E(ld), .CK(clk), .Q(
        text_in_r[60]) );
  EDFFX1 \text_in_r_reg[59]  ( .D(text_in[59]), .E(ld), .CK(clk), .Q(
        text_in_r[59]) );
  EDFFX1 \text_in_r_reg[58]  ( .D(text_in[58]), .E(ld), .CK(clk), .Q(
        text_in_r[58]) );
  EDFFX1 \text_in_r_reg[57]  ( .D(text_in[57]), .E(ld), .CK(clk), .Q(
        text_in_r[57]) );
  EDFFX1 \text_in_r_reg[56]  ( .D(text_in[56]), .E(ld), .CK(clk), .Q(
        text_in_r[56]) );
  EDFFX1 \text_in_r_reg[55]  ( .D(text_in[55]), .E(ld), .CK(clk), .Q(
        text_in_r[55]) );
  EDFFX1 \text_in_r_reg[54]  ( .D(text_in[54]), .E(ld), .CK(clk), .Q(
        text_in_r[54]) );
  EDFFX1 \text_in_r_reg[53]  ( .D(text_in[53]), .E(ld), .CK(clk), .Q(
        text_in_r[53]) );
  EDFFX1 \text_in_r_reg[52]  ( .D(text_in[52]), .E(ld), .CK(clk), .Q(
        text_in_r[52]) );
  EDFFX1 \text_in_r_reg[51]  ( .D(text_in[51]), .E(ld), .CK(clk), .Q(
        text_in_r[51]) );
  EDFFX1 \text_in_r_reg[50]  ( .D(text_in[50]), .E(ld), .CK(clk), .Q(
        text_in_r[50]) );
  EDFFX1 \text_in_r_reg[49]  ( .D(text_in[49]), .E(ld), .CK(clk), .Q(
        text_in_r[49]) );
  EDFFX1 \text_in_r_reg[48]  ( .D(text_in[48]), .E(ld), .CK(clk), .Q(
        text_in_r[48]) );
  EDFFX1 \text_in_r_reg[47]  ( .D(text_in[47]), .E(ld), .CK(clk), .Q(
        text_in_r[47]) );
  EDFFX1 \text_in_r_reg[46]  ( .D(text_in[46]), .E(ld), .CK(clk), .Q(
        text_in_r[46]) );
  EDFFX1 \text_in_r_reg[45]  ( .D(text_in[45]), .E(ld), .CK(clk), .Q(
        text_in_r[45]) );
  EDFFX1 \text_in_r_reg[44]  ( .D(text_in[44]), .E(ld), .CK(clk), .Q(
        text_in_r[44]) );
  EDFFX1 \text_in_r_reg[43]  ( .D(text_in[43]), .E(ld), .CK(clk), .Q(
        text_in_r[43]) );
  EDFFX1 \text_in_r_reg[42]  ( .D(text_in[42]), .E(ld), .CK(clk), .Q(
        text_in_r[42]) );
  EDFFX1 \text_in_r_reg[41]  ( .D(text_in[41]), .E(ld), .CK(clk), .Q(
        text_in_r[41]) );
  EDFFX1 \text_in_r_reg[40]  ( .D(text_in[40]), .E(ld), .CK(clk), .Q(
        text_in_r[40]) );
  EDFFX1 \text_in_r_reg[39]  ( .D(text_in[39]), .E(ld), .CK(clk), .Q(
        text_in_r[39]) );
  EDFFX1 \text_in_r_reg[38]  ( .D(text_in[38]), .E(ld), .CK(clk), .Q(
        text_in_r[38]) );
  EDFFX1 \text_in_r_reg[37]  ( .D(text_in[37]), .E(ld), .CK(clk), .Q(
        text_in_r[37]) );
  EDFFX1 \text_in_r_reg[36]  ( .D(text_in[36]), .E(ld), .CK(clk), .Q(
        text_in_r[36]) );
  EDFFX1 \text_in_r_reg[35]  ( .D(text_in[35]), .E(ld), .CK(clk), .Q(
        text_in_r[35]) );
  EDFFX1 \text_in_r_reg[34]  ( .D(text_in[34]), .E(ld), .CK(clk), .Q(
        text_in_r[34]) );
  EDFFX1 \text_in_r_reg[33]  ( .D(text_in[33]), .E(ld), .CK(clk), .Q(
        text_in_r[33]) );
  EDFFX1 \text_in_r_reg[32]  ( .D(text_in[32]), .E(ld), .CK(clk), .Q(
        text_in_r[32]) );
  EDFFX1 \text_in_r_reg[31]  ( .D(text_in[31]), .E(ld), .CK(clk), .Q(
        text_in_r[31]) );
  EDFFX1 \text_in_r_reg[30]  ( .D(text_in[30]), .E(ld), .CK(clk), .Q(
        text_in_r[30]) );
  EDFFX1 \text_in_r_reg[29]  ( .D(text_in[29]), .E(ld), .CK(clk), .Q(
        text_in_r[29]) );
  EDFFX1 \text_in_r_reg[28]  ( .D(text_in[28]), .E(ld), .CK(clk), .Q(
        text_in_r[28]) );
  EDFFX1 \text_in_r_reg[27]  ( .D(text_in[27]), .E(ld), .CK(clk), .Q(
        text_in_r[27]) );
  EDFFX1 \text_in_r_reg[26]  ( .D(text_in[26]), .E(ld), .CK(clk), .Q(
        text_in_r[26]) );
  EDFFX1 \text_in_r_reg[25]  ( .D(text_in[25]), .E(ld), .CK(clk), .Q(
        text_in_r[25]) );
  EDFFX1 \text_in_r_reg[24]  ( .D(text_in[24]), .E(ld), .CK(clk), .Q(
        text_in_r[24]) );
  EDFFX1 \text_in_r_reg[23]  ( .D(text_in[23]), .E(ld), .CK(clk), .Q(
        text_in_r[23]) );
  EDFFX1 \text_in_r_reg[22]  ( .D(text_in[22]), .E(ld), .CK(clk), .Q(
        text_in_r[22]) );
  EDFFX1 \text_in_r_reg[21]  ( .D(text_in[21]), .E(ld), .CK(clk), .Q(
        text_in_r[21]) );
  EDFFX1 \text_in_r_reg[20]  ( .D(text_in[20]), .E(ld), .CK(clk), .Q(
        text_in_r[20]) );
  EDFFX1 \text_in_r_reg[19]  ( .D(text_in[19]), .E(ld), .CK(clk), .Q(
        text_in_r[19]) );
  EDFFX1 \text_in_r_reg[18]  ( .D(text_in[18]), .E(ld), .CK(clk), .Q(
        text_in_r[18]) );
  EDFFX1 \text_in_r_reg[17]  ( .D(text_in[17]), .E(ld), .CK(clk), .Q(
        text_in_r[17]) );
  EDFFX1 \text_in_r_reg[16]  ( .D(text_in[16]), .E(ld), .CK(clk), .Q(
        text_in_r[16]) );
  EDFFX1 \text_in_r_reg[15]  ( .D(text_in[15]), .E(ld), .CK(clk), .Q(
        text_in_r[15]) );
  EDFFX1 \text_in_r_reg[14]  ( .D(text_in[14]), .E(ld), .CK(clk), .Q(
        text_in_r[14]) );
  EDFFX1 \text_in_r_reg[13]  ( .D(text_in[13]), .E(ld), .CK(clk), .Q(
        text_in_r[13]) );
  EDFFX1 \text_in_r_reg[12]  ( .D(text_in[12]), .E(ld), .CK(clk), .Q(
        text_in_r[12]) );
  EDFFX1 \text_in_r_reg[11]  ( .D(text_in[11]), .E(ld), .CK(clk), .Q(
        text_in_r[11]) );
  EDFFX1 \text_in_r_reg[10]  ( .D(text_in[10]), .E(ld), .CK(clk), .Q(
        text_in_r[10]) );
  EDFFX1 \text_in_r_reg[9]  ( .D(text_in[9]), .E(ld), .CK(clk), .Q(
        text_in_r[9]) );
  EDFFX1 \text_in_r_reg[8]  ( .D(text_in[8]), .E(ld), .CK(clk), .Q(
        text_in_r[8]) );
  EDFFX1 \text_in_r_reg[7]  ( .D(text_in[7]), .E(ld), .CK(clk), .Q(
        text_in_r[7]) );
  EDFFX1 \text_in_r_reg[6]  ( .D(text_in[6]), .E(ld), .CK(clk), .Q(
        text_in_r[6]) );
  EDFFX1 \text_in_r_reg[5]  ( .D(text_in[5]), .E(ld), .CK(clk), .Q(
        text_in_r[5]) );
  EDFFX1 \text_in_r_reg[4]  ( .D(text_in[4]), .E(ld), .CK(clk), .Q(
        text_in_r[4]) );
  EDFFX1 \text_in_r_reg[3]  ( .D(text_in[3]), .E(ld), .CK(clk), .Q(
        text_in_r[3]) );
  EDFFX1 \text_in_r_reg[2]  ( .D(text_in[2]), .E(ld), .CK(clk), .Q(
        text_in_r[2]) );
  EDFFX1 \text_in_r_reg[1]  ( .D(text_in[1]), .E(ld), .CK(clk), .Q(
        text_in_r[1]) );
  EDFFX1 \text_in_r_reg[0]  ( .D(text_in[0]), .E(ld), .CK(clk), .Q(
        text_in_r[0]) );
  DFFX1 \dcnt_reg[2]  ( .D(n145), .CK(clk), .Q(n730) );
  DFFHQX1 \dcnt_reg[3]  ( .D(n1), .CK(clk), .Q(dcnt[3]) );
  DFFHQX1 \sa00_reg[0]  ( .D(N272), .CK(clk), .Q(sa00[0]) );
  DFFHQX1 \sa30_reg[0]  ( .D(N224), .CK(clk), .Q(sa30[0]) );
  DFFHQX1 \sa31_reg[0]  ( .D(N160), .CK(clk), .Q(sa31[0]) );
  DFFHQX1 \sa32_reg[0]  ( .D(N96), .CK(clk), .Q(sa32[0]) );
  DFFHQX1 \sa33_reg[0]  ( .D(N32), .CK(clk), .Q(sa33[0]) );
  DFFHQX1 \sa12_reg[0]  ( .D(N128), .CK(clk), .Q(sa12[0]) );
  DFFHQX1 \sa11_reg[0]  ( .D(N192), .CK(clk), .Q(sa11[0]) );
  DFFHQX1 \sa10_reg[0]  ( .D(N256), .CK(clk), .Q(sa10[0]) );
  DFFHQX1 \sa01_reg[0]  ( .D(N208), .CK(clk), .Q(sa01[0]) );
  DFFHQX1 \sa21_reg[0]  ( .D(N176), .CK(clk), .Q(sa21[0]) );
  DFFHQX1 \sa03_reg[0]  ( .D(N80), .CK(clk), .Q(sa03[0]) );
  DFFHQX1 \sa23_reg[0]  ( .D(N48), .CK(clk), .Q(sa23[0]) );
  DFFHQX1 \sa13_reg[0]  ( .D(N64), .CK(clk), .Q(sa13[0]) );
  DFFHQX1 \sa02_reg[0]  ( .D(N144), .CK(clk), .Q(sa02[0]) );
  DFFHQX1 \sa22_reg[0]  ( .D(N112), .CK(clk), .Q(sa22[0]) );
  DFFHQX1 \sa20_reg[0]  ( .D(N240), .CK(clk), .Q(sa20[0]) );
  DFFHQX1 \dcnt_reg[1]  ( .D(n146), .CK(clk), .Q(dcnt[1]) );
  DFFHQX1 \dcnt_reg[0]  ( .D(n147), .CK(clk), .Q(dcnt[0]) );
  DFFHQX1 \sa20_reg[7]  ( .D(N247), .CK(clk), .Q(sa20[7]) );
  DFFHQX1 \sa23_reg[7]  ( .D(N55), .CK(clk), .Q(sa23[7]) );
  DFFHQX1 \sa01_reg[7]  ( .D(N215), .CK(clk), .Q(sa01[7]) );
  DFFHQX1 \sa21_reg[7]  ( .D(N183), .CK(clk), .Q(sa21[7]) );
  DFFHQX1 \sa11_reg[7]  ( .D(N199), .CK(clk), .Q(sa11[7]) );
  DFFHQX1 \sa03_reg[7]  ( .D(N87), .CK(clk), .Q(sa03[7]) );
  DFFHQX1 \sa13_reg[7]  ( .D(N71), .CK(clk), .Q(sa13[7]) );
  DFFHQX1 \sa31_reg[7]  ( .D(N167), .CK(clk), .Q(sa31[7]) );
  DFFHQX1 \sa33_reg[7]  ( .D(N39), .CK(clk), .Q(sa33[7]) );
  DFFHQX1 \sa02_reg[7]  ( .D(N151), .CK(clk), .Q(sa02[7]) );
  DFFHQX1 \sa12_reg[7]  ( .D(N135), .CK(clk), .Q(sa12[7]) );
  DFFHQX1 \sa22_reg[7]  ( .D(N119), .CK(clk), .Q(sa22[7]) );
  DFFHQX1 \sa00_reg[7]  ( .D(N279), .CK(clk), .Q(sa00[7]) );
  DFFHQX1 \sa10_reg[7]  ( .D(N263), .CK(clk), .Q(sa10[7]) );
  DFFHQX1 \sa30_reg[7]  ( .D(N231), .CK(clk), .Q(sa30[7]) );
  DFFHQX1 \sa32_reg[7]  ( .D(N103), .CK(clk), .Q(sa32[7]) );
  DFFHQX1 \sa01_reg[5]  ( .D(N213), .CK(clk), .Q(sa01[5]) );
  DFFHQX1 \sa21_reg[5]  ( .D(N181), .CK(clk), .Q(sa21[5]) );
  DFFHQX1 \sa31_reg[5]  ( .D(N165), .CK(clk), .Q(sa31[5]) );
  DFFHQX1 \sa11_reg[5]  ( .D(N197), .CK(clk), .Q(sa11[5]) );
  DFFHQX1 \sa03_reg[5]  ( .D(N85), .CK(clk), .Q(sa03[5]) );
  DFFHQX1 \sa23_reg[5]  ( .D(N53), .CK(clk), .Q(sa23[5]) );
  DFFHQX1 \sa33_reg[5]  ( .D(N37), .CK(clk), .Q(sa33[5]) );
  DFFHQX1 \sa13_reg[5]  ( .D(N69), .CK(clk), .Q(sa13[5]) );
  DFFHQX1 \sa02_reg[5]  ( .D(N149), .CK(clk), .Q(sa02[5]) );
  DFFHQX1 \sa22_reg[5]  ( .D(N117), .CK(clk), .Q(sa22[5]) );
  DFFHQX1 \sa32_reg[5]  ( .D(N101), .CK(clk), .Q(sa32[5]) );
  DFFHQX1 \sa12_reg[5]  ( .D(N133), .CK(clk), .Q(sa12[5]) );
  DFFHQX1 \sa20_reg[5]  ( .D(N245), .CK(clk), .Q(sa20[5]) );
  DFFHQX1 \sa00_reg[5]  ( .D(N277), .CK(clk), .Q(sa00[5]) );
  DFFHQX1 \sa10_reg[5]  ( .D(N261), .CK(clk), .Q(sa10[5]) );
  DFFHQX1 \sa30_reg[5]  ( .D(N229), .CK(clk), .Q(sa30[5]) );
  DFFHQX1 \sa31_reg[3]  ( .D(N163), .CK(clk), .Q(sa31[3]) );
  DFFHQX1 \sa11_reg[3]  ( .D(N195), .CK(clk), .Q(sa11[3]) );
  DFFHQX1 \sa01_reg[3]  ( .D(N211), .CK(clk), .Q(sa01[3]) );
  DFFHQX1 \sa21_reg[3]  ( .D(N179), .CK(clk), .Q(sa21[3]) );
  DFFHQX1 \sa03_reg[3]  ( .D(N83), .CK(clk), .Q(sa03[3]) );
  DFFHQX1 \sa33_reg[3]  ( .D(N35), .CK(clk), .Q(sa33[3]) );
  DFFHQX1 \sa23_reg[3]  ( .D(N51), .CK(clk), .Q(sa23[3]) );
  DFFHQX1 \sa13_reg[3]  ( .D(N67), .CK(clk), .Q(sa13[3]) );
  DFFHQX1 \sa02_reg[3]  ( .D(N147), .CK(clk), .Q(sa02[3]) );
  DFFHQX1 \sa22_reg[3]  ( .D(N115), .CK(clk), .Q(sa22[3]) );
  DFFHQX1 \sa32_reg[3]  ( .D(N99), .CK(clk), .Q(sa32[3]) );
  DFFHQX1 \sa12_reg[3]  ( .D(N131), .CK(clk), .Q(sa12[3]) );
  DFFHQX1 \sa00_reg[3]  ( .D(N275), .CK(clk), .Q(sa00[3]) );
  DFFHQX1 \sa10_reg[3]  ( .D(N259), .CK(clk), .Q(sa10[3]) );
  DFFHQX1 \sa30_reg[3]  ( .D(N227), .CK(clk), .Q(sa30[3]) );
  DFFHQX1 \sa20_reg[3]  ( .D(N243), .CK(clk), .Q(sa20[3]) );
  DFFHQX1 \sa01_reg[2]  ( .D(N210), .CK(clk), .Q(sa01[2]) );
  DFFHQX1 \sa21_reg[2]  ( .D(N178), .CK(clk), .Q(sa21[2]) );
  DFFHQX1 \sa31_reg[2]  ( .D(N162), .CK(clk), .Q(sa31[2]) );
  DFFHQX1 \sa11_reg[2]  ( .D(N194), .CK(clk), .Q(sa11[2]) );
  DFFHQX1 \sa03_reg[2]  ( .D(N82), .CK(clk), .Q(sa03[2]) );
  DFFHQX1 \sa23_reg[2]  ( .D(N50), .CK(clk), .Q(sa23[2]) );
  DFFHQX1 \sa33_reg[2]  ( .D(N34), .CK(clk), .Q(sa33[2]) );
  DFFHQX1 \sa13_reg[2]  ( .D(N66), .CK(clk), .Q(sa13[2]) );
  DFFHQX1 \sa02_reg[2]  ( .D(N146), .CK(clk), .Q(sa02[2]) );
  DFFHQX1 \sa22_reg[2]  ( .D(N114), .CK(clk), .Q(sa22[2]) );
  DFFHQX1 \sa32_reg[2]  ( .D(N98), .CK(clk), .Q(sa32[2]) );
  DFFHQX1 \sa12_reg[2]  ( .D(N130), .CK(clk), .Q(sa12[2]) );
  DFFHQX1 \sa20_reg[2]  ( .D(N242), .CK(clk), .Q(sa20[2]) );
  DFFHQX1 \sa00_reg[2]  ( .D(N274), .CK(clk), .Q(sa00[2]) );
  DFFHQX1 \sa10_reg[2]  ( .D(N258), .CK(clk), .Q(sa10[2]) );
  DFFHQX1 \sa30_reg[2]  ( .D(N226), .CK(clk), .Q(sa30[2]) );
  DFFHQX1 \sa31_reg[4]  ( .D(N164), .CK(clk), .Q(sa31[4]) );
  DFFHQX1 \sa11_reg[4]  ( .D(N196), .CK(clk), .Q(sa11[4]) );
  DFFHQX1 \sa01_reg[4]  ( .D(N212), .CK(clk), .Q(sa01[4]) );
  DFFHQX1 \sa21_reg[4]  ( .D(N180), .CK(clk), .Q(sa21[4]) );
  DFFHQX1 \sa03_reg[4]  ( .D(N84), .CK(clk), .Q(sa03[4]) );
  DFFHQX1 \sa33_reg[4]  ( .D(N36), .CK(clk), .Q(sa33[4]) );
  DFFHQX1 \sa23_reg[4]  ( .D(N52), .CK(clk), .Q(sa23[4]) );
  DFFHQX1 \sa13_reg[4]  ( .D(N68), .CK(clk), .Q(sa13[4]) );
  DFFHQX1 \sa02_reg[4]  ( .D(N148), .CK(clk), .Q(sa02[4]) );
  DFFHQX1 \sa22_reg[4]  ( .D(N116), .CK(clk), .Q(sa22[4]) );
  DFFHQX1 \sa32_reg[4]  ( .D(N100), .CK(clk), .Q(sa32[4]) );
  DFFHQX1 \sa12_reg[4]  ( .D(N132), .CK(clk), .Q(sa12[4]) );
  DFFHQX1 \sa00_reg[4]  ( .D(N276), .CK(clk), .Q(sa00[4]) );
  DFFHQX1 \sa10_reg[4]  ( .D(N260), .CK(clk), .Q(sa10[4]) );
  DFFHQX1 \sa30_reg[4]  ( .D(N228), .CK(clk), .Q(sa30[4]) );
  DFFHQX1 \sa20_reg[4]  ( .D(N244), .CK(clk), .Q(sa20[4]) );
  DFFX1 ld_r_reg ( .D(ld), .CK(clk), .Q(n731), .QN(n580) );
  DFFHQX1 \sa01_reg[6]  ( .D(N214), .CK(clk), .Q(sa01[6]) );
  DFFHQX1 \sa21_reg[6]  ( .D(N182), .CK(clk), .Q(sa21[6]) );
  DFFHQX1 \sa31_reg[6]  ( .D(N166), .CK(clk), .Q(sa31[6]) );
  DFFHQX1 \sa11_reg[6]  ( .D(N198), .CK(clk), .Q(sa11[6]) );
  DFFHQX1 \sa03_reg[6]  ( .D(N86), .CK(clk), .Q(sa03[6]) );
  DFFHQX1 \sa23_reg[6]  ( .D(N54), .CK(clk), .Q(sa23[6]) );
  DFFHQX1 \sa33_reg[6]  ( .D(N38), .CK(clk), .Q(sa33[6]) );
  DFFHQX1 \sa13_reg[6]  ( .D(N70), .CK(clk), .Q(sa13[6]) );
  DFFHQX1 \sa02_reg[6]  ( .D(N150), .CK(clk), .Q(sa02[6]) );
  DFFHQX1 \sa22_reg[6]  ( .D(N118), .CK(clk), .Q(sa22[6]) );
  DFFHQX1 \sa32_reg[6]  ( .D(N102), .CK(clk), .Q(sa32[6]) );
  DFFHQX1 \sa12_reg[6]  ( .D(N134), .CK(clk), .Q(sa12[6]) );
  DFFHQX1 \sa20_reg[6]  ( .D(N246), .CK(clk), .Q(sa20[6]) );
  DFFHQX1 \sa00_reg[6]  ( .D(N278), .CK(clk), .Q(sa00[6]) );
  DFFHQX1 \sa10_reg[6]  ( .D(N262), .CK(clk), .Q(sa10[6]) );
  DFFHQX1 \sa30_reg[6]  ( .D(N230), .CK(clk), .Q(sa30[6]) );
  XOR2X1 U922 ( .A(w0[24]), .B(sa10_sr[0]), .Y(n166) );
  XOR2X1 U924 ( .A(n166), .B(n165), .Y(sa00_next[0]) );
  XOR2X1 U825 ( .A(w0[0]), .B(sa20_sr[0]), .Y(n237) );
  XOR2X1 U827 ( .A(n237), .B(n236), .Y(sa30_next[0]) );
  XOR2X1 U685 ( .A(w1[0]), .B(sa21_sr[0]), .Y(n327) );
  XOR2X1 U687 ( .A(n327), .B(n326), .Y(sa31_next[0]) );
  XOR2X1 U545 ( .A(w2[0]), .B(sa22_sr[0]), .Y(n417) );
  XOR2X1 U547 ( .A(n417), .B(n416), .Y(sa32_next[0]) );
  XOR2X1 U405 ( .A(w3[0]), .B(sa23_sr[0]), .Y(n507) );
  XOR2X1 U407 ( .A(n507), .B(n506), .Y(sa33_next[0]) );
  XOR2X1 U884 ( .A(w0[15]), .B(sa30_sr[7]), .Y(n194) );
  XOR2X1 U886 ( .A(n194), .B(n193), .Y(sa20_next[7]) );
  XOR2X1 U607 ( .A(w2[16]), .B(sa02_sr[0]), .Y(n372) );
  XOR2X1 U609 ( .A(n372), .B(n371), .Y(sa12_next[0]) );
  XOR2X1 U747 ( .A(w1[16]), .B(sa01_sr[0]), .Y(n282) );
  XOR2X1 U749 ( .A(n282), .B(n281), .Y(sa11_next[0]) );
  XOR2X1 U887 ( .A(w0[16]), .B(sa00_sr[0]), .Y(n192) );
  XOR2X1 U889 ( .A(n192), .B(n191), .Y(sa10_next[0]) );
  XOR2X1 U464 ( .A(w3[15]), .B(sa33_sr[7]), .Y(n464) );
  XOR2X1 U466 ( .A(n464), .B(n463), .Y(sa23_next[7]) );
  XOR2X1 U820 ( .A(w1[31]), .B(sa11_sr[7]), .Y(n239) );
  XOR2X1 U822 ( .A(n239), .B(n238), .Y(sa01_next[7]) );
  XOR2X1 U793 ( .A(n541), .B(n531), .Y(n250) );
  XOR2X1 U794 ( .A(n251), .B(n250), .Y(sa01_next[2]) );
  XOR2X1 U690 ( .A(n543), .B(n541), .Y(n323) );
  XOR2X1 U692 ( .A(n323), .B(n322), .Y(sa31_next[1]) );
  XOR2X1 U752 ( .A(n526), .B(n532), .Y(n278) );
  XOR2X1 U754 ( .A(n278), .B(n277), .Y(sa11_next[1]) );
  XOR2X1 U728 ( .A(n540), .B(n532), .Y(n295) );
  XOR2X1 U729 ( .A(n296), .B(n295), .Y(sa21_next[2]) );
  XOR2X1 U695 ( .A(n540), .B(n321), .Y(n319) );
  XOR2X1 U696 ( .A(n320), .B(n319), .Y(sa31_next[2]) );
  XOR2X1 U756 ( .A(sa11_sr[1]), .B(sa21_sr[1]), .Y(n275) );
  XOR2X1 U758 ( .A(n275), .B(n274), .Y(sa11_next[2]) );
  XOR2X1 U699 ( .A(n543), .B(n539), .Y(n316) );
  XOR2X1 U701 ( .A(n316), .B(n315), .Y(sa31_next[3]) );
  XOR2X1 U761 ( .A(n526), .B(n530), .Y(n271) );
  XOR2X1 U763 ( .A(n271), .B(n270), .Y(sa11_next[3]) );
  XOR2X1 U810 ( .A(w1[29]), .B(sa11_sr[5]), .Y(n243) );
  XOR2X1 U812 ( .A(n243), .B(n242), .Y(sa01_next[5]) );
  XOR2X1 U704 ( .A(n543), .B(n538), .Y(n312) );
  XOR2X1 U706 ( .A(n312), .B(n311), .Y(sa31_next[4]) );
  XOR2X1 U766 ( .A(n526), .B(n529), .Y(n267) );
  XOR2X1 U768 ( .A(n267), .B(n266), .Y(sa11_next[4]) );
  XOR2X1 U815 ( .A(w1[30]), .B(sa11_sr[6]), .Y(n241) );
  XOR2X1 U817 ( .A(n241), .B(n240), .Y(sa01_next[6]) );
  XOR2X1 U738 ( .A(w1[13]), .B(sa31_sr[5]), .Y(n288) );
  XOR2X1 U740 ( .A(n288), .B(n287), .Y(sa21_next[5]) );
  XOR2X1 U710 ( .A(n537), .B(n310), .Y(n308) );
  XOR2X1 U711 ( .A(n309), .B(n308), .Y(sa31_next[5]) );
  XOR2X1 U772 ( .A(n528), .B(n265), .Y(n263) );
  XOR2X1 U773 ( .A(n264), .B(n263), .Y(sa11_next[5]) );
  XOR2X1 U741 ( .A(w1[14]), .B(sa31_sr[6]), .Y(n286) );
  XOR2X1 U743 ( .A(n286), .B(n285), .Y(sa21_next[6]) );
  XOR2X1 U713 ( .A(sa21_sr[6]), .B(sa31_sr[5]), .Y(n306) );
  XOR2X1 U715 ( .A(n306), .B(n305), .Y(sa31_next[6]) );
  XOR2X1 U775 ( .A(sa11_sr[5]), .B(sa21_sr[5]), .Y(n261) );
  XOR2X1 U777 ( .A(n261), .B(n260), .Y(sa11_next[6]) );
  XOR2X1 U804 ( .A(n535), .B(n539), .Y(n245) );
  XOR2X1 U806 ( .A(n245), .B(n244), .Y(sa01_next[4]) );
  XOR2X1 U798 ( .A(n535), .B(n540), .Y(n248) );
  XOR2X1 U800 ( .A(n248), .B(n247), .Y(sa01_next[3]) );
  XOR2X1 U787 ( .A(n535), .B(n542), .Y(n253) );
  XOR2X1 U789 ( .A(n253), .B(n252), .Y(sa01_next[1]) );
  XOR2X1 U782 ( .A(w1[24]), .B(sa11_sr[0]), .Y(n256) );
  XOR2X1 U784 ( .A(n256), .B(n255), .Y(sa01_next[0]) );
  XOR2X1 U744 ( .A(w1[15]), .B(sa31_sr[7]), .Y(n284) );
  XOR2X1 U746 ( .A(n284), .B(n283), .Y(sa21_next[7]) );
  XOR2X1 U779 ( .A(sa11_sr[6]), .B(sa21_sr[6]), .Y(n258) );
  XOR2X1 U781 ( .A(n258), .B(n257), .Y(sa11_next[7]) );
  XOR2X1 U735 ( .A(n534), .B(n538), .Y(n290) );
  XOR2X1 U737 ( .A(n290), .B(n289), .Y(sa21_next[4]) );
  XOR2X1 U731 ( .A(n534), .B(n539), .Y(n293) );
  XOR2X1 U733 ( .A(n293), .B(n292), .Y(sa21_next[3]) );
  XOR2X1 U724 ( .A(n534), .B(n541), .Y(n298) );
  XOR2X1 U726 ( .A(n298), .B(n297), .Y(sa21_next[1]) );
  XOR2X1 U720 ( .A(w1[8]), .B(sa31_sr[0]), .Y(n301) );
  XOR2X1 U722 ( .A(n301), .B(n300), .Y(sa21_next[0]) );
  XOR2X1 U502 ( .A(w3[24]), .B(sa13_sr[0]), .Y(n436) );
  XOR2X1 U504 ( .A(n436), .B(n435), .Y(sa03_next[0]) );
  XOR2X1 U540 ( .A(w3[31]), .B(sa13_sr[7]), .Y(n419) );
  XOR2X1 U542 ( .A(n419), .B(n418), .Y(sa03_next[7]) );
  XOR2X1 U507 ( .A(n571), .B(n578), .Y(n433) );
  XOR2X1 U509 ( .A(n433), .B(n432), .Y(sa03_next[1]) );
  XOR2X1 U513 ( .A(n577), .B(n567), .Y(n430) );
  XOR2X1 U514 ( .A(n431), .B(n430), .Y(sa03_next[2]) );
  XOR2X1 U410 ( .A(n579), .B(n577), .Y(n503) );
  XOR2X1 U412 ( .A(n503), .B(n502), .Y(sa33_next[1]) );
  XOR2X1 U518 ( .A(n571), .B(n576), .Y(n428) );
  XOR2X1 U520 ( .A(n428), .B(n427), .Y(sa03_next[3]) );
  XOR2X1 U448 ( .A(n576), .B(n568), .Y(n475) );
  XOR2X1 U449 ( .A(n476), .B(n475), .Y(sa23_next[2]) );
  XOR2X1 U415 ( .A(n576), .B(n501), .Y(n499) );
  XOR2X1 U416 ( .A(n500), .B(n499), .Y(sa33_next[2]) );
  XOR2X1 U476 ( .A(sa13_sr[1]), .B(sa23_sr[1]), .Y(n455) );
  XOR2X1 U478 ( .A(n455), .B(n454), .Y(sa13_next[2]) );
  XOR2X1 U524 ( .A(n571), .B(n575), .Y(n425) );
  XOR2X1 U526 ( .A(n425), .B(n424), .Y(sa03_next[4]) );
  XOR2X1 U419 ( .A(n579), .B(n575), .Y(n496) );
  XOR2X1 U421 ( .A(n496), .B(n495), .Y(sa33_next[3]) );
  XOR2X1 U530 ( .A(w3[29]), .B(sa13_sr[5]), .Y(n423) );
  XOR2X1 U532 ( .A(n423), .B(n422), .Y(sa03_next[5]) );
  XOR2X1 U424 ( .A(n579), .B(n574), .Y(n492) );
  XOR2X1 U426 ( .A(n492), .B(n491), .Y(sa33_next[4]) );
  XOR2X1 U535 ( .A(w3[30]), .B(sa13_sr[6]), .Y(n421) );
  XOR2X1 U537 ( .A(n421), .B(n420), .Y(sa03_next[6]) );
  XOR2X1 U458 ( .A(w3[13]), .B(sa33_sr[5]), .Y(n468) );
  XOR2X1 U460 ( .A(n468), .B(n467), .Y(sa23_next[5]) );
  XOR2X1 U430 ( .A(n573), .B(n490), .Y(n488) );
  XOR2X1 U431 ( .A(n489), .B(n488), .Y(sa33_next[5]) );
  XOR2X1 U492 ( .A(n564), .B(n445), .Y(n443) );
  XOR2X1 U493 ( .A(n444), .B(n443), .Y(sa13_next[5]) );
  XOR2X1 U461 ( .A(w3[14]), .B(sa33_sr[6]), .Y(n466) );
  XOR2X1 U463 ( .A(n466), .B(n465), .Y(sa23_next[6]) );
  XOR2X1 U433 ( .A(sa23_sr[6]), .B(sa33_sr[5]), .Y(n486) );
  XOR2X1 U435 ( .A(n486), .B(n485), .Y(sa33_next[6]) );
  XOR2X1 U495 ( .A(sa13_sr[5]), .B(sa23_sr[5]), .Y(n441) );
  XOR2X1 U497 ( .A(n441), .B(n440), .Y(sa13_next[6]) );
  XOR2X1 U499 ( .A(sa13_sr[6]), .B(sa23_sr[6]), .Y(n438) );
  XOR2X1 U501 ( .A(n438), .B(n437), .Y(sa13_next[7]) );
  XOR2X1 U455 ( .A(n570), .B(n574), .Y(n470) );
  XOR2X1 U457 ( .A(n470), .B(n469), .Y(sa23_next[4]) );
  XOR2X1 U451 ( .A(n570), .B(n575), .Y(n473) );
  XOR2X1 U453 ( .A(n473), .B(n472), .Y(sa23_next[3]) );
  XOR2X1 U444 ( .A(n570), .B(n577), .Y(n478) );
  XOR2X1 U446 ( .A(n478), .B(n477), .Y(sa23_next[1]) );
  XOR2X1 U440 ( .A(w3[8]), .B(sa33_sr[0]), .Y(n481) );
  XOR2X1 U442 ( .A(n481), .B(n480), .Y(sa23_next[0]) );
  XOR2X1 U717 ( .A(sa21_sr[7]), .B(sa31_sr[6]), .Y(n303) );
  XOR2X1 U719 ( .A(n303), .B(n302), .Y(sa31_next[7]) );
  XOR2X1 U437 ( .A(sa23_sr[7]), .B(sa33_sr[6]), .Y(n483) );
  XOR2X1 U439 ( .A(n483), .B(n482), .Y(sa33_next[7]) );
  XOR2X1 U486 ( .A(n562), .B(n565), .Y(n447) );
  XOR2X1 U488 ( .A(n447), .B(n446), .Y(sa13_next[4]) );
  XOR2X1 U481 ( .A(n562), .B(n566), .Y(n451) );
  XOR2X1 U483 ( .A(n451), .B(n450), .Y(sa13_next[3]) );
  XOR2X1 U472 ( .A(n562), .B(n568), .Y(n458) );
  XOR2X1 U474 ( .A(n458), .B(n457), .Y(sa13_next[1]) );
  XOR2X1 U467 ( .A(w3[16]), .B(sa03_sr[0]), .Y(n462) );
  XOR2X1 U469 ( .A(n462), .B(n461), .Y(sa13_next[0]) );
  XOR2X1 U642 ( .A(w2[24]), .B(sa12_sr[0]), .Y(n346) );
  XOR2X1 U644 ( .A(n346), .B(n345), .Y(sa02_next[0]) );
  XOR2X1 U647 ( .A(n553), .B(n560), .Y(n343) );
  XOR2X1 U649 ( .A(n343), .B(n342), .Y(sa02_next[1]) );
  XOR2X1 U653 ( .A(n559), .B(n549), .Y(n340) );
  XOR2X1 U654 ( .A(n341), .B(n340), .Y(sa02_next[2]) );
  XOR2X1 U550 ( .A(n561), .B(n559), .Y(n413) );
  XOR2X1 U552 ( .A(n413), .B(n412), .Y(sa32_next[1]) );
  XOR2X1 U612 ( .A(n544), .B(n550), .Y(n368) );
  XOR2X1 U614 ( .A(n368), .B(n367), .Y(sa12_next[1]) );
  XOR2X1 U658 ( .A(n553), .B(n558), .Y(n338) );
  XOR2X1 U660 ( .A(n338), .B(n337), .Y(sa02_next[3]) );
  XOR2X1 U555 ( .A(n558), .B(n411), .Y(n409) );
  XOR2X1 U556 ( .A(n410), .B(n409), .Y(sa32_next[2]) );
  XOR2X1 U616 ( .A(sa12_sr[1]), .B(sa22_sr[1]), .Y(n365) );
  XOR2X1 U618 ( .A(n365), .B(n364), .Y(sa12_next[2]) );
  XOR2X1 U664 ( .A(n553), .B(n557), .Y(n335) );
  XOR2X1 U666 ( .A(n335), .B(n334), .Y(sa02_next[4]) );
  XOR2X1 U559 ( .A(n561), .B(n557), .Y(n406) );
  XOR2X1 U561 ( .A(n406), .B(n405), .Y(sa32_next[3]) );
  XOR2X1 U621 ( .A(n544), .B(n548), .Y(n361) );
  XOR2X1 U623 ( .A(n361), .B(n360), .Y(sa12_next[3]) );
  XOR2X1 U670 ( .A(w2[29]), .B(sa12_sr[5]), .Y(n333) );
  XOR2X1 U672 ( .A(n333), .B(n332), .Y(sa02_next[5]) );
  XOR2X1 U626 ( .A(n544), .B(n547), .Y(n357) );
  XOR2X1 U628 ( .A(n357), .B(n356), .Y(sa12_next[4]) );
  XOR2X1 U675 ( .A(w2[30]), .B(sa12_sr[6]), .Y(n331) );
  XOR2X1 U677 ( .A(n331), .B(n330), .Y(sa02_next[6]) );
  XOR2X1 U632 ( .A(n546), .B(n355), .Y(n353) );
  XOR2X1 U633 ( .A(n354), .B(n353), .Y(sa12_next[5]) );
  XOR2X1 U680 ( .A(w2[31]), .B(sa12_sr[7]), .Y(n329) );
  XOR2X1 U682 ( .A(n329), .B(n328), .Y(sa02_next[7]) );
  XOR2X1 U635 ( .A(sa12_sr[5]), .B(sa22_sr[5]), .Y(n351) );
  XOR2X1 U637 ( .A(n351), .B(n350), .Y(sa12_next[6]) );
  XOR2X1 U639 ( .A(sa12_sr[6]), .B(sa22_sr[6]), .Y(n348) );
  XOR2X1 U641 ( .A(n348), .B(n347), .Y(sa12_next[7]) );
  XOR2X1 U604 ( .A(w2[15]), .B(sa32_sr[7]), .Y(n374) );
  XOR2X1 U606 ( .A(n374), .B(n373), .Y(sa22_next[7]) );
  XOR2X1 U927 ( .A(n517), .B(n524), .Y(n163) );
  XOR2X1 U929 ( .A(n163), .B(n162), .Y(sa00_next[1]) );
  XOR2X1 U892 ( .A(n508), .B(n514), .Y(n188) );
  XOR2X1 U894 ( .A(n188), .B(n187), .Y(sa10_next[1]) );
  XOR2X1 U868 ( .A(n522), .B(n514), .Y(n205) );
  XOR2X1 U869 ( .A(n206), .B(n205), .Y(sa20_next[2]) );
  XOR2X1 U830 ( .A(n525), .B(n523), .Y(n233) );
  XOR2X1 U832 ( .A(n233), .B(n232), .Y(sa30_next[1]) );
  XOR2X1 U933 ( .A(n523), .B(n513), .Y(n160) );
  XOR2X1 U934 ( .A(n161), .B(n160), .Y(sa00_next[2]) );
  XOR2X1 U896 ( .A(sa10_sr[1]), .B(sa20_sr[1]), .Y(n185) );
  XOR2X1 U898 ( .A(n185), .B(n184), .Y(sa10_next[2]) );
  XOR2X1 U835 ( .A(n522), .B(n231), .Y(n229) );
  XOR2X1 U836 ( .A(n230), .B(n229), .Y(sa30_next[2]) );
  XOR2X1 U938 ( .A(n517), .B(n522), .Y(n158) );
  XOR2X1 U940 ( .A(n158), .B(n157), .Y(sa00_next[3]) );
  XOR2X1 U901 ( .A(n508), .B(n512), .Y(n181) );
  XOR2X1 U903 ( .A(n181), .B(n180), .Y(sa10_next[3]) );
  XOR2X1 U839 ( .A(n525), .B(n521), .Y(n226) );
  XOR2X1 U841 ( .A(n226), .B(n225), .Y(sa30_next[3]) );
  XOR2X1 U944 ( .A(n517), .B(n521), .Y(n155) );
  XOR2X1 U946 ( .A(n155), .B(n154), .Y(sa00_next[4]) );
  XOR2X1 U906 ( .A(n508), .B(n511), .Y(n177) );
  XOR2X1 U908 ( .A(n177), .B(n176), .Y(sa10_next[4]) );
  XOR2X1 U878 ( .A(w0[13]), .B(sa30_sr[5]), .Y(n198) );
  XOR2X1 U880 ( .A(n198), .B(n197), .Y(sa20_next[5]) );
  XOR2X1 U844 ( .A(n525), .B(n520), .Y(n222) );
  XOR2X1 U846 ( .A(n222), .B(n221), .Y(sa30_next[4]) );
  XOR2X1 U950 ( .A(w0[29]), .B(sa10_sr[5]), .Y(n153) );
  XOR2X1 U952 ( .A(n153), .B(n152), .Y(sa00_next[5]) );
  XOR2X1 U912 ( .A(n510), .B(n175), .Y(n173) );
  XOR2X1 U913 ( .A(n174), .B(n173), .Y(sa10_next[5]) );
  XOR2X1 U881 ( .A(w0[14]), .B(sa30_sr[6]), .Y(n196) );
  XOR2X1 U883 ( .A(n196), .B(n195), .Y(sa20_next[6]) );
  XOR2X1 U850 ( .A(n519), .B(n220), .Y(n218) );
  XOR2X1 U851 ( .A(n219), .B(n218), .Y(sa30_next[5]) );
  XOR2X1 U955 ( .A(w0[30]), .B(sa10_sr[6]), .Y(n151) );
  XOR2X1 U957 ( .A(n151), .B(n150), .Y(sa00_next[6]) );
  XOR2X1 U915 ( .A(sa10_sr[5]), .B(sa20_sr[5]), .Y(n171) );
  XOR2X1 U917 ( .A(n171), .B(n170), .Y(sa10_next[6]) );
  XOR2X1 U853 ( .A(sa20_sr[6]), .B(sa30_sr[5]), .Y(n216) );
  XOR2X1 U855 ( .A(n216), .B(n215), .Y(sa30_next[6]) );
  XOR2X1 U960 ( .A(w0[31]), .B(sa10_sr[7]), .Y(n149) );
  XOR2X1 U962 ( .A(n149), .B(n148), .Y(sa00_next[7]) );
  XOR2X1 U919 ( .A(sa10_sr[6]), .B(sa20_sr[6]), .Y(n168) );
  XOR2X1 U921 ( .A(n168), .B(n167), .Y(sa10_next[7]) );
  XOR2X1 U875 ( .A(n516), .B(n520), .Y(n200) );
  XOR2X1 U877 ( .A(n200), .B(n199), .Y(sa20_next[4]) );
  XOR2X1 U871 ( .A(n516), .B(n521), .Y(n203) );
  XOR2X1 U873 ( .A(n203), .B(n202), .Y(sa20_next[3]) );
  XOR2X1 U864 ( .A(n516), .B(n523), .Y(n208) );
  XOR2X1 U866 ( .A(n208), .B(n207), .Y(sa20_next[1]) );
  XOR2X1 U860 ( .A(w0[8]), .B(sa30_sr[0]), .Y(n211) );
  XOR2X1 U862 ( .A(n211), .B(n210), .Y(sa20_next[0]) );
  XOR2X1 U857 ( .A(sa20_sr[7]), .B(sa30_sr[6]), .Y(n213) );
  XOR2X1 U859 ( .A(n213), .B(n212), .Y(sa30_next[7]) );
  XOR2X1 U580 ( .A(w2[8]), .B(sa32_sr[0]), .Y(n391) );
  XOR2X1 U582 ( .A(n391), .B(n390), .Y(sa22_next[0]) );
  XOR2X1 U584 ( .A(n552), .B(n559), .Y(n388) );
  XOR2X1 U586 ( .A(n388), .B(n387), .Y(sa22_next[1]) );
  XOR2X1 U588 ( .A(n558), .B(n550), .Y(n385) );
  XOR2X1 U589 ( .A(n386), .B(n385), .Y(sa22_next[2]) );
  XOR2X1 U591 ( .A(n552), .B(n557), .Y(n383) );
  XOR2X1 U593 ( .A(n383), .B(n382), .Y(sa22_next[3]) );
  XOR2X1 U595 ( .A(n552), .B(n556), .Y(n380) );
  XOR2X1 U597 ( .A(n380), .B(n379), .Y(sa22_next[4]) );
  XOR2X1 U564 ( .A(n561), .B(n556), .Y(n402) );
  XOR2X1 U566 ( .A(n402), .B(n401), .Y(sa32_next[4]) );
  XOR2X1 U598 ( .A(w2[13]), .B(sa32_sr[5]), .Y(n378) );
  XOR2X1 U600 ( .A(n378), .B(n377), .Y(sa22_next[5]) );
  XOR2X1 U570 ( .A(n555), .B(n400), .Y(n398) );
  XOR2X1 U571 ( .A(n399), .B(n398), .Y(sa32_next[5]) );
  XOR2X1 U601 ( .A(w2[14]), .B(sa32_sr[6]), .Y(n376) );
  XOR2X1 U603 ( .A(n376), .B(n375), .Y(sa22_next[6]) );
  XOR2X1 U573 ( .A(sa22_sr[6]), .B(sa32_sr[5]), .Y(n396) );
  XOR2X1 U575 ( .A(n396), .B(n395), .Y(sa32_next[6]) );
  XOR2X1 U577 ( .A(sa22_sr[7]), .B(sa32_sr[6]), .Y(n393) );
  XOR2X1 U579 ( .A(n393), .B(n392), .Y(sa32_next[7]) );
  XOR2X1 U712 ( .A(w1[6]), .B(sa01_sr[5]), .Y(n307) );
  XOR2X1 U714 ( .A(n536), .B(n307), .Y(n305) );
  XOR2X1 U797 ( .A(w1[27]), .B(sa11_sr[3]), .Y(n249) );
  XOR2X1 U799 ( .A(n530), .B(n249), .Y(n247) );
  XOR2X1 U517 ( .A(w3[27]), .B(sa13_sr[3]), .Y(n429) );
  XOR2X1 U519 ( .A(n566), .B(n429), .Y(n427) );
  XOR2X1 U432 ( .A(w3[6]), .B(sa03_sr[5]), .Y(n487) );
  XOR2X1 U434 ( .A(n572), .B(n487), .Y(n485) );
  XOR2X1 U657 ( .A(w2[27]), .B(sa12_sr[3]), .Y(n339) );
  XOR2X1 U659 ( .A(n548), .B(n339), .Y(n337) );
  XOR2X1 U572 ( .A(w2[6]), .B(sa02_sr[5]), .Y(n397) );
  XOR2X1 U574 ( .A(n554), .B(n397), .Y(n395) );
  XOR2X1 U937 ( .A(w0[27]), .B(sa10_sr[3]), .Y(n159) );
  XOR2X1 U939 ( .A(n512), .B(n159), .Y(n157) );
  XOR2X1 U852 ( .A(w0[6]), .B(sa00_sr[5]), .Y(n217) );
  XOR2X1 U854 ( .A(n518), .B(n217), .Y(n215) );
  XOR2X1 U730 ( .A(w1[11]), .B(sa31_sr[3]), .Y(n294) );
  XOR2X1 U732 ( .A(n531), .B(n294), .Y(n292) );
  XOR2X1 U450 ( .A(w3[11]), .B(sa33_sr[3]), .Y(n474) );
  XOR2X1 U452 ( .A(n567), .B(n474), .Y(n472) );
  XOR2X1 U590 ( .A(w2[11]), .B(sa32_sr[3]), .Y(n384) );
  XOR2X1 U592 ( .A(n549), .B(n384), .Y(n382) );
  XOR2X1 U870 ( .A(w0[11]), .B(sa30_sr[3]), .Y(n204) );
  XOR2X1 U872 ( .A(n513), .B(n204), .Y(n202) );
  XOR2X1 U689 ( .A(sa21_sr[1]), .B(sa31_sr[0]), .Y(n324) );
  XOR2X1 U688 ( .A(w1[1]), .B(sa01_sr[0]), .Y(n325) );
  XOR2X1 U691 ( .A(n325), .B(n324), .Y(n322) );
  XOR2X1 U409 ( .A(sa23_sr[1]), .B(sa33_sr[0]), .Y(n504) );
  XOR2X1 U408 ( .A(w3[1]), .B(sa03_sr[0]), .Y(n505) );
  XOR2X1 U411 ( .A(n505), .B(n504), .Y(n502) );
  XOR2X1 U549 ( .A(sa22_sr[1]), .B(sa32_sr[0]), .Y(n414) );
  XOR2X1 U548 ( .A(w2[1]), .B(sa02_sr[0]), .Y(n415) );
  XOR2X1 U551 ( .A(n415), .B(n414), .Y(n412) );
  XOR2X1 U829 ( .A(sa20_sr[1]), .B(sa30_sr[0]), .Y(n234) );
  XOR2X1 U828 ( .A(w0[1]), .B(sa00_sr[0]), .Y(n235) );
  XOR2X1 U831 ( .A(n235), .B(n234), .Y(n232) );
  XOR2X1 U774 ( .A(w1[22]), .B(sa01_sr[6]), .Y(n262) );
  XOR2X1 U776 ( .A(n527), .B(n262), .Y(n260) );
  XOR2X1 U786 ( .A(w1[25]), .B(sa11_sr[1]), .Y(n254) );
  XOR2X1 U788 ( .A(n532), .B(n254), .Y(n252) );
  XOR2X1 U506 ( .A(w3[25]), .B(sa13_sr[1]), .Y(n434) );
  XOR2X1 U508 ( .A(n568), .B(n434), .Y(n432) );
  XOR2X1 U494 ( .A(w3[22]), .B(sa03_sr[6]), .Y(n442) );
  XOR2X1 U496 ( .A(n563), .B(n442), .Y(n440) );
  XOR2X1 U646 ( .A(w2[25]), .B(sa12_sr[1]), .Y(n344) );
  XOR2X1 U648 ( .A(n550), .B(n344), .Y(n342) );
  XOR2X1 U634 ( .A(w2[22]), .B(sa02_sr[6]), .Y(n352) );
  XOR2X1 U636 ( .A(n545), .B(n352), .Y(n350) );
  XOR2X1 U926 ( .A(w0[25]), .B(sa10_sr[1]), .Y(n164) );
  XOR2X1 U928 ( .A(n514), .B(n164), .Y(n162) );
  XOR2X1 U914 ( .A(w0[22]), .B(sa00_sr[6]), .Y(n172) );
  XOR2X1 U916 ( .A(n509), .B(n172), .Y(n170) );
  XOR2XL U755 ( .A(w1[18]), .B(sa01_sr[2]), .Y(n276) );
  XOR2X1 U757 ( .A(n531), .B(n276), .Y(n274) );
  XOR2XL U475 ( .A(w3[18]), .B(sa03_sr[2]), .Y(n456) );
  XOR2X1 U477 ( .A(n567), .B(n456), .Y(n454) );
  XOR2XL U615 ( .A(w2[18]), .B(sa02_sr[2]), .Y(n366) );
  XOR2X1 U617 ( .A(n549), .B(n366), .Y(n364) );
  XOR2XL U895 ( .A(w0[18]), .B(sa00_sr[2]), .Y(n186) );
  XOR2X1 U897 ( .A(n513), .B(n186), .Y(n184) );
  XOR2X1 U751 ( .A(sa11_sr[0]), .B(sa21_sr[0]), .Y(n279) );
  XOR2X1 U750 ( .A(w1[17]), .B(sa01_sr[1]), .Y(n280) );
  XOR2X1 U753 ( .A(n280), .B(n279), .Y(n277) );
  XOR2X1 U765 ( .A(sa11_sr[3]), .B(sa21_sr[3]), .Y(n268) );
  XOR2XL U764 ( .A(w1[20]), .B(sa01_sr[4]), .Y(n269) );
  XOR2X1 U767 ( .A(n269), .B(n268), .Y(n266) );
  XOR2X1 U485 ( .A(sa13_sr[3]), .B(sa23_sr[3]), .Y(n448) );
  XOR2XL U484 ( .A(w3[20]), .B(sa03_sr[4]), .Y(n449) );
  XOR2X1 U487 ( .A(n449), .B(n448), .Y(n446) );
  XOR2X1 U471 ( .A(sa13_sr[0]), .B(sa23_sr[0]), .Y(n459) );
  XOR2X1 U470 ( .A(w3[17]), .B(sa03_sr[1]), .Y(n460) );
  XOR2X1 U473 ( .A(n460), .B(n459), .Y(n457) );
  XOR2X1 U611 ( .A(sa12_sr[0]), .B(sa22_sr[0]), .Y(n369) );
  XOR2X1 U610 ( .A(w2[17]), .B(sa02_sr[1]), .Y(n370) );
  XOR2X1 U613 ( .A(n370), .B(n369), .Y(n367) );
  XOR2X1 U625 ( .A(sa12_sr[3]), .B(sa22_sr[3]), .Y(n358) );
  XOR2XL U624 ( .A(w2[20]), .B(sa02_sr[4]), .Y(n359) );
  XOR2X1 U627 ( .A(n359), .B(n358), .Y(n356) );
  XOR2X1 U891 ( .A(sa10_sr[0]), .B(sa20_sr[0]), .Y(n189) );
  XOR2X1 U890 ( .A(w0[17]), .B(sa00_sr[1]), .Y(n190) );
  XOR2X1 U893 ( .A(n190), .B(n189), .Y(n187) );
  XOR2X1 U905 ( .A(sa10_sr[3]), .B(sa20_sr[3]), .Y(n178) );
  XOR2XL U904 ( .A(w0[20]), .B(sa00_sr[4]), .Y(n179) );
  XOR2X1 U907 ( .A(n179), .B(n178), .Y(n176) );
  XOR2X1 U723 ( .A(w1[9]), .B(sa31_sr[1]), .Y(n299) );
  XOR2X1 U725 ( .A(n533), .B(n299), .Y(n297) );
  XOR2X1 U443 ( .A(w3[9]), .B(sa33_sr[1]), .Y(n479) );
  XOR2X1 U445 ( .A(n569), .B(n479), .Y(n477) );
  XOR2X1 U583 ( .A(w2[9]), .B(sa32_sr[1]), .Y(n389) );
  XOR2X1 U585 ( .A(n551), .B(n389), .Y(n387) );
  XOR2X1 U863 ( .A(w0[9]), .B(sa30_sr[1]), .Y(n209) );
  XOR2X1 U865 ( .A(n515), .B(n209), .Y(n207) );
  XOR2XL U698 ( .A(sa21_sr[3]), .B(sa31_sr[2]), .Y(n317) );
  XOR2XL U697 ( .A(w1[3]), .B(sa01_sr[2]), .Y(n318) );
  XOR2X1 U700 ( .A(n318), .B(n317), .Y(n315) );
  XOR2XL U734 ( .A(w1[12]), .B(sa31_sr[4]), .Y(n291) );
  XOR2X1 U736 ( .A(n530), .B(n291), .Y(n289) );
  XOR2XL U418 ( .A(sa23_sr[3]), .B(sa33_sr[2]), .Y(n497) );
  XOR2XL U417 ( .A(w3[3]), .B(sa03_sr[2]), .Y(n498) );
  XOR2X1 U420 ( .A(n498), .B(n497), .Y(n495) );
  XOR2XL U454 ( .A(w3[12]), .B(sa33_sr[4]), .Y(n471) );
  XOR2X1 U456 ( .A(n566), .B(n471), .Y(n469) );
  XOR2XL U558 ( .A(sa22_sr[3]), .B(sa32_sr[2]), .Y(n407) );
  XOR2XL U557 ( .A(w2[3]), .B(sa02_sr[2]), .Y(n408) );
  XOR2X1 U560 ( .A(n408), .B(n407), .Y(n405) );
  XOR2XL U594 ( .A(w2[12]), .B(sa32_sr[4]), .Y(n381) );
  XOR2X1 U596 ( .A(n548), .B(n381), .Y(n379) );
  XOR2XL U838 ( .A(sa20_sr[3]), .B(sa30_sr[2]), .Y(n227) );
  XOR2XL U837 ( .A(w0[3]), .B(sa00_sr[2]), .Y(n228) );
  XOR2X1 U840 ( .A(n228), .B(n227), .Y(n225) );
  XOR2XL U874 ( .A(w0[12]), .B(sa30_sr[4]), .Y(n201) );
  XOR2X1 U876 ( .A(n512), .B(n201), .Y(n199) );
  XOR2X1 U703 ( .A(sa21_sr[4]), .B(sa31_sr[3]), .Y(n313) );
  XOR2X1 U702 ( .A(w1[4]), .B(sa01_sr[3]), .Y(n314) );
  XOR2X1 U705 ( .A(n314), .B(n313), .Y(n311) );
  XOR2X1 U423 ( .A(sa23_sr[4]), .B(sa33_sr[3]), .Y(n493) );
  XOR2X1 U422 ( .A(w3[4]), .B(sa03_sr[3]), .Y(n494) );
  XOR2X1 U425 ( .A(n494), .B(n493), .Y(n491) );
  XOR2X1 U563 ( .A(sa22_sr[4]), .B(sa32_sr[3]), .Y(n403) );
  XOR2X1 U562 ( .A(w2[4]), .B(sa02_sr[3]), .Y(n404) );
  XOR2X1 U565 ( .A(n404), .B(n403), .Y(n401) );
  XOR2X1 U843 ( .A(sa20_sr[4]), .B(sa30_sr[3]), .Y(n223) );
  XOR2X1 U842 ( .A(w0[4]), .B(sa00_sr[3]), .Y(n224) );
  XOR2X1 U845 ( .A(n224), .B(n223), .Y(n221) );
  XOR2XL U760 ( .A(sa11_sr[2]), .B(sa21_sr[2]), .Y(n272) );
  XOR2X1 U759 ( .A(w1[19]), .B(sa01_sr[3]), .Y(n273) );
  XOR2X1 U762 ( .A(n273), .B(n272), .Y(n270) );
  XOR2XL U480 ( .A(sa13_sr[2]), .B(sa23_sr[2]), .Y(n452) );
  XOR2X1 U479 ( .A(w3[19]), .B(sa03_sr[3]), .Y(n453) );
  XOR2X1 U482 ( .A(n453), .B(n452), .Y(n450) );
  XOR2XL U620 ( .A(sa12_sr[2]), .B(sa22_sr[2]), .Y(n362) );
  XOR2X1 U619 ( .A(w2[19]), .B(sa02_sr[3]), .Y(n363) );
  XOR2X1 U622 ( .A(n363), .B(n362), .Y(n360) );
  XOR2XL U900 ( .A(sa10_sr[2]), .B(sa20_sr[2]), .Y(n182) );
  XOR2X1 U899 ( .A(w0[19]), .B(sa00_sr[3]), .Y(n183) );
  XOR2X1 U902 ( .A(n183), .B(n182), .Y(n180) );
  XOR2X1 U778 ( .A(w1[23]), .B(sa01_sr[7]), .Y(n259) );
  XOR2X1 U780 ( .A(n534), .B(n259), .Y(n257) );
  XOR2X1 U498 ( .A(w3[23]), .B(sa03_sr[7]), .Y(n439) );
  XOR2X1 U500 ( .A(n570), .B(n439), .Y(n437) );
  XOR2X1 U716 ( .A(w1[7]), .B(sa01_sr[6]), .Y(n304) );
  XOR2X1 U718 ( .A(n535), .B(n304), .Y(n302) );
  XOR2X1 U436 ( .A(w3[7]), .B(sa03_sr[6]), .Y(n484) );
  XOR2X1 U438 ( .A(n571), .B(n484), .Y(n482) );
  XOR2X1 U638 ( .A(w2[23]), .B(sa02_sr[7]), .Y(n349) );
  XOR2X1 U640 ( .A(n552), .B(n349), .Y(n347) );
  XOR2X1 U918 ( .A(w0[23]), .B(sa00_sr[7]), .Y(n169) );
  XOR2X1 U920 ( .A(n516), .B(n169), .Y(n167) );
  XOR2X1 U856 ( .A(w0[7]), .B(sa00_sr[6]), .Y(n214) );
  XOR2X1 U858 ( .A(n517), .B(n214), .Y(n212) );
  XOR2X1 U576 ( .A(w2[7]), .B(sa02_sr[6]), .Y(n394) );
  XOR2X1 U578 ( .A(n553), .B(n394), .Y(n392) );
  XOR2XL U803 ( .A(w1[28]), .B(sa11_sr[4]), .Y(n246) );
  XOR2X1 U805 ( .A(n529), .B(n246), .Y(n244) );
  XOR2XL U523 ( .A(w3[28]), .B(sa13_sr[4]), .Y(n426) );
  XOR2X1 U525 ( .A(n565), .B(n426), .Y(n424) );
  XOR2XL U663 ( .A(w2[28]), .B(sa12_sr[4]), .Y(n336) );
  XOR2X1 U665 ( .A(n547), .B(n336), .Y(n334) );
  XOR2XL U943 ( .A(w0[28]), .B(sa10_sr[4]), .Y(n156) );
  XOR2X1 U945 ( .A(n511), .B(n156), .Y(n154) );
  XOR2XL U792 ( .A(w1[26]), .B(sa11_sr[2]), .Y(n251) );
  XOR2XL U512 ( .A(w3[26]), .B(sa13_sr[2]), .Y(n431) );
  XOR2XL U652 ( .A(w2[26]), .B(sa12_sr[2]), .Y(n341) );
  XOR2XL U932 ( .A(w0[26]), .B(sa10_sr[2]), .Y(n161) );
  XOR2XL U727 ( .A(w1[10]), .B(sa31_sr[2]), .Y(n296) );
  XOR2XL U447 ( .A(w3[10]), .B(sa33_sr[2]), .Y(n476) );
  XOR2XL U587 ( .A(w2[10]), .B(sa32_sr[2]), .Y(n386) );
  XOR2XL U867 ( .A(w0[10]), .B(sa30_sr[2]), .Y(n206) );
  XOR2X1 U693 ( .A(w1[2]), .B(sa01_sr[1]), .Y(n321) );
  XOR2X1 U770 ( .A(w1[21]), .B(sa01_sr[5]), .Y(n265) );
  XOR2X1 U413 ( .A(w3[2]), .B(sa03_sr[1]), .Y(n501) );
  XOR2X1 U490 ( .A(w3[21]), .B(sa03_sr[5]), .Y(n445) );
  XOR2X1 U553 ( .A(w2[2]), .B(sa02_sr[1]), .Y(n411) );
  XOR2X1 U630 ( .A(w2[21]), .B(sa02_sr[5]), .Y(n355) );
  XOR2X1 U833 ( .A(w0[2]), .B(sa00_sr[1]), .Y(n231) );
  XOR2X1 U910 ( .A(w0[21]), .B(sa00_sr[5]), .Y(n175) );
  XOR2XL U708 ( .A(w1[5]), .B(sa01_sr[4]), .Y(n310) );
  XOR2XL U428 ( .A(w3[5]), .B(sa03_sr[4]), .Y(n490) );
  XOR2XL U568 ( .A(w2[5]), .B(sa02_sr[4]), .Y(n400) );
  XOR2XL U848 ( .A(w0[5]), .B(sa00_sr[4]), .Y(n220) );
  DFFHQX1 done_reg ( .D(N21), .CK(clk), .Q(done) );
  DFFHQX1 \text_out_reg[127]  ( .D(N376), .CK(clk), .Q(text_out[127]) );
  DFFHQX1 \text_out_reg[126]  ( .D(N377), .CK(clk), .Q(text_out[126]) );
  DFFHQX1 \text_out_reg[125]  ( .D(N378), .CK(clk), .Q(text_out[125]) );
  DFFHQX1 \text_out_reg[124]  ( .D(N379), .CK(clk), .Q(text_out[124]) );
  DFFHQX1 \text_out_reg[123]  ( .D(N380), .CK(clk), .Q(text_out[123]) );
  DFFHQX1 \text_out_reg[122]  ( .D(N381), .CK(clk), .Q(text_out[122]) );
  DFFHQX1 \text_out_reg[121]  ( .D(N382), .CK(clk), .Q(text_out[121]) );
  DFFHQX1 \text_out_reg[120]  ( .D(N383), .CK(clk), .Q(text_out[120]) );
  DFFHQX1 \text_out_reg[95]  ( .D(N384), .CK(clk), .Q(text_out[95]) );
  DFFHQX1 \text_out_reg[94]  ( .D(N385), .CK(clk), .Q(text_out[94]) );
  DFFHQX1 \text_out_reg[93]  ( .D(N386), .CK(clk), .Q(text_out[93]) );
  DFFHQX1 \text_out_reg[92]  ( .D(N387), .CK(clk), .Q(text_out[92]) );
  DFFHQX1 \text_out_reg[91]  ( .D(N388), .CK(clk), .Q(text_out[91]) );
  DFFHQX1 \text_out_reg[90]  ( .D(N389), .CK(clk), .Q(text_out[90]) );
  DFFHQX1 \text_out_reg[89]  ( .D(N390), .CK(clk), .Q(text_out[89]) );
  DFFHQX1 \text_out_reg[88]  ( .D(N391), .CK(clk), .Q(text_out[88]) );
  DFFHQX1 \text_out_reg[63]  ( .D(N392), .CK(clk), .Q(text_out[63]) );
  DFFHQX1 \text_out_reg[62]  ( .D(N393), .CK(clk), .Q(text_out[62]) );
  DFFHQX1 \text_out_reg[61]  ( .D(N394), .CK(clk), .Q(text_out[61]) );
  DFFHQX1 \text_out_reg[60]  ( .D(N395), .CK(clk), .Q(text_out[60]) );
  DFFHQX1 \text_out_reg[59]  ( .D(N396), .CK(clk), .Q(text_out[59]) );
  DFFHQX1 \text_out_reg[58]  ( .D(N397), .CK(clk), .Q(text_out[58]) );
  DFFHQX1 \text_out_reg[57]  ( .D(N398), .CK(clk), .Q(text_out[57]) );
  DFFHQX1 \text_out_reg[56]  ( .D(N399), .CK(clk), .Q(text_out[56]) );
  DFFHQX1 \text_out_reg[31]  ( .D(N400), .CK(clk), .Q(text_out[31]) );
  DFFHQX1 \text_out_reg[30]  ( .D(N401), .CK(clk), .Q(text_out[30]) );
  DFFHQX1 \text_out_reg[29]  ( .D(N402), .CK(clk), .Q(text_out[29]) );
  DFFHQX1 \text_out_reg[28]  ( .D(N403), .CK(clk), .Q(text_out[28]) );
  DFFHQX1 \text_out_reg[27]  ( .D(N404), .CK(clk), .Q(text_out[27]) );
  DFFHQX1 \text_out_reg[26]  ( .D(N405), .CK(clk), .Q(text_out[26]) );
  DFFHQX1 \text_out_reg[25]  ( .D(N406), .CK(clk), .Q(text_out[25]) );
  DFFHQX1 \text_out_reg[24]  ( .D(N407), .CK(clk), .Q(text_out[24]) );
  DFFHQX1 \text_out_reg[119]  ( .D(N408), .CK(clk), .Q(text_out[119]) );
  DFFHQX1 \text_out_reg[118]  ( .D(N409), .CK(clk), .Q(text_out[118]) );
  DFFHQX1 \text_out_reg[117]  ( .D(N410), .CK(clk), .Q(text_out[117]) );
  DFFHQX1 \text_out_reg[116]  ( .D(N411), .CK(clk), .Q(text_out[116]) );
  DFFHQX1 \text_out_reg[115]  ( .D(N412), .CK(clk), .Q(text_out[115]) );
  DFFHQX1 \text_out_reg[114]  ( .D(N413), .CK(clk), .Q(text_out[114]) );
  DFFHQX1 \text_out_reg[113]  ( .D(N414), .CK(clk), .Q(text_out[113]) );
  DFFHQX1 \text_out_reg[112]  ( .D(N415), .CK(clk), .Q(text_out[112]) );
  DFFHQX1 \text_out_reg[87]  ( .D(N416), .CK(clk), .Q(text_out[87]) );
  DFFHQX1 \text_out_reg[86]  ( .D(N417), .CK(clk), .Q(text_out[86]) );
  DFFHQX1 \text_out_reg[85]  ( .D(N418), .CK(clk), .Q(text_out[85]) );
  DFFHQX1 \text_out_reg[84]  ( .D(N419), .CK(clk), .Q(text_out[84]) );
  DFFHQX1 \text_out_reg[83]  ( .D(N420), .CK(clk), .Q(text_out[83]) );
  DFFHQX1 \text_out_reg[82]  ( .D(N421), .CK(clk), .Q(text_out[82]) );
  DFFHQX1 \text_out_reg[81]  ( .D(N422), .CK(clk), .Q(text_out[81]) );
  DFFHQX1 \text_out_reg[80]  ( .D(N423), .CK(clk), .Q(text_out[80]) );
  DFFHQX1 \text_out_reg[55]  ( .D(N424), .CK(clk), .Q(text_out[55]) );
  DFFHQX1 \text_out_reg[54]  ( .D(N425), .CK(clk), .Q(text_out[54]) );
  DFFHQX1 \text_out_reg[53]  ( .D(N426), .CK(clk), .Q(text_out[53]) );
  DFFHQX1 \text_out_reg[52]  ( .D(N427), .CK(clk), .Q(text_out[52]) );
  DFFHQX1 \text_out_reg[51]  ( .D(N428), .CK(clk), .Q(text_out[51]) );
  DFFHQX1 \text_out_reg[50]  ( .D(N429), .CK(clk), .Q(text_out[50]) );
  DFFHQX1 \text_out_reg[49]  ( .D(N430), .CK(clk), .Q(text_out[49]) );
  DFFHQX1 \text_out_reg[48]  ( .D(N431), .CK(clk), .Q(text_out[48]) );
  DFFHQX1 \text_out_reg[23]  ( .D(N432), .CK(clk), .Q(text_out[23]) );
  DFFHQX1 \text_out_reg[22]  ( .D(N433), .CK(clk), .Q(text_out[22]) );
  DFFHQX1 \text_out_reg[21]  ( .D(N434), .CK(clk), .Q(text_out[21]) );
  DFFHQX1 \text_out_reg[20]  ( .D(N435), .CK(clk), .Q(text_out[20]) );
  DFFHQX1 \text_out_reg[19]  ( .D(N436), .CK(clk), .Q(text_out[19]) );
  DFFHQX1 \text_out_reg[18]  ( .D(N437), .CK(clk), .Q(text_out[18]) );
  DFFHQX1 \text_out_reg[17]  ( .D(N438), .CK(clk), .Q(text_out[17]) );
  DFFHQX1 \text_out_reg[16]  ( .D(N439), .CK(clk), .Q(text_out[16]) );
  DFFHQX1 \text_out_reg[111]  ( .D(N440), .CK(clk), .Q(text_out[111]) );
  DFFHQX1 \text_out_reg[110]  ( .D(N441), .CK(clk), .Q(text_out[110]) );
  DFFHQX1 \text_out_reg[109]  ( .D(N442), .CK(clk), .Q(text_out[109]) );
  DFFHQX1 \text_out_reg[108]  ( .D(N443), .CK(clk), .Q(text_out[108]) );
  DFFHQX1 \text_out_reg[107]  ( .D(N444), .CK(clk), .Q(text_out[107]) );
  DFFHQX1 \text_out_reg[106]  ( .D(N445), .CK(clk), .Q(text_out[106]) );
  DFFHQX1 \text_out_reg[105]  ( .D(N446), .CK(clk), .Q(text_out[105]) );
  DFFHQX1 \text_out_reg[104]  ( .D(N447), .CK(clk), .Q(text_out[104]) );
  DFFHQX1 \text_out_reg[79]  ( .D(N448), .CK(clk), .Q(text_out[79]) );
  DFFHQX1 \text_out_reg[78]  ( .D(N449), .CK(clk), .Q(text_out[78]) );
  DFFHQX1 \text_out_reg[77]  ( .D(N450), .CK(clk), .Q(text_out[77]) );
  DFFHQX1 \text_out_reg[76]  ( .D(N451), .CK(clk), .Q(text_out[76]) );
  DFFHQX1 \text_out_reg[75]  ( .D(N452), .CK(clk), .Q(text_out[75]) );
  DFFHQX1 \text_out_reg[74]  ( .D(N453), .CK(clk), .Q(text_out[74]) );
  DFFHQX1 \text_out_reg[73]  ( .D(N454), .CK(clk), .Q(text_out[73]) );
  DFFHQX1 \text_out_reg[72]  ( .D(N455), .CK(clk), .Q(text_out[72]) );
  DFFHQX1 \text_out_reg[47]  ( .D(N456), .CK(clk), .Q(text_out[47]) );
  DFFHQX1 \text_out_reg[46]  ( .D(N457), .CK(clk), .Q(text_out[46]) );
  DFFHQX1 \text_out_reg[45]  ( .D(N458), .CK(clk), .Q(text_out[45]) );
  DFFHQX1 \text_out_reg[44]  ( .D(N459), .CK(clk), .Q(text_out[44]) );
  DFFHQX1 \text_out_reg[43]  ( .D(N460), .CK(clk), .Q(text_out[43]) );
  DFFHQX1 \text_out_reg[42]  ( .D(N461), .CK(clk), .Q(text_out[42]) );
  DFFHQX1 \text_out_reg[41]  ( .D(N462), .CK(clk), .Q(text_out[41]) );
  DFFHQX1 \text_out_reg[40]  ( .D(N463), .CK(clk), .Q(text_out[40]) );
  DFFHQX1 \text_out_reg[15]  ( .D(N464), .CK(clk), .Q(text_out[15]) );
  DFFHQX1 \text_out_reg[14]  ( .D(N465), .CK(clk), .Q(text_out[14]) );
  DFFHQX1 \text_out_reg[13]  ( .D(N466), .CK(clk), .Q(text_out[13]) );
  DFFHQX1 \text_out_reg[12]  ( .D(N467), .CK(clk), .Q(text_out[12]) );
  DFFHQX1 \text_out_reg[11]  ( .D(N468), .CK(clk), .Q(text_out[11]) );
  DFFHQX1 \text_out_reg[10]  ( .D(N469), .CK(clk), .Q(text_out[10]) );
  DFFHQX1 \text_out_reg[9]  ( .D(N470), .CK(clk), .Q(text_out[9]) );
  DFFHQX1 \text_out_reg[8]  ( .D(N471), .CK(clk), .Q(text_out[8]) );
  DFFHQX1 \text_out_reg[103]  ( .D(N472), .CK(clk), .Q(text_out[103]) );
  DFFHQX1 \text_out_reg[102]  ( .D(N473), .CK(clk), .Q(text_out[102]) );
  DFFHQX1 \text_out_reg[101]  ( .D(N474), .CK(clk), .Q(text_out[101]) );
  DFFHQX1 \text_out_reg[100]  ( .D(N475), .CK(clk), .Q(text_out[100]) );
  DFFHQX1 \text_out_reg[99]  ( .D(N476), .CK(clk), .Q(text_out[99]) );
  DFFHQX1 \text_out_reg[98]  ( .D(N477), .CK(clk), .Q(text_out[98]) );
  DFFHQX1 \text_out_reg[97]  ( .D(N478), .CK(clk), .Q(text_out[97]) );
  DFFHQX1 \text_out_reg[96]  ( .D(N479), .CK(clk), .Q(text_out[96]) );
  DFFHQX1 \text_out_reg[71]  ( .D(N480), .CK(clk), .Q(text_out[71]) );
  DFFHQX1 \text_out_reg[70]  ( .D(N481), .CK(clk), .Q(text_out[70]) );
  DFFHQX1 \text_out_reg[69]  ( .D(N482), .CK(clk), .Q(text_out[69]) );
  DFFHQX1 \text_out_reg[68]  ( .D(N483), .CK(clk), .Q(text_out[68]) );
  DFFHQX1 \text_out_reg[67]  ( .D(N484), .CK(clk), .Q(text_out[67]) );
  DFFHQX1 \text_out_reg[66]  ( .D(N485), .CK(clk), .Q(text_out[66]) );
  DFFHQX1 \text_out_reg[65]  ( .D(N486), .CK(clk), .Q(text_out[65]) );
  DFFHQX1 \text_out_reg[64]  ( .D(N487), .CK(clk), .Q(text_out[64]) );
  DFFHQX1 \text_out_reg[39]  ( .D(N488), .CK(clk), .Q(text_out[39]) );
  DFFHQX1 \text_out_reg[38]  ( .D(N489), .CK(clk), .Q(text_out[38]) );
  DFFHQX1 \text_out_reg[37]  ( .D(N490), .CK(clk), .Q(text_out[37]) );
  DFFHQX1 \text_out_reg[36]  ( .D(N491), .CK(clk), .Q(text_out[36]) );
  DFFHQX1 \text_out_reg[35]  ( .D(N492), .CK(clk), .Q(text_out[35]) );
  DFFHQX1 \text_out_reg[34]  ( .D(N493), .CK(clk), .Q(text_out[34]) );
  DFFHQX1 \text_out_reg[33]  ( .D(N494), .CK(clk), .Q(text_out[33]) );
  DFFHQX1 \text_out_reg[32]  ( .D(N495), .CK(clk), .Q(text_out[32]) );
  DFFHQX1 \text_out_reg[7]  ( .D(N496), .CK(clk), .Q(text_out[7]) );
  DFFHQX1 \text_out_reg[6]  ( .D(N497), .CK(clk), .Q(text_out[6]) );
  DFFHQX1 \text_out_reg[5]  ( .D(N498), .CK(clk), .Q(text_out[5]) );
  DFFHQX1 \text_out_reg[4]  ( .D(N499), .CK(clk), .Q(text_out[4]) );
  DFFHQX1 \text_out_reg[3]  ( .D(N500), .CK(clk), .Q(text_out[3]) );
  DFFHQX1 \text_out_reg[2]  ( .D(N501), .CK(clk), .Q(text_out[2]) );
  DFFHQX1 \text_out_reg[1]  ( .D(N502), .CK(clk), .Q(text_out[1]) );
  DFFHQX1 \text_out_reg[0]  ( .D(N503), .CK(clk), .Q(text_out[0]) );
  XOR2X1 U694 ( .A(sa21_sr[2]), .B(sa31_sr[1]), .Y(n320) );
  XOR2X1 U414 ( .A(sa23_sr[2]), .B(sa33_sr[1]), .Y(n500) );
  XOR2X1 U554 ( .A(sa22_sr[2]), .B(sa32_sr[1]), .Y(n410) );
  XOR2X1 U834 ( .A(sa20_sr[2]), .B(sa30_sr[1]), .Y(n230) );
  XOR2XL U709 ( .A(sa21_sr[5]), .B(sa31_sr[4]), .Y(n309) );
  XOR2XL U429 ( .A(sa23_sr[5]), .B(sa33_sr[4]), .Y(n489) );
  XOR2XL U569 ( .A(sa22_sr[5]), .B(sa32_sr[4]), .Y(n399) );
  XOR2XL U849 ( .A(sa20_sr[5]), .B(sa30_sr[4]), .Y(n219) );
  XOR2XL U771 ( .A(sa11_sr[4]), .B(sa21_sr[4]), .Y(n264) );
  XOR2XL U491 ( .A(sa13_sr[4]), .B(sa23_sr[4]), .Y(n444) );
  XOR2XL U631 ( .A(sa12_sr[4]), .B(sa22_sr[4]), .Y(n354) );
  XOR2XL U911 ( .A(sa10_sr[4]), .B(sa20_sr[4]), .Y(n174) );
  XOR2X1 U819 ( .A(sa01_sr[5]), .B(sa11_sr[5]), .Y(n537) );
  XOR2X1 U539 ( .A(sa03_sr[5]), .B(sa13_sr[5]), .Y(n573) );
  XOR2X1 U679 ( .A(sa02_sr[5]), .B(sa12_sr[5]), .Y(n555) );
  XOR2X1 U959 ( .A(sa00_sr[5]), .B(sa10_sr[5]), .Y(n519) );
  XOR2X1 U847 ( .A(sa00_sr[7]), .B(sa30_sr[7]), .Y(n525) );
  XOR2X1 U707 ( .A(sa01_sr[7]), .B(sa31_sr[7]), .Y(n543) );
  XOR2X1 U567 ( .A(sa02_sr[7]), .B(sa32_sr[7]), .Y(n561) );
  XOR2X1 U427 ( .A(sa03_sr[7]), .B(sa33_sr[7]), .Y(n579) );
  XOR2X1 U629 ( .A(sa12_sr[7]), .B(sa22_sr[7]), .Y(n544) );
  XOR2X1 U769 ( .A(sa11_sr[7]), .B(sa21_sr[7]), .Y(n526) );
  XOR2X1 U909 ( .A(sa10_sr[7]), .B(sa20_sr[7]), .Y(n508) );
  XOR2X1 U489 ( .A(sa13_sr[7]), .B(sa23_sr[7]), .Y(n562) );
  XOR2X1 U801 ( .A(sa21_sr[3]), .B(sa31_sr[3]), .Y(n530) );
  XOR2X1 U521 ( .A(sa23_sr[3]), .B(sa33_sr[3]), .Y(n566) );
  XOR2X1 U661 ( .A(sa22_sr[3]), .B(sa32_sr[3]), .Y(n548) );
  XOR2X1 U941 ( .A(sa20_sr[3]), .B(sa30_sr[3]), .Y(n512) );
  XOR2X1 U823 ( .A(sa01_sr[6]), .B(sa11_sr[6]), .Y(n536) );
  XOR2X1 U543 ( .A(sa03_sr[6]), .B(sa13_sr[6]), .Y(n572) );
  XOR2X1 U683 ( .A(sa02_sr[6]), .B(sa12_sr[6]), .Y(n554) );
  XOR2X1 U963 ( .A(sa00_sr[6]), .B(sa10_sr[6]), .Y(n518) );
  XOR2X1 U795 ( .A(sa21_sr[2]), .B(sa31_sr[2]), .Y(n531) );
  XOR2X1 U515 ( .A(sa23_sr[2]), .B(sa33_sr[2]), .Y(n567) );
  XOR2X1 U655 ( .A(sa22_sr[2]), .B(sa32_sr[2]), .Y(n549) );
  XOR2X1 U935 ( .A(sa20_sr[2]), .B(sa30_sr[2]), .Y(n513) );
  XOR2XL U802 ( .A(sa01_sr[2]), .B(sa11_sr[2]), .Y(n540) );
  XOR2XL U522 ( .A(sa03_sr[2]), .B(sa13_sr[2]), .Y(n576) );
  XOR2XL U662 ( .A(sa02_sr[2]), .B(sa12_sr[2]), .Y(n558) );
  XOR2XL U942 ( .A(sa00_sr[2]), .B(sa10_sr[2]), .Y(n522) );
  XOR2X1 U958 ( .A(sa20_sr[6]), .B(sa30_sr[6]), .Y(n509) );
  XOR2X1 U538 ( .A(sa23_sr[6]), .B(sa33_sr[6]), .Y(n563) );
  XOR2X1 U790 ( .A(sa21_sr[1]), .B(sa31_sr[1]), .Y(n532) );
  XOR2X1 U813 ( .A(sa21_sr[5]), .B(sa31_sr[5]), .Y(n528) );
  XOR2X1 U818 ( .A(sa21_sr[6]), .B(sa31_sr[6]), .Y(n527) );
  XOR2X1 U510 ( .A(sa23_sr[1]), .B(sa33_sr[1]), .Y(n568) );
  XOR2X1 U533 ( .A(sa23_sr[5]), .B(sa33_sr[5]), .Y(n564) );
  XOR2X1 U650 ( .A(sa22_sr[1]), .B(sa32_sr[1]), .Y(n550) );
  XOR2X1 U673 ( .A(sa22_sr[5]), .B(sa32_sr[5]), .Y(n546) );
  XOR2X1 U678 ( .A(sa22_sr[6]), .B(sa32_sr[6]), .Y(n545) );
  XOR2X1 U930 ( .A(sa20_sr[1]), .B(sa30_sr[1]), .Y(n514) );
  XOR2X1 U953 ( .A(sa20_sr[5]), .B(sa30_sr[5]), .Y(n510) );
  XOR2X1 U796 ( .A(sa01_sr[1]), .B(sa11_sr[1]), .Y(n541) );
  XOR2X1 U516 ( .A(sa03_sr[1]), .B(sa13_sr[1]), .Y(n577) );
  XOR2X1 U656 ( .A(sa02_sr[1]), .B(sa12_sr[1]), .Y(n559) );
  XOR2X1 U936 ( .A(sa00_sr[1]), .B(sa10_sr[1]), .Y(n523) );
  XOR2X1 U925 ( .A(sa20_sr[0]), .B(sa30_sr[0]), .Y(n515) );
  XOR2X1 U645 ( .A(sa22_sr[0]), .B(sa32_sr[0]), .Y(n551) );
  XOR2X1 U785 ( .A(sa21_sr[0]), .B(sa31_sr[0]), .Y(n533) );
  XOR2X1 U505 ( .A(sa23_sr[0]), .B(sa33_sr[0]), .Y(n569) );
  XOR2X1 U949 ( .A(sa00_sr[7]), .B(sa10_sr[7]), .Y(n517) );
  XOR2X1 U529 ( .A(sa03_sr[7]), .B(sa13_sr[7]), .Y(n571) );
  XOR2X1 U824 ( .A(sa21_sr[7]), .B(sa31_sr[7]), .Y(n534) );
  XOR2X1 U809 ( .A(sa01_sr[7]), .B(sa11_sr[7]), .Y(n535) );
  XOR2X1 U544 ( .A(sa23_sr[7]), .B(sa33_sr[7]), .Y(n570) );
  XOR2X1 U669 ( .A(sa02_sr[7]), .B(sa12_sr[7]), .Y(n553) );
  XOR2X1 U684 ( .A(sa22_sr[7]), .B(sa32_sr[7]), .Y(n552) );
  XOR2X1 U964 ( .A(sa20_sr[7]), .B(sa30_sr[7]), .Y(n516) );
  XOR2X1 U807 ( .A(sa21_sr[4]), .B(sa31_sr[4]), .Y(n529) );
  XOR2X1 U527 ( .A(sa23_sr[4]), .B(sa33_sr[4]), .Y(n565) );
  XOR2X1 U667 ( .A(sa22_sr[4]), .B(sa32_sr[4]), .Y(n547) );
  XOR2X1 U947 ( .A(sa20_sr[4]), .B(sa30_sr[4]), .Y(n511) );
  XOR2XL U814 ( .A(sa01_sr[4]), .B(sa11_sr[4]), .Y(n538) );
  XOR2XL U534 ( .A(sa03_sr[4]), .B(sa13_sr[4]), .Y(n574) );
  XOR2XL U674 ( .A(sa02_sr[4]), .B(sa12_sr[4]), .Y(n556) );
  XOR2XL U954 ( .A(sa00_sr[4]), .B(sa10_sr[4]), .Y(n520) );
  XOR2X1 U931 ( .A(sa00_sr[0]), .B(sa10_sr[0]), .Y(n524) );
  XOR2X1 U791 ( .A(sa01_sr[0]), .B(sa11_sr[0]), .Y(n542) );
  XOR2X1 U651 ( .A(sa02_sr[0]), .B(sa12_sr[0]), .Y(n560) );
  XOR2X1 U511 ( .A(sa03_sr[0]), .B(sa13_sr[0]), .Y(n578) );
  XOR2X1 U808 ( .A(sa01_sr[3]), .B(sa11_sr[3]), .Y(n539) );
  XOR2X1 U528 ( .A(sa03_sr[3]), .B(sa13_sr[3]), .Y(n575) );
  XOR2X1 U668 ( .A(sa02_sr[3]), .B(sa12_sr[3]), .Y(n557) );
  XOR2X1 U948 ( .A(sa00_sr[3]), .B(sa10_sr[3]), .Y(n521) );
  XOR2X1 U821 ( .A(n534), .B(n536), .Y(n238) );
  XOR2X1 U541 ( .A(n570), .B(n572), .Y(n418) );
  XOR2X1 U681 ( .A(n552), .B(n554), .Y(n328) );
  XOR2X1 U961 ( .A(n516), .B(n518), .Y(n148) );
  XOR2X1 U885 ( .A(n517), .B(n509), .Y(n193) );
  XOR2X1 U465 ( .A(n571), .B(n563), .Y(n463) );
  XOR2X1 U816 ( .A(n537), .B(n527), .Y(n240) );
  XOR2X1 U742 ( .A(n536), .B(n528), .Y(n285) );
  XOR2X1 U745 ( .A(n535), .B(n527), .Y(n283) );
  XOR2X1 U536 ( .A(n573), .B(n563), .Y(n420) );
  XOR2X1 U462 ( .A(n572), .B(n564), .Y(n465) );
  XOR2X1 U676 ( .A(n555), .B(n545), .Y(n330) );
  XOR2X1 U602 ( .A(n554), .B(n546), .Y(n375) );
  XOR2X1 U605 ( .A(n553), .B(n545), .Y(n373) );
  XOR2X1 U882 ( .A(n518), .B(n510), .Y(n195) );
  XOR2X1 U956 ( .A(n519), .B(n509), .Y(n150) );
  XOR2X1 U923 ( .A(n517), .B(n515), .Y(n165) );
  XOR2X1 U608 ( .A(n544), .B(n551), .Y(n371) );
  XOR2X1 U748 ( .A(n526), .B(n533), .Y(n281) );
  XOR2X1 U888 ( .A(n508), .B(n515), .Y(n191) );
  XOR2X1 U783 ( .A(n535), .B(n533), .Y(n255) );
  XOR2X1 U503 ( .A(n571), .B(n569), .Y(n435) );
  XOR2X1 U468 ( .A(n562), .B(n569), .Y(n461) );
  XOR2X1 U643 ( .A(n553), .B(n551), .Y(n345) );
  XOR2X1 U739 ( .A(n537), .B(n529), .Y(n287) );
  XOR2X1 U459 ( .A(n573), .B(n565), .Y(n467) );
  XOR2X1 U599 ( .A(n555), .B(n547), .Y(n377) );
  XOR2X1 U879 ( .A(n519), .B(n511), .Y(n197) );
  XOR2X1 U826 ( .A(n525), .B(n524), .Y(n236) );
  XOR2X1 U686 ( .A(n543), .B(n542), .Y(n326) );
  XOR2X1 U546 ( .A(n561), .B(n560), .Y(n416) );
  XOR2X1 U406 ( .A(n579), .B(n578), .Y(n506) );
  XOR2X1 U721 ( .A(n534), .B(n542), .Y(n300) );
  XOR2X1 U441 ( .A(n570), .B(n578), .Y(n480) );
  XOR2X1 U581 ( .A(n552), .B(n560), .Y(n390) );
  XOR2X1 U861 ( .A(n516), .B(n524), .Y(n210) );
  XOR2X1 U811 ( .A(n538), .B(n528), .Y(n242) );
  XOR2X1 U531 ( .A(n574), .B(n564), .Y(n422) );
  XOR2X1 U671 ( .A(n556), .B(n546), .Y(n332) );
  XOR2X1 U951 ( .A(n520), .B(n510), .Y(n152) );
  DFFHQX2 \sa00_reg[1]  ( .D(N273), .CK(clk), .Q(sa00[1]) );
  DFFHQX2 \sa01_reg[1]  ( .D(N209), .CK(clk), .Q(sa01[1]) );
  DFFHQX2 \sa02_reg[1]  ( .D(N145), .CK(clk), .Q(sa02[1]) );
  DFFHQX2 \sa03_reg[1]  ( .D(N81), .CK(clk), .Q(sa03[1]) );
  DFFHQX2 \sa10_reg[1]  ( .D(N257), .CK(clk), .Q(sa10[1]) );
  DFFHQX2 \sa11_reg[1]  ( .D(N193), .CK(clk), .Q(sa11[1]) );
  DFFHQX2 \sa12_reg[1]  ( .D(N129), .CK(clk), .Q(sa12[1]) );
  DFFHQX2 \sa13_reg[1]  ( .D(N65), .CK(clk), .Q(sa13[1]) );
  DFFHQX2 \sa20_reg[1]  ( .D(N241), .CK(clk), .Q(sa20[1]) );
  DFFHQX2 \sa21_reg[1]  ( .D(N177), .CK(clk), .Q(sa21[1]) );
  DFFHQX2 \sa22_reg[1]  ( .D(N113), .CK(clk), .Q(sa22[1]) );
  DFFHQX2 \sa23_reg[1]  ( .D(N49), .CK(clk), .Q(sa23[1]) );
  DFFHQX2 \sa30_reg[1]  ( .D(N225), .CK(clk), .Q(sa30[1]) );
  DFFHQX2 \sa31_reg[1]  ( .D(N161), .CK(clk), .Q(sa31[1]) );
  DFFHQX2 \sa32_reg[1]  ( .D(N97), .CK(clk), .Q(sa32[1]) );
  DFFHQX2 \sa33_reg[1]  ( .D(N33), .CK(clk), .Q(sa33[1]) );
  CLKINVX3 U965 ( .A(n590), .Y(n582) );
  CLKINVX3 U966 ( .A(n580), .Y(n587) );
  CLKINVX3 U967 ( .A(n589), .Y(n585) );
  CLKINVX3 U968 ( .A(n589), .Y(n583) );
  CLKINVX3 U969 ( .A(n590), .Y(n581) );
  CLKINVX3 U970 ( .A(n590), .Y(n588) );
  CLKINVX3 U971 ( .A(n580), .Y(n586) );
  CLKINVX3 U972 ( .A(n589), .Y(n584) );
  INVX1 U973 ( .A(n731), .Y(n590) );
  INVX1 U974 ( .A(n731), .Y(n589) );
  OAI21XL U975 ( .A0(dcnt[0]), .A1(n591), .B0(n592), .Y(n147) );
  OAI21XL U976 ( .A0(n593), .A1(n591), .B0(n592), .Y(n146) );
  AOI21X1 U977 ( .A0(dcnt[1]), .A1(dcnt[0]), .B0(n594), .Y(n593) );
  AOI21X1 U978 ( .A0(n595), .A1(n596), .B0(n591), .Y(n145) );
  NAND2X1 U979 ( .A(n730), .B(n597), .Y(n596) );
  OAI31X1 U980 ( .A0(n598), .A1(n599), .A2(n591), .B0(n592), .Y(n1) );
  NAND2X1 U981 ( .A(ld), .B(rst), .Y(n592) );
  OAI211X1 U982 ( .A0(dcnt[3]), .A1(n595), .B0(n600), .C0(rst), .Y(n591) );
  INVX1 U983 ( .A(ld), .Y(n600) );
  INVX1 U984 ( .A(n599), .Y(n595) );
  NOR2X1 U985 ( .A(n597), .B(n730), .Y(n599) );
  INVX1 U986 ( .A(n594), .Y(n597) );
  NOR2X1 U987 ( .A(dcnt[1]), .B(dcnt[0]), .Y(n594) );
  INVX1 U988 ( .A(dcnt[3]), .Y(n598) );
  MX2X1 U989 ( .A(sa32_next[3]), .B(n601), .S0(n581), .Y(N99) );
  XOR2X1 U990 ( .A(w2[3]), .B(text_in_r[35]), .Y(n601) );
  MX2X1 U991 ( .A(sa32_next[2]), .B(n602), .S0(n581), .Y(N98) );
  XOR2X1 U992 ( .A(w2[2]), .B(text_in_r[34]), .Y(n602) );
  MX2X1 U993 ( .A(sa32_next[1]), .B(n603), .S0(n581), .Y(N97) );
  XOR2X1 U994 ( .A(w2[1]), .B(text_in_r[33]), .Y(n603) );
  MX2X1 U995 ( .A(sa32_next[0]), .B(n604), .S0(n581), .Y(N96) );
  XOR2X1 U996 ( .A(w2[0]), .B(text_in_r[32]), .Y(n604) );
  MX2X1 U997 ( .A(sa03_next[7]), .B(n605), .S0(n581), .Y(N87) );
  XOR2X1 U998 ( .A(w3[31]), .B(text_in_r[31]), .Y(n605) );
  MX2X1 U999 ( .A(sa03_next[6]), .B(n606), .S0(n581), .Y(N86) );
  XOR2X1 U1000 ( .A(w3[30]), .B(text_in_r[30]), .Y(n606) );
  MX2X1 U1001 ( .A(sa03_next[5]), .B(n607), .S0(n581), .Y(N85) );
  XOR2X1 U1002 ( .A(w3[29]), .B(text_in_r[29]), .Y(n607) );
  MX2X1 U1003 ( .A(sa03_next[4]), .B(n608), .S0(n581), .Y(N84) );
  XOR2X1 U1004 ( .A(w3[28]), .B(text_in_r[28]), .Y(n608) );
  MX2X1 U1005 ( .A(sa03_next[3]), .B(n609), .S0(n581), .Y(N83) );
  XOR2X1 U1006 ( .A(w3[27]), .B(text_in_r[27]), .Y(n609) );
  MX2X1 U1007 ( .A(sa03_next[2]), .B(n610), .S0(n581), .Y(N82) );
  XOR2X1 U1008 ( .A(w3[26]), .B(text_in_r[26]), .Y(n610) );
  MX2X1 U1009 ( .A(sa03_next[1]), .B(n611), .S0(n581), .Y(N81) );
  XOR2X1 U1010 ( .A(w3[25]), .B(text_in_r[25]), .Y(n611) );
  MX2X1 U1011 ( .A(sa03_next[0]), .B(n612), .S0(n581), .Y(N80) );
  XOR2X1 U1012 ( .A(w3[24]), .B(text_in_r[24]), .Y(n612) );
  MX2X1 U1013 ( .A(sa13_next[7]), .B(n613), .S0(n581), .Y(N71) );
  XOR2X1 U1014 ( .A(w3[23]), .B(text_in_r[23]), .Y(n613) );
  MX2X1 U1015 ( .A(sa13_next[6]), .B(n614), .S0(n582), .Y(N70) );
  XOR2X1 U1016 ( .A(w3[22]), .B(text_in_r[22]), .Y(n614) );
  MX2X1 U1017 ( .A(sa13_next[5]), .B(n615), .S0(n582), .Y(N69) );
  XOR2X1 U1018 ( .A(w3[21]), .B(text_in_r[21]), .Y(n615) );
  MX2X1 U1019 ( .A(sa13_next[4]), .B(n616), .S0(n582), .Y(N68) );
  XOR2X1 U1020 ( .A(w3[20]), .B(text_in_r[20]), .Y(n616) );
  MX2X1 U1021 ( .A(sa13_next[3]), .B(n617), .S0(n582), .Y(N67) );
  XOR2X1 U1022 ( .A(w3[19]), .B(text_in_r[19]), .Y(n617) );
  MX2X1 U1023 ( .A(sa13_next[2]), .B(n618), .S0(n582), .Y(N66) );
  XOR2X1 U1024 ( .A(w3[18]), .B(text_in_r[18]), .Y(n618) );
  MX2X1 U1025 ( .A(sa13_next[1]), .B(n619), .S0(n582), .Y(N65) );
  XOR2X1 U1026 ( .A(w3[17]), .B(text_in_r[17]), .Y(n619) );
  MX2X1 U1027 ( .A(sa13_next[0]), .B(n620), .S0(n582), .Y(N64) );
  XOR2X1 U1028 ( .A(w3[16]), .B(text_in_r[16]), .Y(n620) );
  MX2X1 U1029 ( .A(sa23_next[7]), .B(n621), .S0(n582), .Y(N55) );
  XOR2X1 U1030 ( .A(w3[15]), .B(text_in_r[15]), .Y(n621) );
  MX2X1 U1031 ( .A(sa23_next[6]), .B(n622), .S0(n582), .Y(N54) );
  XOR2X1 U1032 ( .A(w3[14]), .B(text_in_r[14]), .Y(n622) );
  MX2X1 U1033 ( .A(sa23_next[5]), .B(n623), .S0(n582), .Y(N53) );
  XOR2X1 U1034 ( .A(w3[13]), .B(text_in_r[13]), .Y(n623) );
  MX2X1 U1035 ( .A(sa23_next[4]), .B(n624), .S0(n582), .Y(N52) );
  XOR2X1 U1036 ( .A(w3[12]), .B(text_in_r[12]), .Y(n624) );
  MX2X1 U1037 ( .A(sa23_next[3]), .B(n625), .S0(n582), .Y(N51) );
  XOR2X1 U1038 ( .A(w3[11]), .B(text_in_r[11]), .Y(n625) );
  XOR2X1 U1039 ( .A(w3[0]), .B(sa33_sr[0]), .Y(N503) );
  XOR2X1 U1040 ( .A(w3[1]), .B(sa33_sr[1]), .Y(N502) );
  XOR2X1 U1041 ( .A(w3[2]), .B(sa33_sr[2]), .Y(N501) );
  XOR2X1 U1042 ( .A(w3[3]), .B(sa33_sr[3]), .Y(N500) );
  MX2X1 U1043 ( .A(sa23_next[2]), .B(n626), .S0(n582), .Y(N50) );
  XOR2X1 U1044 ( .A(w3[10]), .B(text_in_r[10]), .Y(n626) );
  XOR2X1 U1045 ( .A(w3[4]), .B(sa33_sr[4]), .Y(N499) );
  XOR2X1 U1046 ( .A(w3[5]), .B(sa33_sr[5]), .Y(N498) );
  XOR2X1 U1047 ( .A(w3[6]), .B(sa33_sr[6]), .Y(N497) );
  XOR2X1 U1048 ( .A(w3[7]), .B(sa33_sr[7]), .Y(N496) );
  XOR2X1 U1049 ( .A(w2[0]), .B(sa32_sr[0]), .Y(N495) );
  XOR2X1 U1050 ( .A(w2[1]), .B(sa32_sr[1]), .Y(N494) );
  XOR2X1 U1051 ( .A(w2[2]), .B(sa32_sr[2]), .Y(N493) );
  XOR2X1 U1052 ( .A(w2[3]), .B(sa32_sr[3]), .Y(N492) );
  XOR2X1 U1053 ( .A(w2[4]), .B(sa32_sr[4]), .Y(N491) );
  XOR2X1 U1054 ( .A(w2[5]), .B(sa32_sr[5]), .Y(N490) );
  MX2X1 U1055 ( .A(sa23_next[1]), .B(n627), .S0(n583), .Y(N49) );
  XOR2X1 U1056 ( .A(w3[9]), .B(text_in_r[9]), .Y(n627) );
  XOR2X1 U1057 ( .A(w2[6]), .B(sa32_sr[6]), .Y(N489) );
  XOR2X1 U1058 ( .A(w2[7]), .B(sa32_sr[7]), .Y(N488) );
  XOR2X1 U1059 ( .A(w1[0]), .B(sa31_sr[0]), .Y(N487) );
  XOR2X1 U1060 ( .A(w1[1]), .B(sa31_sr[1]), .Y(N486) );
  XOR2X1 U1061 ( .A(w1[2]), .B(sa31_sr[2]), .Y(N485) );
  XOR2X1 U1062 ( .A(w1[3]), .B(sa31_sr[3]), .Y(N484) );
  XOR2X1 U1063 ( .A(w1[4]), .B(sa31_sr[4]), .Y(N483) );
  XOR2X1 U1064 ( .A(w1[5]), .B(sa31_sr[5]), .Y(N482) );
  XOR2X1 U1065 ( .A(w1[6]), .B(sa31_sr[6]), .Y(N481) );
  XOR2X1 U1066 ( .A(w1[7]), .B(sa31_sr[7]), .Y(N480) );
  MX2X1 U1067 ( .A(sa23_next[0]), .B(n628), .S0(n583), .Y(N48) );
  XOR2X1 U1068 ( .A(w3[8]), .B(text_in_r[8]), .Y(n628) );
  XOR2X1 U1069 ( .A(w0[0]), .B(sa30_sr[0]), .Y(N479) );
  XOR2X1 U1070 ( .A(w0[1]), .B(sa30_sr[1]), .Y(N478) );
  XOR2X1 U1071 ( .A(w0[2]), .B(sa30_sr[2]), .Y(N477) );
  XOR2X1 U1072 ( .A(w0[3]), .B(sa30_sr[3]), .Y(N476) );
  XOR2X1 U1073 ( .A(w0[4]), .B(sa30_sr[4]), .Y(N475) );
  XOR2X1 U1074 ( .A(w0[5]), .B(sa30_sr[5]), .Y(N474) );
  XOR2X1 U1075 ( .A(w0[6]), .B(sa30_sr[6]), .Y(N473) );
  XOR2X1 U1076 ( .A(w0[7]), .B(sa30_sr[7]), .Y(N472) );
  XOR2X1 U1077 ( .A(w3[8]), .B(sa23_sr[0]), .Y(N471) );
  XOR2X1 U1078 ( .A(w3[9]), .B(sa23_sr[1]), .Y(N470) );
  XOR2X1 U1079 ( .A(w3[10]), .B(sa23_sr[2]), .Y(N469) );
  XOR2X1 U1080 ( .A(w3[11]), .B(sa23_sr[3]), .Y(N468) );
  XOR2X1 U1081 ( .A(w3[12]), .B(sa23_sr[4]), .Y(N467) );
  XOR2X1 U1082 ( .A(w3[13]), .B(sa23_sr[5]), .Y(N466) );
  XOR2X1 U1083 ( .A(w3[14]), .B(sa23_sr[6]), .Y(N465) );
  XOR2X1 U1084 ( .A(w3[15]), .B(sa23_sr[7]), .Y(N464) );
  XOR2X1 U1085 ( .A(w2[8]), .B(sa22_sr[0]), .Y(N463) );
  XOR2X1 U1086 ( .A(w2[9]), .B(sa22_sr[1]), .Y(N462) );
  XOR2X1 U1087 ( .A(w2[10]), .B(sa22_sr[2]), .Y(N461) );
  XOR2X1 U1088 ( .A(w2[11]), .B(sa22_sr[3]), .Y(N460) );
  XOR2X1 U1089 ( .A(w2[12]), .B(sa22_sr[4]), .Y(N459) );
  XOR2X1 U1090 ( .A(w2[13]), .B(sa22_sr[5]), .Y(N458) );
  XOR2X1 U1091 ( .A(w2[14]), .B(sa22_sr[6]), .Y(N457) );
  XOR2X1 U1092 ( .A(w2[15]), .B(sa22_sr[7]), .Y(N456) );
  XOR2X1 U1093 ( .A(w1[8]), .B(sa21_sr[0]), .Y(N455) );
  XOR2X1 U1094 ( .A(w1[9]), .B(sa21_sr[1]), .Y(N454) );
  XOR2X1 U1095 ( .A(w1[10]), .B(sa21_sr[2]), .Y(N453) );
  XOR2X1 U1096 ( .A(w1[11]), .B(sa21_sr[3]), .Y(N452) );
  XOR2X1 U1097 ( .A(w1[12]), .B(sa21_sr[4]), .Y(N451) );
  XOR2X1 U1098 ( .A(w1[13]), .B(sa21_sr[5]), .Y(N450) );
  XOR2X1 U1099 ( .A(w1[14]), .B(sa21_sr[6]), .Y(N449) );
  XOR2X1 U1100 ( .A(w1[15]), .B(sa21_sr[7]), .Y(N448) );
  XOR2X1 U1101 ( .A(w0[8]), .B(sa20_sr[0]), .Y(N447) );
  XOR2X1 U1102 ( .A(w0[9]), .B(sa20_sr[1]), .Y(N446) );
  XOR2X1 U1103 ( .A(w0[10]), .B(sa20_sr[2]), .Y(N445) );
  XOR2X1 U1104 ( .A(w0[11]), .B(sa20_sr[3]), .Y(N444) );
  XOR2X1 U1105 ( .A(w0[12]), .B(sa20_sr[4]), .Y(N443) );
  XOR2X1 U1106 ( .A(w0[13]), .B(sa20_sr[5]), .Y(N442) );
  XOR2X1 U1107 ( .A(w0[14]), .B(sa20_sr[6]), .Y(N441) );
  XOR2X1 U1108 ( .A(w0[15]), .B(sa20_sr[7]), .Y(N440) );
  XOR2X1 U1109 ( .A(w3[16]), .B(sa13_sr[0]), .Y(N439) );
  XOR2X1 U1110 ( .A(w3[17]), .B(sa13_sr[1]), .Y(N438) );
  XOR2X1 U1111 ( .A(w3[18]), .B(sa13_sr[2]), .Y(N437) );
  XOR2X1 U1112 ( .A(w3[19]), .B(sa13_sr[3]), .Y(N436) );
  XOR2X1 U1113 ( .A(w3[20]), .B(sa13_sr[4]), .Y(N435) );
  XOR2X1 U1114 ( .A(w3[21]), .B(sa13_sr[5]), .Y(N434) );
  XOR2X1 U1115 ( .A(w3[22]), .B(sa13_sr[6]), .Y(N433) );
  XOR2X1 U1116 ( .A(w3[23]), .B(sa13_sr[7]), .Y(N432) );
  XOR2X1 U1117 ( .A(w2[16]), .B(sa12_sr[0]), .Y(N431) );
  XOR2X1 U1118 ( .A(w2[17]), .B(sa12_sr[1]), .Y(N430) );
  XOR2X1 U1119 ( .A(w2[18]), .B(sa12_sr[2]), .Y(N429) );
  XOR2X1 U1120 ( .A(w2[19]), .B(sa12_sr[3]), .Y(N428) );
  XOR2X1 U1121 ( .A(w2[20]), .B(sa12_sr[4]), .Y(N427) );
  XOR2X1 U1122 ( .A(w2[21]), .B(sa12_sr[5]), .Y(N426) );
  XOR2X1 U1123 ( .A(w2[22]), .B(sa12_sr[6]), .Y(N425) );
  XOR2X1 U1124 ( .A(w2[23]), .B(sa12_sr[7]), .Y(N424) );
  XOR2X1 U1125 ( .A(w1[16]), .B(sa11_sr[0]), .Y(N423) );
  XOR2X1 U1126 ( .A(w1[17]), .B(sa11_sr[1]), .Y(N422) );
  XOR2X1 U1127 ( .A(w1[18]), .B(sa11_sr[2]), .Y(N421) );
  XOR2X1 U1128 ( .A(w1[19]), .B(sa11_sr[3]), .Y(N420) );
  XOR2X1 U1129 ( .A(w1[20]), .B(sa11_sr[4]), .Y(N419) );
  XOR2X1 U1130 ( .A(w1[21]), .B(sa11_sr[5]), .Y(N418) );
  XOR2X1 U1131 ( .A(w1[22]), .B(sa11_sr[6]), .Y(N417) );
  XOR2X1 U1132 ( .A(w1[23]), .B(sa11_sr[7]), .Y(N416) );
  XOR2X1 U1133 ( .A(w0[16]), .B(sa10_sr[0]), .Y(N415) );
  XOR2X1 U1134 ( .A(w0[17]), .B(sa10_sr[1]), .Y(N414) );
  XOR2X1 U1135 ( .A(w0[18]), .B(sa10_sr[2]), .Y(N413) );
  XOR2X1 U1136 ( .A(w0[19]), .B(sa10_sr[3]), .Y(N412) );
  XOR2X1 U1137 ( .A(w0[20]), .B(sa10_sr[4]), .Y(N411) );
  XOR2X1 U1138 ( .A(w0[21]), .B(sa10_sr[5]), .Y(N410) );
  XOR2X1 U1139 ( .A(w0[22]), .B(sa10_sr[6]), .Y(N409) );
  XOR2X1 U1140 ( .A(w0[23]), .B(sa10_sr[7]), .Y(N408) );
  XOR2X1 U1141 ( .A(w3[24]), .B(sa03_sr[0]), .Y(N407) );
  XOR2X1 U1142 ( .A(w3[25]), .B(sa03_sr[1]), .Y(N406) );
  XOR2X1 U1143 ( .A(w3[26]), .B(sa03_sr[2]), .Y(N405) );
  XOR2X1 U1144 ( .A(w3[27]), .B(sa03_sr[3]), .Y(N404) );
  XOR2X1 U1145 ( .A(w3[28]), .B(sa03_sr[4]), .Y(N403) );
  XOR2X1 U1146 ( .A(w3[29]), .B(sa03_sr[5]), .Y(N402) );
  XOR2X1 U1147 ( .A(w3[30]), .B(sa03_sr[6]), .Y(N401) );
  XOR2X1 U1148 ( .A(w3[31]), .B(sa03_sr[7]), .Y(N400) );
  XOR2X1 U1149 ( .A(w2[24]), .B(sa02_sr[0]), .Y(N399) );
  XOR2X1 U1150 ( .A(w2[25]), .B(sa02_sr[1]), .Y(N398) );
  XOR2X1 U1151 ( .A(w2[26]), .B(sa02_sr[2]), .Y(N397) );
  XOR2X1 U1152 ( .A(w2[27]), .B(sa02_sr[3]), .Y(N396) );
  XOR2X1 U1153 ( .A(w2[28]), .B(sa02_sr[4]), .Y(N395) );
  XOR2X1 U1154 ( .A(w2[29]), .B(sa02_sr[5]), .Y(N394) );
  XOR2X1 U1155 ( .A(w2[30]), .B(sa02_sr[6]), .Y(N393) );
  XOR2X1 U1156 ( .A(w2[31]), .B(sa02_sr[7]), .Y(N392) );
  XOR2X1 U1157 ( .A(w1[24]), .B(sa01_sr[0]), .Y(N391) );
  XOR2X1 U1158 ( .A(w1[25]), .B(sa01_sr[1]), .Y(N390) );
  MX2X1 U1159 ( .A(sa33_next[7]), .B(n629), .S0(n583), .Y(N39) );
  XOR2X1 U1160 ( .A(w3[7]), .B(text_in_r[7]), .Y(n629) );
  XOR2X1 U1161 ( .A(w1[26]), .B(sa01_sr[2]), .Y(N389) );
  XOR2X1 U1162 ( .A(w1[27]), .B(sa01_sr[3]), .Y(N388) );
  XOR2X1 U1163 ( .A(w1[28]), .B(sa01_sr[4]), .Y(N387) );
  XOR2X1 U1164 ( .A(w1[29]), .B(sa01_sr[5]), .Y(N386) );
  XOR2X1 U1165 ( .A(w1[30]), .B(sa01_sr[6]), .Y(N385) );
  XOR2X1 U1166 ( .A(w1[31]), .B(sa01_sr[7]), .Y(N384) );
  XOR2X1 U1167 ( .A(w0[24]), .B(sa00_sr[0]), .Y(N383) );
  XOR2X1 U1168 ( .A(w0[25]), .B(sa00_sr[1]), .Y(N382) );
  XOR2X1 U1169 ( .A(w0[26]), .B(sa00_sr[2]), .Y(N381) );
  XOR2X1 U1170 ( .A(w0[27]), .B(sa00_sr[3]), .Y(N380) );
  MX2X1 U1171 ( .A(sa33_next[6]), .B(n630), .S0(n583), .Y(N38) );
  XOR2X1 U1172 ( .A(w3[6]), .B(text_in_r[6]), .Y(n630) );
  XOR2X1 U1173 ( .A(w0[28]), .B(sa00_sr[4]), .Y(N379) );
  XOR2X1 U1174 ( .A(w0[29]), .B(sa00_sr[5]), .Y(N378) );
  XOR2X1 U1175 ( .A(w0[30]), .B(sa00_sr[6]), .Y(N377) );
  XOR2X1 U1176 ( .A(w0[31]), .B(sa00_sr[7]), .Y(N376) );
  MX2X1 U1177 ( .A(sa33_next[5]), .B(n631), .S0(n583), .Y(N37) );
  XOR2X1 U1178 ( .A(w3[5]), .B(text_in_r[5]), .Y(n631) );
  MX2X1 U1179 ( .A(sa33_next[4]), .B(n632), .S0(n583), .Y(N36) );
  XOR2X1 U1180 ( .A(w3[4]), .B(text_in_r[4]), .Y(n632) );
  MX2X1 U1181 ( .A(sa33_next[3]), .B(n633), .S0(n583), .Y(N35) );
  XOR2X1 U1182 ( .A(w3[3]), .B(text_in_r[3]), .Y(n633) );
  MX2X1 U1183 ( .A(sa33_next[2]), .B(n634), .S0(n583), .Y(N34) );
  XOR2X1 U1184 ( .A(w3[2]), .B(text_in_r[2]), .Y(n634) );
  MX2X1 U1185 ( .A(sa33_next[1]), .B(n635), .S0(n583), .Y(N33) );
  XOR2X1 U1186 ( .A(w3[1]), .B(text_in_r[1]), .Y(n635) );
  MX2X1 U1187 ( .A(sa33_next[0]), .B(n636), .S0(n583), .Y(N32) );
  XOR2X1 U1188 ( .A(w3[0]), .B(text_in_r[0]), .Y(n636) );
  MX2X1 U1189 ( .A(sa00_next[7]), .B(n637), .S0(n583), .Y(N279) );
  XOR2X1 U1190 ( .A(w0[31]), .B(text_in_r[127]), .Y(n637) );
  MX2X1 U1191 ( .A(sa00_next[6]), .B(n638), .S0(n583), .Y(N278) );
  XOR2X1 U1192 ( .A(w0[30]), .B(text_in_r[126]), .Y(n638) );
  MX2X1 U1193 ( .A(sa00_next[5]), .B(n639), .S0(n583), .Y(N277) );
  XOR2X1 U1194 ( .A(w0[29]), .B(text_in_r[125]), .Y(n639) );
  MX2X1 U1195 ( .A(sa00_next[4]), .B(n640), .S0(n584), .Y(N276) );
  XOR2X1 U1196 ( .A(w0[28]), .B(text_in_r[124]), .Y(n640) );
  MX2X1 U1197 ( .A(sa00_next[3]), .B(n641), .S0(n584), .Y(N275) );
  XOR2X1 U1198 ( .A(w0[27]), .B(text_in_r[123]), .Y(n641) );
  MX2X1 U1199 ( .A(sa00_next[2]), .B(n642), .S0(n584), .Y(N274) );
  XOR2X1 U1200 ( .A(w0[26]), .B(text_in_r[122]), .Y(n642) );
  MX2X1 U1201 ( .A(sa00_next[1]), .B(n643), .S0(n584), .Y(N273) );
  XOR2X1 U1202 ( .A(w0[25]), .B(text_in_r[121]), .Y(n643) );
  MX2X1 U1203 ( .A(sa00_next[0]), .B(n644), .S0(n584), .Y(N272) );
  XOR2X1 U1204 ( .A(w0[24]), .B(text_in_r[120]), .Y(n644) );
  MX2X1 U1205 ( .A(sa10_next[7]), .B(n645), .S0(n584), .Y(N263) );
  XOR2X1 U1206 ( .A(w0[23]), .B(text_in_r[119]), .Y(n645) );
  MX2X1 U1207 ( .A(sa10_next[6]), .B(n646), .S0(n584), .Y(N262) );
  XOR2X1 U1208 ( .A(w0[22]), .B(text_in_r[118]), .Y(n646) );
  MX2X1 U1209 ( .A(sa10_next[5]), .B(n647), .S0(n584), .Y(N261) );
  XOR2X1 U1210 ( .A(w0[21]), .B(text_in_r[117]), .Y(n647) );
  MX2X1 U1211 ( .A(sa10_next[4]), .B(n648), .S0(n584), .Y(N260) );
  XOR2X1 U1212 ( .A(w0[20]), .B(text_in_r[116]), .Y(n648) );
  MX2X1 U1213 ( .A(sa10_next[3]), .B(n649), .S0(n584), .Y(N259) );
  XOR2X1 U1214 ( .A(w0[19]), .B(text_in_r[115]), .Y(n649) );
  MX2X1 U1215 ( .A(sa10_next[2]), .B(n650), .S0(n584), .Y(N258) );
  XOR2X1 U1216 ( .A(w0[18]), .B(text_in_r[114]), .Y(n650) );
  MX2X1 U1217 ( .A(sa10_next[1]), .B(n651), .S0(n584), .Y(N257) );
  XOR2X1 U1218 ( .A(w0[17]), .B(text_in_r[113]), .Y(n651) );
  MX2X1 U1219 ( .A(sa10_next[0]), .B(n652), .S0(n584), .Y(N256) );
  XOR2X1 U1220 ( .A(w0[16]), .B(text_in_r[112]), .Y(n652) );
  MX2X1 U1221 ( .A(sa20_next[7]), .B(n653), .S0(n585), .Y(N247) );
  XOR2X1 U1222 ( .A(w0[15]), .B(text_in_r[111]), .Y(n653) );
  MX2X1 U1223 ( .A(sa20_next[6]), .B(n654), .S0(n585), .Y(N246) );
  XOR2X1 U1224 ( .A(w0[14]), .B(text_in_r[110]), .Y(n654) );
  MX2X1 U1225 ( .A(sa20_next[5]), .B(n655), .S0(n585), .Y(N245) );
  XOR2X1 U1226 ( .A(w0[13]), .B(text_in_r[109]), .Y(n655) );
  MX2X1 U1227 ( .A(sa20_next[4]), .B(n656), .S0(n585), .Y(N244) );
  XOR2X1 U1228 ( .A(w0[12]), .B(text_in_r[108]), .Y(n656) );
  MX2X1 U1229 ( .A(sa20_next[3]), .B(n657), .S0(n585), .Y(N243) );
  XOR2X1 U1230 ( .A(w0[11]), .B(text_in_r[107]), .Y(n657) );
  MX2X1 U1231 ( .A(sa20_next[2]), .B(n658), .S0(n585), .Y(N242) );
  XOR2X1 U1232 ( .A(w0[10]), .B(text_in_r[106]), .Y(n658) );
  MX2X1 U1233 ( .A(sa20_next[1]), .B(n659), .S0(n585), .Y(N241) );
  XOR2X1 U1234 ( .A(w0[9]), .B(text_in_r[105]), .Y(n659) );
  MX2X1 U1235 ( .A(sa20_next[0]), .B(n660), .S0(n585), .Y(N240) );
  XOR2X1 U1236 ( .A(w0[8]), .B(text_in_r[104]), .Y(n660) );
  MX2X1 U1237 ( .A(sa30_next[7]), .B(n661), .S0(n585), .Y(N231) );
  XOR2X1 U1238 ( .A(w0[7]), .B(text_in_r[103]), .Y(n661) );
  MX2X1 U1239 ( .A(sa30_next[6]), .B(n662), .S0(n585), .Y(N230) );
  XOR2X1 U1240 ( .A(w0[6]), .B(text_in_r[102]), .Y(n662) );
  MX2X1 U1241 ( .A(sa30_next[5]), .B(n663), .S0(n585), .Y(N229) );
  XOR2X1 U1242 ( .A(w0[5]), .B(text_in_r[101]), .Y(n663) );
  MX2X1 U1243 ( .A(sa30_next[4]), .B(n664), .S0(n585), .Y(N228) );
  XOR2X1 U1244 ( .A(w0[4]), .B(text_in_r[100]), .Y(n664) );
  MX2X1 U1245 ( .A(sa30_next[3]), .B(n665), .S0(n585), .Y(N227) );
  XOR2X1 U1246 ( .A(w0[3]), .B(text_in_r[99]), .Y(n665) );
  MX2X1 U1247 ( .A(sa30_next[2]), .B(n666), .S0(n586), .Y(N226) );
  XOR2X1 U1248 ( .A(w0[2]), .B(text_in_r[98]), .Y(n666) );
  MX2X1 U1249 ( .A(sa30_next[1]), .B(n667), .S0(n586), .Y(N225) );
  XOR2X1 U1250 ( .A(w0[1]), .B(text_in_r[97]), .Y(n667) );
  MX2X1 U1251 ( .A(sa30_next[0]), .B(n668), .S0(n586), .Y(N224) );
  XOR2X1 U1252 ( .A(w0[0]), .B(text_in_r[96]), .Y(n668) );
  MX2X1 U1253 ( .A(sa01_next[7]), .B(n669), .S0(n586), .Y(N215) );
  XOR2X1 U1254 ( .A(w1[31]), .B(text_in_r[95]), .Y(n669) );
  MX2X1 U1255 ( .A(sa01_next[6]), .B(n670), .S0(n586), .Y(N214) );
  XOR2X1 U1256 ( .A(w1[30]), .B(text_in_r[94]), .Y(n670) );
  MX2X1 U1257 ( .A(sa01_next[5]), .B(n671), .S0(n586), .Y(N213) );
  XOR2X1 U1258 ( .A(w1[29]), .B(text_in_r[93]), .Y(n671) );
  MX2X1 U1259 ( .A(sa01_next[4]), .B(n672), .S0(n586), .Y(N212) );
  XOR2X1 U1260 ( .A(w1[28]), .B(text_in_r[92]), .Y(n672) );
  MX2X1 U1261 ( .A(sa01_next[3]), .B(n673), .S0(n586), .Y(N211) );
  XOR2X1 U1262 ( .A(w1[27]), .B(text_in_r[91]), .Y(n673) );
  MX2X1 U1263 ( .A(sa01_next[2]), .B(n674), .S0(n586), .Y(N210) );
  XOR2X1 U1264 ( .A(w1[26]), .B(text_in_r[90]), .Y(n674) );
  NOR3BX1 U1265 ( .AN(dcnt[0]), .B(n675), .C(dcnt[1]), .Y(N21) );
  OR3XL U1266 ( .A(n730), .B(ld), .C(dcnt[3]), .Y(n675) );
  MX2X1 U1267 ( .A(sa01_next[1]), .B(n676), .S0(n586), .Y(N209) );
  XOR2X1 U1268 ( .A(w1[25]), .B(text_in_r[89]), .Y(n676) );
  MX2X1 U1269 ( .A(sa01_next[0]), .B(n677), .S0(n586), .Y(N208) );
  XOR2X1 U1270 ( .A(w1[24]), .B(text_in_r[88]), .Y(n677) );
  MX2X1 U1271 ( .A(sa11_next[7]), .B(n678), .S0(n586), .Y(N199) );
  XOR2X1 U1272 ( .A(w1[23]), .B(text_in_r[87]), .Y(n678) );
  MX2X1 U1273 ( .A(sa11_next[6]), .B(n679), .S0(n586), .Y(N198) );
  XOR2X1 U1274 ( .A(w1[22]), .B(text_in_r[86]), .Y(n679) );
  MX2X1 U1275 ( .A(sa11_next[5]), .B(n680), .S0(n587), .Y(N197) );
  XOR2X1 U1276 ( .A(w1[21]), .B(text_in_r[85]), .Y(n680) );
  MX2X1 U1277 ( .A(sa11_next[4]), .B(n681), .S0(n587), .Y(N196) );
  XOR2X1 U1278 ( .A(w1[20]), .B(text_in_r[84]), .Y(n681) );
  MX2X1 U1279 ( .A(sa11_next[3]), .B(n682), .S0(n587), .Y(N195) );
  XOR2X1 U1280 ( .A(w1[19]), .B(text_in_r[83]), .Y(n682) );
  MX2X1 U1281 ( .A(sa11_next[2]), .B(n683), .S0(n587), .Y(N194) );
  XOR2X1 U1282 ( .A(w1[18]), .B(text_in_r[82]), .Y(n683) );
  MX2X1 U1283 ( .A(sa11_next[1]), .B(n684), .S0(n587), .Y(N193) );
  XOR2X1 U1284 ( .A(w1[17]), .B(text_in_r[81]), .Y(n684) );
  MX2X1 U1285 ( .A(sa11_next[0]), .B(n685), .S0(n587), .Y(N192) );
  XOR2X1 U1286 ( .A(w1[16]), .B(text_in_r[80]), .Y(n685) );
  MX2X1 U1287 ( .A(sa21_next[7]), .B(n686), .S0(n587), .Y(N183) );
  XOR2X1 U1288 ( .A(w1[15]), .B(text_in_r[79]), .Y(n686) );
  MX2X1 U1289 ( .A(sa21_next[6]), .B(n687), .S0(n587), .Y(N182) );
  XOR2X1 U1290 ( .A(w1[14]), .B(text_in_r[78]), .Y(n687) );
  MX2X1 U1291 ( .A(sa21_next[5]), .B(n688), .S0(n587), .Y(N181) );
  XOR2X1 U1292 ( .A(w1[13]), .B(text_in_r[77]), .Y(n688) );
  MX2X1 U1293 ( .A(sa21_next[4]), .B(n689), .S0(n587), .Y(N180) );
  XOR2X1 U1294 ( .A(w1[12]), .B(text_in_r[76]), .Y(n689) );
  MX2X1 U1295 ( .A(sa21_next[3]), .B(n690), .S0(n587), .Y(N179) );
  XOR2X1 U1296 ( .A(w1[11]), .B(text_in_r[75]), .Y(n690) );
  MX2X1 U1297 ( .A(sa21_next[2]), .B(n691), .S0(n587), .Y(N178) );
  XOR2X1 U1298 ( .A(w1[10]), .B(text_in_r[74]), .Y(n691) );
  MX2X1 U1299 ( .A(sa21_next[1]), .B(n692), .S0(n587), .Y(N177) );
  XOR2X1 U1300 ( .A(w1[9]), .B(text_in_r[73]), .Y(n692) );
  MX2X1 U1301 ( .A(sa21_next[0]), .B(n693), .S0(n588), .Y(N176) );
  XOR2X1 U1302 ( .A(w1[8]), .B(text_in_r[72]), .Y(n693) );
  MX2X1 U1303 ( .A(sa31_next[7]), .B(n694), .S0(n588), .Y(N167) );
  XOR2X1 U1304 ( .A(w1[7]), .B(text_in_r[71]), .Y(n694) );
  MX2X1 U1305 ( .A(sa31_next[6]), .B(n695), .S0(n588), .Y(N166) );
  XOR2X1 U1306 ( .A(w1[6]), .B(text_in_r[70]), .Y(n695) );
  MX2X1 U1307 ( .A(sa31_next[5]), .B(n696), .S0(n588), .Y(N165) );
  XOR2X1 U1308 ( .A(w1[5]), .B(text_in_r[69]), .Y(n696) );
  MX2X1 U1309 ( .A(sa31_next[4]), .B(n697), .S0(n588), .Y(N164) );
  XOR2X1 U1310 ( .A(w1[4]), .B(text_in_r[68]), .Y(n697) );
  MX2X1 U1311 ( .A(sa31_next[3]), .B(n698), .S0(n588), .Y(N163) );
  XOR2X1 U1312 ( .A(w1[3]), .B(text_in_r[67]), .Y(n698) );
  MX2X1 U1313 ( .A(sa31_next[2]), .B(n699), .S0(n588), .Y(N162) );
  XOR2X1 U1314 ( .A(w1[2]), .B(text_in_r[66]), .Y(n699) );
  MX2X1 U1315 ( .A(sa31_next[1]), .B(n700), .S0(n588), .Y(N161) );
  XOR2X1 U1316 ( .A(w1[1]), .B(text_in_r[65]), .Y(n700) );
  MX2X1 U1317 ( .A(sa31_next[0]), .B(n701), .S0(n588), .Y(N160) );
  XOR2X1 U1318 ( .A(w1[0]), .B(text_in_r[64]), .Y(n701) );
  MX2X1 U1319 ( .A(sa02_next[7]), .B(n702), .S0(n588), .Y(N151) );
  XOR2X1 U1320 ( .A(w2[31]), .B(text_in_r[63]), .Y(n702) );
  MX2X1 U1321 ( .A(sa02_next[6]), .B(n703), .S0(n588), .Y(N150) );
  XOR2X1 U1322 ( .A(w2[30]), .B(text_in_r[62]), .Y(n703) );
  MX2X1 U1323 ( .A(sa02_next[5]), .B(n704), .S0(n588), .Y(N149) );
  XOR2X1 U1324 ( .A(w2[29]), .B(text_in_r[61]), .Y(n704) );
  MX2X1 U1325 ( .A(sa02_next[4]), .B(n705), .S0(n588), .Y(N148) );
  XOR2X1 U1326 ( .A(w2[28]), .B(text_in_r[60]), .Y(n705) );
  MX2X1 U1327 ( .A(sa02_next[3]), .B(n706), .S0(n581), .Y(N147) );
  XOR2X1 U1328 ( .A(w2[27]), .B(text_in_r[59]), .Y(n706) );
  MX2X1 U1329 ( .A(sa02_next[2]), .B(n707), .S0(n582), .Y(N146) );
  XOR2X1 U1330 ( .A(w2[26]), .B(text_in_r[58]), .Y(n707) );
  MX2X1 U1331 ( .A(sa02_next[1]), .B(n708), .S0(n588), .Y(N145) );
  XOR2X1 U1332 ( .A(w2[25]), .B(text_in_r[57]), .Y(n708) );
  MX2X1 U1333 ( .A(sa02_next[0]), .B(n709), .S0(n731), .Y(N144) );
  XOR2X1 U1334 ( .A(w2[24]), .B(text_in_r[56]), .Y(n709) );
  MX2X1 U1335 ( .A(sa12_next[7]), .B(n710), .S0(n587), .Y(N135) );
  XOR2X1 U1336 ( .A(w2[23]), .B(text_in_r[55]), .Y(n710) );
  MX2X1 U1337 ( .A(sa12_next[6]), .B(n711), .S0(n586), .Y(N134) );
  XOR2X1 U1338 ( .A(w2[22]), .B(text_in_r[54]), .Y(n711) );
  MX2X1 U1339 ( .A(sa12_next[5]), .B(n712), .S0(n584), .Y(N133) );
  XOR2X1 U1340 ( .A(w2[21]), .B(text_in_r[53]), .Y(n712) );
  MX2X1 U1341 ( .A(sa12_next[4]), .B(n713), .S0(n583), .Y(N132) );
  XOR2X1 U1342 ( .A(w2[20]), .B(text_in_r[52]), .Y(n713) );
  MX2X1 U1343 ( .A(sa12_next[3]), .B(n714), .S0(n585), .Y(N131) );
  XOR2X1 U1344 ( .A(w2[19]), .B(text_in_r[51]), .Y(n714) );
  MX2X1 U1345 ( .A(sa12_next[2]), .B(n715), .S0(n581), .Y(N130) );
  XOR2X1 U1346 ( .A(w2[18]), .B(text_in_r[50]), .Y(n715) );
  MX2X1 U1347 ( .A(sa12_next[1]), .B(n716), .S0(n582), .Y(N129) );
  XOR2X1 U1348 ( .A(w2[17]), .B(text_in_r[49]), .Y(n716) );
  MX2X1 U1349 ( .A(sa12_next[0]), .B(n717), .S0(n588), .Y(N128) );
  XOR2X1 U1350 ( .A(w2[16]), .B(text_in_r[48]), .Y(n717) );
  MX2X1 U1351 ( .A(sa22_next[7]), .B(n718), .S0(n731), .Y(N119) );
  XOR2X1 U1352 ( .A(w2[15]), .B(text_in_r[47]), .Y(n718) );
  MX2X1 U1353 ( .A(sa22_next[6]), .B(n719), .S0(n731), .Y(N118) );
  XOR2X1 U1354 ( .A(w2[14]), .B(text_in_r[46]), .Y(n719) );
  MX2X1 U1355 ( .A(sa22_next[5]), .B(n720), .S0(n731), .Y(N117) );
  XOR2X1 U1356 ( .A(w2[13]), .B(text_in_r[45]), .Y(n720) );
  MX2X1 U1357 ( .A(sa22_next[4]), .B(n721), .S0(n731), .Y(N116) );
  XOR2X1 U1358 ( .A(w2[12]), .B(text_in_r[44]), .Y(n721) );
  MX2X1 U1359 ( .A(sa22_next[3]), .B(n722), .S0(n731), .Y(N115) );
  XOR2X1 U1360 ( .A(w2[11]), .B(text_in_r[43]), .Y(n722) );
  MX2X1 U1361 ( .A(sa22_next[2]), .B(n723), .S0(n731), .Y(N114) );
  XOR2X1 U1362 ( .A(w2[10]), .B(text_in_r[42]), .Y(n723) );
  MX2X1 U1363 ( .A(sa22_next[1]), .B(n724), .S0(n731), .Y(N113) );
  XOR2X1 U1364 ( .A(w2[9]), .B(text_in_r[41]), .Y(n724) );
  MX2X1 U1365 ( .A(sa22_next[0]), .B(n725), .S0(n731), .Y(N112) );
  XOR2X1 U1366 ( .A(w2[8]), .B(text_in_r[40]), .Y(n725) );
  MX2X1 U1367 ( .A(sa32_next[7]), .B(n726), .S0(n731), .Y(N103) );
  XOR2X1 U1368 ( .A(w2[7]), .B(text_in_r[39]), .Y(n726) );
  MX2X1 U1369 ( .A(sa32_next[6]), .B(n727), .S0(n731), .Y(N102) );
  XOR2X1 U1370 ( .A(w2[6]), .B(text_in_r[38]), .Y(n727) );
  MX2X1 U1371 ( .A(sa32_next[5]), .B(n728), .S0(n731), .Y(N101) );
  XOR2X1 U1372 ( .A(w2[5]), .B(text_in_r[37]), .Y(n728) );
  MX2X1 U1373 ( .A(sa32_next[4]), .B(n729), .S0(n731), .Y(N100) );
  XOR2X1 U1374 ( .A(w2[4]), .B(text_in_r[36]), .Y(n729) );
  MX2X1 \u0/U130  ( .A(\u0/N10 ), .B(key[127]), .S0(ld), .Y(\u0/n1 ) );
  MX2X1 \u0/U129  ( .A(\u0/N78 ), .B(key[93]), .S0(ld), .Y(\u0/n10 ) );
  MX2X1 \u0/U128  ( .A(\u0/N232 ), .B(key[7]), .S0(ld), .Y(\u0/n100 ) );
  MX2X1 \u0/U127  ( .A(\u0/N35 ), .B(key[102]), .S0(ld), .Y(\u0/n101 ) );
  MX2X1 \u0/U126  ( .A(\u0/N101 ), .B(key[70]), .S0(ld), .Y(\u0/n102 ) );
  MX2X1 \u0/U125  ( .A(\u0/N167 ), .B(key[38]), .S0(ld), .Y(\u0/n103 ) );
  MX2X1 \u0/U124  ( .A(\u0/N233 ), .B(key[6]), .S0(ld), .Y(\u0/n104 ) );
  MX2X1 \u0/U123  ( .A(\u0/N36 ), .B(key[101]), .S0(ld), .Y(\u0/n105 ) );
  MX2X1 \u0/U122  ( .A(\u0/N102 ), .B(key[69]), .S0(ld), .Y(\u0/n106 ) );
  MX2X1 \u0/U121  ( .A(\u0/N168 ), .B(key[37]), .S0(ld), .Y(\u0/n107 ) );
  MX2X1 \u0/U120  ( .A(\u0/N234 ), .B(key[5]), .S0(ld), .Y(\u0/n108 ) );
  MX2X1 \u0/U119  ( .A(\u0/N37 ), .B(key[100]), .S0(ld), .Y(\u0/n109 ) );
  MX2X1 \u0/U118  ( .A(\u0/N144 ), .B(key[61]), .S0(ld), .Y(\u0/n11 ) );
  MX2X1 \u0/U117  ( .A(\u0/N103 ), .B(key[68]), .S0(ld), .Y(\u0/n110 ) );
  MX2X1 \u0/U116  ( .A(\u0/N169 ), .B(key[36]), .S0(ld), .Y(\u0/n111 ) );
  MX2X1 \u0/U115  ( .A(\u0/N235 ), .B(key[4]), .S0(ld), .Y(\u0/n112 ) );
  MX2X1 \u0/U114  ( .A(\u0/N38 ), .B(key[99]), .S0(ld), .Y(\u0/n113 ) );
  MX2X1 \u0/U113  ( .A(\u0/N104 ), .B(key[67]), .S0(ld), .Y(\u0/n114 ) );
  MX2X1 \u0/U112  ( .A(\u0/N170 ), .B(key[35]), .S0(ld), .Y(\u0/n115 ) );
  MX2X1 \u0/U111  ( .A(\u0/N236 ), .B(key[3]), .S0(ld), .Y(\u0/n116 ) );
  MX2X1 \u0/U110  ( .A(\u0/N39 ), .B(key[98]), .S0(ld), .Y(\u0/n117 ) );
  MX2X1 \u0/U109  ( .A(\u0/N105 ), .B(key[66]), .S0(ld), .Y(\u0/n118 ) );
  MX2X1 \u0/U108  ( .A(\u0/N171 ), .B(key[34]), .S0(ld), .Y(\u0/n119 ) );
  MX2X1 \u0/U107  ( .A(\u0/N210 ), .B(key[29]), .S0(ld), .Y(\u0/n12 ) );
  MX2X1 \u0/U106  ( .A(\u0/N237 ), .B(key[2]), .S0(ld), .Y(\u0/n120 ) );
  MX2X1 \u0/U105  ( .A(\u0/N40 ), .B(key[97]), .S0(ld), .Y(\u0/n121 ) );
  MX2X1 \u0/U104  ( .A(\u0/N106 ), .B(key[65]), .S0(ld), .Y(\u0/n122 ) );
  MX2X1 \u0/U103  ( .A(\u0/N172 ), .B(key[33]), .S0(ld), .Y(\u0/n123 ) );
  MX2X1 \u0/U102  ( .A(\u0/N238 ), .B(key[1]), .S0(ld), .Y(\u0/n124 ) );
  MX2X1 \u0/U101  ( .A(\u0/N41 ), .B(key[96]), .S0(ld), .Y(\u0/n125 ) );
  MX2X1 \u0/U100  ( .A(\u0/N107 ), .B(key[64]), .S0(ld), .Y(\u0/n126 ) );
  MX2X1 \u0/U99  ( .A(\u0/N173 ), .B(key[32]), .S0(ld), .Y(\u0/n127 ) );
  MX2X1 \u0/U98  ( .A(\u0/N239 ), .B(key[0]), .S0(ld), .Y(\u0/n128 ) );
  MX2X1 \u0/U97  ( .A(\u0/N13 ), .B(key[124]), .S0(ld), .Y(\u0/n13 ) );
  MX2X1 \u0/U96  ( .A(\u0/N79 ), .B(key[92]), .S0(ld), .Y(\u0/n14 ) );
  MX2X1 \u0/U95  ( .A(\u0/N145 ), .B(key[60]), .S0(ld), .Y(\u0/n15 ) );
  MX2X1 \u0/U94  ( .A(\u0/N211 ), .B(key[28]), .S0(ld), .Y(\u0/n16 ) );
  MX2X1 \u0/U93  ( .A(\u0/N14 ), .B(key[123]), .S0(ld), .Y(\u0/n17 ) );
  MX2X1 \u0/U92  ( .A(\u0/N80 ), .B(key[91]), .S0(ld), .Y(\u0/n18 ) );
  MX2X1 \u0/U91  ( .A(\u0/N146 ), .B(key[59]), .S0(ld), .Y(\u0/n19 ) );
  MX2X1 \u0/U90  ( .A(\u0/N76 ), .B(key[95]), .S0(ld), .Y(\u0/n2 ) );
  MX2X1 \u0/U89  ( .A(\u0/N212 ), .B(key[27]), .S0(ld), .Y(\u0/n20 ) );
  MX2X1 \u0/U88  ( .A(\u0/N15 ), .B(key[122]), .S0(ld), .Y(\u0/n21 ) );
  MX2X1 \u0/U87  ( .A(\u0/N81 ), .B(key[90]), .S0(ld), .Y(\u0/n22 ) );
  MX2X1 \u0/U86  ( .A(\u0/N147 ), .B(key[58]), .S0(ld), .Y(\u0/n23 ) );
  MX2X1 \u0/U85  ( .A(\u0/N213 ), .B(key[26]), .S0(ld), .Y(\u0/n24 ) );
  MX2X1 \u0/U84  ( .A(\u0/N16 ), .B(key[121]), .S0(ld), .Y(\u0/n25 ) );
  MX2X1 \u0/U83  ( .A(\u0/N82 ), .B(key[89]), .S0(ld), .Y(\u0/n26 ) );
  MX2X1 \u0/U82  ( .A(\u0/N148 ), .B(key[57]), .S0(ld), .Y(\u0/n27 ) );
  MX2X1 \u0/U81  ( .A(\u0/N214 ), .B(key[25]), .S0(ld), .Y(\u0/n28 ) );
  MX2X1 \u0/U80  ( .A(\u0/N17 ), .B(key[120]), .S0(ld), .Y(\u0/n29 ) );
  MX2X1 \u0/U79  ( .A(\u0/N142 ), .B(key[63]), .S0(ld), .Y(\u0/n3 ) );
  MX2X1 \u0/U78  ( .A(\u0/N83 ), .B(key[88]), .S0(ld), .Y(\u0/n30 ) );
  MX2X1 \u0/U77  ( .A(\u0/N149 ), .B(key[56]), .S0(ld), .Y(\u0/n31 ) );
  MX2X1 \u0/U76  ( .A(\u0/N215 ), .B(key[24]), .S0(ld), .Y(\u0/n32 ) );
  MX2X1 \u0/U75  ( .A(\u0/N18 ), .B(key[119]), .S0(ld), .Y(\u0/n33 ) );
  MX2X1 \u0/U74  ( .A(\u0/N84 ), .B(key[87]), .S0(ld), .Y(\u0/n34 ) );
  MX2X1 \u0/U73  ( .A(\u0/N150 ), .B(key[55]), .S0(ld), .Y(\u0/n35 ) );
  MX2X1 \u0/U72  ( .A(\u0/N216 ), .B(key[23]), .S0(ld), .Y(\u0/n36 ) );
  MX2X1 \u0/U71  ( .A(\u0/N19 ), .B(key[118]), .S0(ld), .Y(\u0/n37 ) );
  MX2X1 \u0/U70  ( .A(\u0/N85 ), .B(key[86]), .S0(ld), .Y(\u0/n38 ) );
  MX2X1 \u0/U69  ( .A(\u0/N151 ), .B(key[54]), .S0(ld), .Y(\u0/n39 ) );
  MX2X1 \u0/U68  ( .A(\u0/N208 ), .B(key[31]), .S0(ld), .Y(\u0/n4 ) );
  MX2X1 \u0/U67  ( .A(\u0/N217 ), .B(key[22]), .S0(ld), .Y(\u0/n40 ) );
  MX2X1 \u0/U66  ( .A(\u0/N20 ), .B(key[117]), .S0(ld), .Y(\u0/n41 ) );
  MX2X1 \u0/U65  ( .A(\u0/N86 ), .B(key[85]), .S0(ld), .Y(\u0/n42 ) );
  MX2X1 \u0/U64  ( .A(\u0/N152 ), .B(key[53]), .S0(ld), .Y(\u0/n43 ) );
  MX2X1 \u0/U63  ( .A(\u0/N218 ), .B(key[21]), .S0(ld), .Y(\u0/n44 ) );
  MX2X1 \u0/U62  ( .A(\u0/N21 ), .B(key[116]), .S0(ld), .Y(\u0/n45 ) );
  MX2X1 \u0/U61  ( .A(\u0/N87 ), .B(key[84]), .S0(ld), .Y(\u0/n46 ) );
  MX2X1 \u0/U60  ( .A(\u0/N153 ), .B(key[52]), .S0(ld), .Y(\u0/n47 ) );
  MX2X1 \u0/U59  ( .A(\u0/N219 ), .B(key[20]), .S0(ld), .Y(\u0/n48 ) );
  MX2X1 \u0/U58  ( .A(\u0/N22 ), .B(key[115]), .S0(ld), .Y(\u0/n49 ) );
  MX2X1 \u0/U57  ( .A(\u0/N11 ), .B(key[126]), .S0(ld), .Y(\u0/n5 ) );
  MX2X1 \u0/U56  ( .A(\u0/N88 ), .B(key[83]), .S0(ld), .Y(\u0/n50 ) );
  MX2X1 \u0/U55  ( .A(\u0/N154 ), .B(key[51]), .S0(ld), .Y(\u0/n51 ) );
  MX2X1 \u0/U54  ( .A(\u0/N220 ), .B(key[19]), .S0(ld), .Y(\u0/n52 ) );
  MX2X1 \u0/U53  ( .A(\u0/N23 ), .B(key[114]), .S0(ld), .Y(\u0/n53 ) );
  MX2X1 \u0/U52  ( .A(\u0/N89 ), .B(key[82]), .S0(ld), .Y(\u0/n54 ) );
  MX2X1 \u0/U51  ( .A(\u0/N155 ), .B(key[50]), .S0(ld), .Y(\u0/n55 ) );
  MX2X1 \u0/U50  ( .A(\u0/N221 ), .B(key[18]), .S0(ld), .Y(\u0/n56 ) );
  MX2X1 \u0/U49  ( .A(\u0/N24 ), .B(key[113]), .S0(ld), .Y(\u0/n57 ) );
  MX2X1 \u0/U48  ( .A(\u0/N90 ), .B(key[81]), .S0(ld), .Y(\u0/n58 ) );
  MX2X1 \u0/U47  ( .A(\u0/N156 ), .B(key[49]), .S0(ld), .Y(\u0/n59 ) );
  MX2X1 \u0/U46  ( .A(\u0/N77 ), .B(key[94]), .S0(ld), .Y(\u0/n6 ) );
  MX2X1 \u0/U45  ( .A(\u0/N222 ), .B(key[17]), .S0(ld), .Y(\u0/n60 ) );
  MX2X1 \u0/U44  ( .A(\u0/N25 ), .B(key[112]), .S0(ld), .Y(\u0/n61 ) );
  MX2X1 \u0/U43  ( .A(\u0/N91 ), .B(key[80]), .S0(ld), .Y(\u0/n62 ) );
  MX2X1 \u0/U42  ( .A(\u0/N157 ), .B(key[48]), .S0(ld), .Y(\u0/n63 ) );
  MX2X1 \u0/U41  ( .A(\u0/N223 ), .B(key[16]), .S0(ld), .Y(\u0/n64 ) );
  MX2X1 \u0/U40  ( .A(\u0/N26 ), .B(key[111]), .S0(ld), .Y(\u0/n65 ) );
  MX2X1 \u0/U39  ( .A(\u0/N92 ), .B(key[79]), .S0(ld), .Y(\u0/n66 ) );
  MX2X1 \u0/U38  ( .A(\u0/N158 ), .B(key[47]), .S0(ld), .Y(\u0/n67 ) );
  MX2X1 \u0/U37  ( .A(\u0/N224 ), .B(key[15]), .S0(ld), .Y(\u0/n68 ) );
  MX2X1 \u0/U36  ( .A(\u0/N27 ), .B(key[110]), .S0(ld), .Y(\u0/n69 ) );
  MX2X1 \u0/U35  ( .A(\u0/N143 ), .B(key[62]), .S0(ld), .Y(\u0/n7 ) );
  MX2X1 \u0/U34  ( .A(\u0/N93 ), .B(key[78]), .S0(ld), .Y(\u0/n70 ) );
  MX2X1 \u0/U33  ( .A(\u0/N159 ), .B(key[46]), .S0(ld), .Y(\u0/n71 ) );
  MX2X1 \u0/U32  ( .A(\u0/N225 ), .B(key[14]), .S0(ld), .Y(\u0/n72 ) );
  MX2X1 \u0/U31  ( .A(\u0/N28 ), .B(key[109]), .S0(ld), .Y(\u0/n73 ) );
  MX2X1 \u0/U30  ( .A(\u0/N94 ), .B(key[77]), .S0(ld), .Y(\u0/n74 ) );
  MX2X1 \u0/U29  ( .A(\u0/N160 ), .B(key[45]), .S0(ld), .Y(\u0/n75 ) );
  MX2X1 \u0/U28  ( .A(\u0/N226 ), .B(key[13]), .S0(ld), .Y(\u0/n76 ) );
  MX2X1 \u0/U27  ( .A(\u0/N29 ), .B(key[108]), .S0(ld), .Y(\u0/n77 ) );
  MX2X1 \u0/U26  ( .A(\u0/N95 ), .B(key[76]), .S0(ld), .Y(\u0/n78 ) );
  MX2X1 \u0/U25  ( .A(\u0/N161 ), .B(key[44]), .S0(ld), .Y(\u0/n79 ) );
  MX2X1 \u0/U24  ( .A(\u0/N209 ), .B(key[30]), .S0(ld), .Y(\u0/n8 ) );
  MX2X1 \u0/U23  ( .A(\u0/N227 ), .B(key[12]), .S0(ld), .Y(\u0/n80 ) );
  MX2X1 \u0/U22  ( .A(\u0/N30 ), .B(key[107]), .S0(ld), .Y(\u0/n81 ) );
  MX2X1 \u0/U21  ( .A(\u0/N96 ), .B(key[75]), .S0(ld), .Y(\u0/n82 ) );
  MX2X1 \u0/U20  ( .A(\u0/N162 ), .B(key[43]), .S0(ld), .Y(\u0/n83 ) );
  MX2X1 \u0/U19  ( .A(\u0/N228 ), .B(key[11]), .S0(ld), .Y(\u0/n84 ) );
  MX2X1 \u0/U18  ( .A(\u0/N31 ), .B(key[106]), .S0(ld), .Y(\u0/n85 ) );
  MX2X1 \u0/U17  ( .A(\u0/N97 ), .B(key[74]), .S0(ld), .Y(\u0/n86 ) );
  MX2X1 \u0/U16  ( .A(\u0/N163 ), .B(key[42]), .S0(ld), .Y(\u0/n87 ) );
  MX2X1 \u0/U15  ( .A(\u0/N229 ), .B(key[10]), .S0(ld), .Y(\u0/n88 ) );
  MX2X1 \u0/U14  ( .A(\u0/N32 ), .B(key[105]), .S0(ld), .Y(\u0/n89 ) );
  MX2X1 \u0/U13  ( .A(\u0/N12 ), .B(key[125]), .S0(ld), .Y(\u0/n9 ) );
  MX2X1 \u0/U12  ( .A(\u0/N98 ), .B(key[73]), .S0(ld), .Y(\u0/n90 ) );
  MX2X1 \u0/U11  ( .A(\u0/N164 ), .B(key[41]), .S0(ld), .Y(\u0/n91 ) );
  MX2X1 \u0/U10  ( .A(\u0/N230 ), .B(key[9]), .S0(ld), .Y(\u0/n92 ) );
  MX2X1 \u0/U9  ( .A(\u0/N33 ), .B(key[104]), .S0(ld), .Y(\u0/n93 ) );
  MX2X1 \u0/U8  ( .A(\u0/N99 ), .B(key[72]), .S0(ld), .Y(\u0/n94 ) );
  MX2X1 \u0/U7  ( .A(\u0/N165 ), .B(key[40]), .S0(ld), .Y(\u0/n95 ) );
  MX2X1 \u0/U6  ( .A(\u0/N231 ), .B(key[8]), .S0(ld), .Y(\u0/n96 ) );
  MX2X1 \u0/U5  ( .A(\u0/N34 ), .B(key[103]), .S0(ld), .Y(\u0/n97 ) );
  MX2X1 \u0/U4  ( .A(\u0/N100 ), .B(key[71]), .S0(ld), .Y(\u0/n98 ) );
  MX2X1 \u0/U3  ( .A(\u0/N166 ), .B(key[39]), .S0(ld), .Y(\u0/n99 ) );
  DFFHQX1 \u0/w_reg[3][6]  ( .D(\u0/n104 ), .CK(clk), .Q(w3[6]) );
  DFFHQX1 \u0/w_reg[3][30]  ( .D(\u0/n8 ), .CK(clk), .Q(w3[30]) );
  DFFHQX1 \u0/w_reg[3][22]  ( .D(\u0/n40 ), .CK(clk), .Q(w3[22]) );
  DFFHQX1 \u0/w_reg[3][14]  ( .D(\u0/n72 ), .CK(clk), .Q(w3[14]) );
  XOR2X1 \u0/U283  ( .A(w0[4]), .B(\u0/subword [4]), .Y(\u0/N37 ) );
  XOR2X1 \u0/U273  ( .A(w0[2]), .B(\u0/subword [2]), .Y(\u0/N39 ) );
  XOR2X1 \u0/U363  ( .A(w0[20]), .B(\u0/subword [20]), .Y(\u0/N21 ) );
  XOR2X1 \u0/U353  ( .A(w0[18]), .B(\u0/subword [18]), .Y(\u0/N23 ) );
  XOR2X1 \u0/U323  ( .A(w0[12]), .B(\u0/subword [12]), .Y(\u0/N29 ) );
  XOR2X1 \u0/U313  ( .A(w0[10]), .B(\u0/subword [10]), .Y(\u0/N31 ) );
  XOR2X1 \u0/U338  ( .A(w0[15]), .B(\u0/subword [15]), .Y(\u0/N26 ) );
  XOR2X1 \u0/U378  ( .A(w0[23]), .B(\u0/subword [23]), .Y(\u0/N18 ) );
  XOR2X1 \u0/U298  ( .A(w0[7]), .B(\u0/subword [7]), .Y(\u0/N34 ) );
  XOR2X1 \u0/U293  ( .A(w0[6]), .B(\u0/subword [6]), .Y(\u0/N35 ) );
  XOR2X1 \u0/U288  ( .A(w0[5]), .B(\u0/subword [5]), .Y(\u0/N36 ) );
  XOR2X1 \u0/U278  ( .A(w0[3]), .B(\u0/subword [3]), .Y(\u0/N38 ) );
  XOR2X1 \u0/U268  ( .A(w0[1]), .B(\u0/subword [1]), .Y(\u0/N40 ) );
  XOR2X1 \u0/U373  ( .A(w0[22]), .B(\u0/subword [22]), .Y(\u0/N19 ) );
  XOR2X1 \u0/U368  ( .A(w0[21]), .B(\u0/subword [21]), .Y(\u0/N20 ) );
  XOR2X1 \u0/U358  ( .A(w0[19]), .B(\u0/subword [19]), .Y(\u0/N22 ) );
  XOR2X1 \u0/U348  ( .A(w0[17]), .B(\u0/subword [17]), .Y(\u0/N24 ) );
  XOR2X1 \u0/U333  ( .A(w0[14]), .B(\u0/subword [14]), .Y(\u0/N27 ) );
  XOR2X1 \u0/U328  ( .A(w0[13]), .B(\u0/subword [13]), .Y(\u0/N28 ) );
  XOR2X1 \u0/U318  ( .A(w0[11]), .B(\u0/subword [11]), .Y(\u0/N30 ) );
  XOR2X1 \u0/U308  ( .A(w0[9]), .B(\u0/subword [9]), .Y(\u0/N32 ) );
  XOR2X1 \u0/U263  ( .A(w0[0]), .B(\u0/subword [0]), .Y(\u0/N41 ) );
  XOR2X1 \u0/U343  ( .A(w0[16]), .B(\u0/subword [16]), .Y(\u0/N25 ) );
  XOR2X1 \u0/U303  ( .A(w0[8]), .B(\u0/subword [8]), .Y(\u0/N33 ) );
  XOR2X1 \u0/U417  ( .A(w1[31]), .B(\u0/N10 ), .Y(\u0/N76 ) );
  XOR2X1 \u0/U412  ( .A(w1[30]), .B(\u0/N11 ), .Y(\u0/N77 ) );
  XOR2X1 \u0/U407  ( .A(w1[29]), .B(\u0/N12 ), .Y(\u0/N78 ) );
  XOR2X1 \u0/U402  ( .A(w1[28]), .B(\u0/N13 ), .Y(\u0/N79 ) );
  XOR2X1 \u0/U397  ( .A(w1[27]), .B(\u0/N14 ), .Y(\u0/N80 ) );
  XOR2X1 \u0/U392  ( .A(w1[26]), .B(\u0/N15 ), .Y(\u0/N81 ) );
  XOR2X1 \u0/U387  ( .A(w1[25]), .B(\u0/N16 ), .Y(\u0/N82 ) );
  XOR2X1 \u0/U382  ( .A(w1[24]), .B(\u0/N17 ), .Y(\u0/N83 ) );
  XOR2X1 \u0/U281  ( .A(w2[4]), .B(\u0/N103 ), .Y(\u0/N169 ) );
  XOR2X1 \u0/U271  ( .A(w2[2]), .B(\u0/N105 ), .Y(\u0/N171 ) );
  XOR2X1 \u0/U361  ( .A(w2[20]), .B(\u0/N87 ), .Y(\u0/N153 ) );
  XOR2X1 \u0/U351  ( .A(w2[18]), .B(\u0/N89 ), .Y(\u0/N155 ) );
  XOR2X1 \u0/U321  ( .A(w2[12]), .B(\u0/N95 ), .Y(\u0/N161 ) );
  XOR2X1 \u0/U311  ( .A(w2[10]), .B(\u0/N97 ), .Y(\u0/N163 ) );
  XOR2X1 \u0/U337  ( .A(w1[15]), .B(\u0/N26 ), .Y(\u0/N92 ) );
  XOR2X1 \u0/U377  ( .A(w1[23]), .B(\u0/N18 ), .Y(\u0/N84 ) );
  XOR2X1 \u0/U297  ( .A(w1[7]), .B(\u0/N34 ), .Y(\u0/N100 ) );
  XOR2X1 \u0/U292  ( .A(w1[6]), .B(\u0/N35 ), .Y(\u0/N101 ) );
  XOR2X1 \u0/U287  ( .A(w1[5]), .B(\u0/N36 ), .Y(\u0/N102 ) );
  XOR2X1 \u0/U282  ( .A(w1[4]), .B(\u0/N37 ), .Y(\u0/N103 ) );
  XOR2X1 \u0/U277  ( .A(w1[3]), .B(\u0/N38 ), .Y(\u0/N104 ) );
  XOR2X1 \u0/U272  ( .A(w1[2]), .B(\u0/N39 ), .Y(\u0/N105 ) );
  XOR2X1 \u0/U267  ( .A(w1[1]), .B(\u0/N40 ), .Y(\u0/N106 ) );
  XOR2X1 \u0/U262  ( .A(w1[0]), .B(\u0/N41 ), .Y(\u0/N107 ) );
  XOR2X1 \u0/U372  ( .A(w1[22]), .B(\u0/N19 ), .Y(\u0/N85 ) );
  XOR2X1 \u0/U367  ( .A(w1[21]), .B(\u0/N20 ), .Y(\u0/N86 ) );
  XOR2X1 \u0/U362  ( .A(w1[20]), .B(\u0/N21 ), .Y(\u0/N87 ) );
  XOR2X1 \u0/U357  ( .A(w1[19]), .B(\u0/N22 ), .Y(\u0/N88 ) );
  XOR2X1 \u0/U352  ( .A(w1[18]), .B(\u0/N23 ), .Y(\u0/N89 ) );
  XOR2X1 \u0/U347  ( .A(w1[17]), .B(\u0/N24 ), .Y(\u0/N90 ) );
  XOR2X1 \u0/U342  ( .A(w1[16]), .B(\u0/N25 ), .Y(\u0/N91 ) );
  XOR2X1 \u0/U332  ( .A(w1[14]), .B(\u0/N27 ), .Y(\u0/N93 ) );
  XOR2X1 \u0/U327  ( .A(w1[13]), .B(\u0/N28 ), .Y(\u0/N94 ) );
  XOR2X1 \u0/U322  ( .A(w1[12]), .B(\u0/N29 ), .Y(\u0/N95 ) );
  XOR2X1 \u0/U317  ( .A(w1[11]), .B(\u0/N30 ), .Y(\u0/N96 ) );
  XOR2X1 \u0/U312  ( .A(w1[10]), .B(\u0/N31 ), .Y(\u0/N97 ) );
  XOR2X1 \u0/U307  ( .A(w1[9]), .B(\u0/N32 ), .Y(\u0/N98 ) );
  XOR2X1 \u0/U302  ( .A(w1[8]), .B(\u0/N33 ), .Y(\u0/N99 ) );
  XOR2X1 \u0/U336  ( .A(w2[15]), .B(\u0/N92 ), .Y(\u0/N158 ) );
  XOR2X1 \u0/U376  ( .A(w2[23]), .B(\u0/N84 ), .Y(\u0/N150 ) );
  XOR2X1 \u0/U416  ( .A(w2[31]), .B(\u0/N76 ), .Y(\u0/N142 ) );
  XOR2X1 \u0/U296  ( .A(w2[7]), .B(\u0/N100 ), .Y(\u0/N166 ) );
  XOR2X1 \u0/U291  ( .A(w2[6]), .B(\u0/N101 ), .Y(\u0/N167 ) );
  XOR2X1 \u0/U286  ( .A(w2[5]), .B(\u0/N102 ), .Y(\u0/N168 ) );
  XOR2X1 \u0/U276  ( .A(w2[3]), .B(\u0/N104 ), .Y(\u0/N170 ) );
  XOR2X1 \u0/U266  ( .A(w2[1]), .B(\u0/N106 ), .Y(\u0/N172 ) );
  XOR2X1 \u0/U261  ( .A(w2[0]), .B(\u0/N107 ), .Y(\u0/N173 ) );
  XOR2X1 \u0/U411  ( .A(w2[30]), .B(\u0/N77 ), .Y(\u0/N143 ) );
  XOR2X1 \u0/U406  ( .A(w2[29]), .B(\u0/N78 ), .Y(\u0/N144 ) );
  XOR2X1 \u0/U401  ( .A(w2[28]), .B(\u0/N79 ), .Y(\u0/N145 ) );
  XOR2X1 \u0/U396  ( .A(w2[27]), .B(\u0/N80 ), .Y(\u0/N146 ) );
  XOR2X1 \u0/U391  ( .A(w2[26]), .B(\u0/N81 ), .Y(\u0/N147 ) );
  XOR2X1 \u0/U386  ( .A(w2[25]), .B(\u0/N82 ), .Y(\u0/N148 ) );
  XOR2X1 \u0/U381  ( .A(w2[24]), .B(\u0/N83 ), .Y(\u0/N149 ) );
  XOR2X1 \u0/U371  ( .A(w2[22]), .B(\u0/N85 ), .Y(\u0/N151 ) );
  XOR2X1 \u0/U366  ( .A(w2[21]), .B(\u0/N86 ), .Y(\u0/N152 ) );
  XOR2X1 \u0/U356  ( .A(w2[19]), .B(\u0/N88 ), .Y(\u0/N154 ) );
  XOR2X1 \u0/U346  ( .A(w2[17]), .B(\u0/N90 ), .Y(\u0/N156 ) );
  XOR2X1 \u0/U341  ( .A(w2[16]), .B(\u0/N91 ), .Y(\u0/N157 ) );
  XOR2X1 \u0/U331  ( .A(w2[14]), .B(\u0/N93 ), .Y(\u0/N159 ) );
  XOR2X1 \u0/U326  ( .A(w2[13]), .B(\u0/N94 ), .Y(\u0/N160 ) );
  XOR2X1 \u0/U316  ( .A(w2[11]), .B(\u0/N96 ), .Y(\u0/N162 ) );
  XOR2X1 \u0/U306  ( .A(w2[9]), .B(\u0/N98 ), .Y(\u0/N164 ) );
  XOR2X1 \u0/U301  ( .A(w2[8]), .B(\u0/N99 ), .Y(\u0/N165 ) );
  XOR2X1 \u0/U419  ( .A(\u0/rcon [31]), .B(\u0/n258 ), .Y(\u0/N10 ) );
  XOR2X1 \u0/U418  ( .A(w0[31]), .B(\u0/subword [31]), .Y(\u0/n258 ) );
  XOR2X1 \u0/U414  ( .A(\u0/rcon [30]), .B(\u0/n259 ), .Y(\u0/N11 ) );
  XOR2X1 \u0/U413  ( .A(w0[30]), .B(\u0/subword [30]), .Y(\u0/n259 ) );
  XOR2X1 \u0/U409  ( .A(\u0/rcon [29]), .B(\u0/n260 ), .Y(\u0/N12 ) );
  XOR2X1 \u0/U408  ( .A(w0[29]), .B(\u0/subword [29]), .Y(\u0/n260 ) );
  XOR2X1 \u0/U399  ( .A(\u0/rcon [27]), .B(\u0/n262 ), .Y(\u0/N14 ) );
  XOR2X1 \u0/U398  ( .A(w0[27]), .B(\u0/subword [27]), .Y(\u0/n262 ) );
  XOR2X1 \u0/U389  ( .A(\u0/rcon [25]), .B(\u0/n264 ), .Y(\u0/N16 ) );
  XOR2X1 \u0/U388  ( .A(w0[25]), .B(\u0/subword [25]), .Y(\u0/n264 ) );
  XOR2X1 \u0/U384  ( .A(\u0/rcon [24]), .B(\u0/n265 ), .Y(\u0/N17 ) );
  XOR2X1 \u0/U383  ( .A(w0[24]), .B(\u0/subword [24]), .Y(\u0/n265 ) );
  XOR2X1 \u0/U404  ( .A(\u0/rcon [28]), .B(\u0/n261 ), .Y(\u0/N13 ) );
  XOR2X1 \u0/U403  ( .A(w0[28]), .B(\u0/subword [28]), .Y(\u0/n261 ) );
  XOR2X1 \u0/U394  ( .A(\u0/rcon [26]), .B(\u0/n263 ), .Y(\u0/N15 ) );
  XOR2X1 \u0/U393  ( .A(w0[26]), .B(\u0/subword [26]), .Y(\u0/n263 ) );
  XOR2X1 \u0/U295  ( .A(w3[7]), .B(\u0/N166 ), .Y(\u0/N232 ) );
  XOR2X1 \u0/U290  ( .A(w3[6]), .B(\u0/N167 ), .Y(\u0/N233 ) );
  XOR2X1 \u0/U285  ( .A(w3[5]), .B(\u0/N168 ), .Y(\u0/N234 ) );
  XOR2X1 \u0/U280  ( .A(w3[4]), .B(\u0/N169 ), .Y(\u0/N235 ) );
  XOR2X1 \u0/U275  ( .A(w3[3]), .B(\u0/N170 ), .Y(\u0/N236 ) );
  XOR2X1 \u0/U270  ( .A(w3[2]), .B(\u0/N171 ), .Y(\u0/N237 ) );
  XOR2X1 \u0/U265  ( .A(w3[1]), .B(\u0/N172 ), .Y(\u0/N238 ) );
  XOR2X1 \u0/U415  ( .A(w3[31]), .B(\u0/N142 ), .Y(\u0/N208 ) );
  XOR2X1 \u0/U410  ( .A(w3[30]), .B(\u0/N143 ), .Y(\u0/N209 ) );
  XOR2X1 \u0/U405  ( .A(w3[29]), .B(\u0/N144 ), .Y(\u0/N210 ) );
  XOR2X1 \u0/U400  ( .A(w3[28]), .B(\u0/N145 ), .Y(\u0/N211 ) );
  XOR2X1 \u0/U395  ( .A(w3[27]), .B(\u0/N146 ), .Y(\u0/N212 ) );
  XOR2X1 \u0/U390  ( .A(w3[26]), .B(\u0/N147 ), .Y(\u0/N213 ) );
  XOR2X1 \u0/U385  ( .A(w3[25]), .B(\u0/N148 ), .Y(\u0/N214 ) );
  XOR2X1 \u0/U380  ( .A(w3[24]), .B(\u0/N149 ), .Y(\u0/N215 ) );
  XOR2X1 \u0/U375  ( .A(w3[23]), .B(\u0/N150 ), .Y(\u0/N216 ) );
  XOR2X1 \u0/U370  ( .A(w3[22]), .B(\u0/N151 ), .Y(\u0/N217 ) );
  XOR2X1 \u0/U365  ( .A(w3[21]), .B(\u0/N152 ), .Y(\u0/N218 ) );
  XOR2X1 \u0/U360  ( .A(w3[20]), .B(\u0/N153 ), .Y(\u0/N219 ) );
  XOR2X1 \u0/U355  ( .A(w3[19]), .B(\u0/N154 ), .Y(\u0/N220 ) );
  XOR2X1 \u0/U350  ( .A(w3[18]), .B(\u0/N155 ), .Y(\u0/N221 ) );
  XOR2X1 \u0/U345  ( .A(w3[17]), .B(\u0/N156 ), .Y(\u0/N222 ) );
  XOR2X1 \u0/U340  ( .A(w3[16]), .B(\u0/N157 ), .Y(\u0/N223 ) );
  XOR2X1 \u0/U335  ( .A(w3[15]), .B(\u0/N158 ), .Y(\u0/N224 ) );
  XOR2X1 \u0/U330  ( .A(w3[14]), .B(\u0/N159 ), .Y(\u0/N225 ) );
  XOR2X1 \u0/U325  ( .A(w3[13]), .B(\u0/N160 ), .Y(\u0/N226 ) );
  XOR2X1 \u0/U320  ( .A(w3[12]), .B(\u0/N161 ), .Y(\u0/N227 ) );
  XOR2X1 \u0/U315  ( .A(w3[11]), .B(\u0/N162 ), .Y(\u0/N228 ) );
  XOR2X1 \u0/U310  ( .A(w3[10]), .B(\u0/N163 ), .Y(\u0/N229 ) );
  XOR2X1 \u0/U305  ( .A(w3[9]), .B(\u0/N164 ), .Y(\u0/N230 ) );
  XOR2X1 \u0/U300  ( .A(w3[8]), .B(\u0/N165 ), .Y(\u0/N231 ) );
  XOR2X1 \u0/U260  ( .A(w3[0]), .B(\u0/N173 ), .Y(\u0/N239 ) );
  DFFHQX2 \u0/w_reg[3][1]  ( .D(\u0/n124 ), .CK(clk), .Q(w3[1]) );
  DFFHQX2 \u0/w_reg[3][25]  ( .D(\u0/n28 ), .CK(clk), .Q(w3[25]) );
  DFFHQX2 \u0/w_reg[3][17]  ( .D(\u0/n60 ), .CK(clk), .Q(w3[17]) );
  DFFHQX2 \u0/w_reg[3][9]  ( .D(\u0/n92 ), .CK(clk), .Q(w3[9]) );
  DFFHQX1 \u0/w_reg[3][4]  ( .D(\u0/n112 ), .CK(clk), .Q(w3[4]) );
  DFFHQX1 \u0/w_reg[3][28]  ( .D(\u0/n16 ), .CK(clk), .Q(w3[28]) );
  DFFHQX1 \u0/w_reg[3][20]  ( .D(\u0/n48 ), .CK(clk), .Q(w3[20]) );
  DFFHQX1 \u0/w_reg[3][12]  ( .D(\u0/n80 ), .CK(clk), .Q(w3[12]) );
  DFFHQX1 \u0/w_reg[3][2]  ( .D(\u0/n120 ), .CK(clk), .Q(w3[2]) );
  DFFHQX1 \u0/w_reg[3][26]  ( .D(\u0/n24 ), .CK(clk), .Q(w3[26]) );
  DFFHQX1 \u0/w_reg[3][18]  ( .D(\u0/n56 ), .CK(clk), .Q(w3[18]) );
  DFFHQX1 \u0/w_reg[3][10]  ( .D(\u0/n88 ), .CK(clk), .Q(w3[10]) );
  DFFHQX1 \u0/w_reg[3][3]  ( .D(\u0/n116 ), .CK(clk), .Q(w3[3]) );
  DFFHQX1 \u0/w_reg[3][27]  ( .D(\u0/n20 ), .CK(clk), .Q(w3[27]) );
  DFFHQX1 \u0/w_reg[3][19]  ( .D(\u0/n52 ), .CK(clk), .Q(w3[19]) );
  DFFHQX1 \u0/w_reg[3][11]  ( .D(\u0/n84 ), .CK(clk), .Q(w3[11]) );
  DFFHQX1 \u0/w_reg[3][5]  ( .D(\u0/n108 ), .CK(clk), .Q(w3[5]) );
  DFFHQX1 \u0/w_reg[3][29]  ( .D(\u0/n12 ), .CK(clk), .Q(w3[29]) );
  DFFHQX1 \u0/w_reg[3][21]  ( .D(\u0/n44 ), .CK(clk), .Q(w3[21]) );
  DFFHQX1 \u0/w_reg[3][13]  ( .D(\u0/n76 ), .CK(clk), .Q(w3[13]) );
  DFFHQX1 \u0/w_reg[3][7]  ( .D(\u0/n100 ), .CK(clk), .Q(w3[7]) );
  DFFHQX1 \u0/w_reg[3][31]  ( .D(\u0/n4 ), .CK(clk), .Q(w3[31]) );
  DFFHQX1 \u0/w_reg[3][23]  ( .D(\u0/n36 ), .CK(clk), .Q(w3[23]) );
  DFFHQX1 \u0/w_reg[3][15]  ( .D(\u0/n68 ), .CK(clk), .Q(w3[15]) );
  DFFHQX1 \u0/w_reg[3][24]  ( .D(\u0/n32 ), .CK(clk), .Q(w3[24]) );
  DFFHQX1 \u0/w_reg[3][16]  ( .D(\u0/n64 ), .CK(clk), .Q(w3[16]) );
  DFFHQX1 \u0/w_reg[3][8]  ( .D(\u0/n96 ), .CK(clk), .Q(w3[8]) );
  DFFHQX1 \u0/w_reg[3][0]  ( .D(\u0/n128 ), .CK(clk), .Q(w3[0]) );
  DFFHQX1 \u0/w_reg[0][15]  ( .D(\u0/n65 ), .CK(clk), .Q(w0[15]) );
  DFFHQX1 \u0/w_reg[1][15]  ( .D(\u0/n66 ), .CK(clk), .Q(w1[15]) );
  DFFHQX1 \u0/w_reg[2][15]  ( .D(\u0/n67 ), .CK(clk), .Q(w2[15]) );
  DFFHQX1 \u0/w_reg[0][23]  ( .D(\u0/n33 ), .CK(clk), .Q(w0[23]) );
  DFFHQX1 \u0/w_reg[1][23]  ( .D(\u0/n34 ), .CK(clk), .Q(w1[23]) );
  DFFHQX1 \u0/w_reg[2][23]  ( .D(\u0/n35 ), .CK(clk), .Q(w2[23]) );
  DFFHQX1 \u0/w_reg[0][31]  ( .D(\u0/n1 ), .CK(clk), .Q(w0[31]) );
  DFFHQX1 \u0/w_reg[1][31]  ( .D(\u0/n2 ), .CK(clk), .Q(w1[31]) );
  DFFHQX1 \u0/w_reg[2][31]  ( .D(\u0/n3 ), .CK(clk), .Q(w2[31]) );
  DFFHQX1 \u0/w_reg[0][7]  ( .D(\u0/n97 ), .CK(clk), .Q(w0[7]) );
  DFFHQX1 \u0/w_reg[1][7]  ( .D(\u0/n98 ), .CK(clk), .Q(w1[7]) );
  DFFHQX1 \u0/w_reg[2][7]  ( .D(\u0/n99 ), .CK(clk), .Q(w2[7]) );
  DFFHQX1 \u0/w_reg[0][6]  ( .D(\u0/n101 ), .CK(clk), .Q(w0[6]) );
  DFFHQX1 \u0/w_reg[1][6]  ( .D(\u0/n102 ), .CK(clk), .Q(w1[6]) );
  DFFHQX1 \u0/w_reg[2][6]  ( .D(\u0/n103 ), .CK(clk), .Q(w2[6]) );
  DFFHQX1 \u0/w_reg[0][5]  ( .D(\u0/n105 ), .CK(clk), .Q(w0[5]) );
  DFFHQX1 \u0/w_reg[1][5]  ( .D(\u0/n106 ), .CK(clk), .Q(w1[5]) );
  DFFHQX1 \u0/w_reg[2][5]  ( .D(\u0/n107 ), .CK(clk), .Q(w2[5]) );
  DFFHQX1 \u0/w_reg[0][4]  ( .D(\u0/n109 ), .CK(clk), .Q(w0[4]) );
  DFFHQX1 \u0/w_reg[1][4]  ( .D(\u0/n110 ), .CK(clk), .Q(w1[4]) );
  DFFHQX1 \u0/w_reg[2][4]  ( .D(\u0/n111 ), .CK(clk), .Q(w2[4]) );
  DFFHQX1 \u0/w_reg[0][3]  ( .D(\u0/n113 ), .CK(clk), .Q(w0[3]) );
  DFFHQX1 \u0/w_reg[1][3]  ( .D(\u0/n114 ), .CK(clk), .Q(w1[3]) );
  DFFHQX1 \u0/w_reg[2][3]  ( .D(\u0/n115 ), .CK(clk), .Q(w2[3]) );
  DFFHQX1 \u0/w_reg[0][2]  ( .D(\u0/n117 ), .CK(clk), .Q(w0[2]) );
  DFFHQX1 \u0/w_reg[1][2]  ( .D(\u0/n118 ), .CK(clk), .Q(w1[2]) );
  DFFHQX1 \u0/w_reg[2][2]  ( .D(\u0/n119 ), .CK(clk), .Q(w2[2]) );
  DFFHQX1 \u0/w_reg[0][1]  ( .D(\u0/n121 ), .CK(clk), .Q(w0[1]) );
  DFFHQX1 \u0/w_reg[1][1]  ( .D(\u0/n122 ), .CK(clk), .Q(w1[1]) );
  DFFHQX1 \u0/w_reg[2][1]  ( .D(\u0/n123 ), .CK(clk), .Q(w2[1]) );
  DFFHQX1 \u0/w_reg[0][0]  ( .D(\u0/n125 ), .CK(clk), .Q(w0[0]) );
  DFFHQX1 \u0/w_reg[1][0]  ( .D(\u0/n126 ), .CK(clk), .Q(w1[0]) );
  DFFHQX1 \u0/w_reg[2][0]  ( .D(\u0/n127 ), .CK(clk), .Q(w2[0]) );
  DFFHQX1 \u0/w_reg[0][30]  ( .D(\u0/n5 ), .CK(clk), .Q(w0[30]) );
  DFFHQX1 \u0/w_reg[1][30]  ( .D(\u0/n6 ), .CK(clk), .Q(w1[30]) );
  DFFHQX1 \u0/w_reg[2][30]  ( .D(\u0/n7 ), .CK(clk), .Q(w2[30]) );
  DFFHQX1 \u0/w_reg[0][29]  ( .D(\u0/n9 ), .CK(clk), .Q(w0[29]) );
  DFFHQX1 \u0/w_reg[1][29]  ( .D(\u0/n10 ), .CK(clk), .Q(w1[29]) );
  DFFHQX1 \u0/w_reg[2][29]  ( .D(\u0/n11 ), .CK(clk), .Q(w2[29]) );
  DFFHQX1 \u0/w_reg[0][28]  ( .D(\u0/n13 ), .CK(clk), .Q(w0[28]) );
  DFFHQX1 \u0/w_reg[1][28]  ( .D(\u0/n14 ), .CK(clk), .Q(w1[28]) );
  DFFHQX1 \u0/w_reg[2][28]  ( .D(\u0/n15 ), .CK(clk), .Q(w2[28]) );
  DFFHQX1 \u0/w_reg[0][27]  ( .D(\u0/n17 ), .CK(clk), .Q(w0[27]) );
  DFFHQX1 \u0/w_reg[1][27]  ( .D(\u0/n18 ), .CK(clk), .Q(w1[27]) );
  DFFHQX1 \u0/w_reg[2][27]  ( .D(\u0/n19 ), .CK(clk), .Q(w2[27]) );
  DFFHQX1 \u0/w_reg[0][26]  ( .D(\u0/n21 ), .CK(clk), .Q(w0[26]) );
  DFFHQX1 \u0/w_reg[1][26]  ( .D(\u0/n22 ), .CK(clk), .Q(w1[26]) );
  DFFHQX1 \u0/w_reg[2][26]  ( .D(\u0/n23 ), .CK(clk), .Q(w2[26]) );
  DFFHQX1 \u0/w_reg[0][25]  ( .D(\u0/n25 ), .CK(clk), .Q(w0[25]) );
  DFFHQX1 \u0/w_reg[1][25]  ( .D(\u0/n26 ), .CK(clk), .Q(w1[25]) );
  DFFHQX1 \u0/w_reg[2][25]  ( .D(\u0/n27 ), .CK(clk), .Q(w2[25]) );
  DFFHQX1 \u0/w_reg[0][24]  ( .D(\u0/n29 ), .CK(clk), .Q(w0[24]) );
  DFFHQX1 \u0/w_reg[1][24]  ( .D(\u0/n30 ), .CK(clk), .Q(w1[24]) );
  DFFHQX1 \u0/w_reg[2][24]  ( .D(\u0/n31 ), .CK(clk), .Q(w2[24]) );
  DFFHQX1 \u0/w_reg[0][22]  ( .D(\u0/n37 ), .CK(clk), .Q(w0[22]) );
  DFFHQX1 \u0/w_reg[1][22]  ( .D(\u0/n38 ), .CK(clk), .Q(w1[22]) );
  DFFHQX1 \u0/w_reg[2][22]  ( .D(\u0/n39 ), .CK(clk), .Q(w2[22]) );
  DFFHQX1 \u0/w_reg[0][21]  ( .D(\u0/n41 ), .CK(clk), .Q(w0[21]) );
  DFFHQX1 \u0/w_reg[1][21]  ( .D(\u0/n42 ), .CK(clk), .Q(w1[21]) );
  DFFHQX1 \u0/w_reg[2][21]  ( .D(\u0/n43 ), .CK(clk), .Q(w2[21]) );
  DFFHQX1 \u0/w_reg[0][20]  ( .D(\u0/n45 ), .CK(clk), .Q(w0[20]) );
  DFFHQX1 \u0/w_reg[1][20]  ( .D(\u0/n46 ), .CK(clk), .Q(w1[20]) );
  DFFHQX1 \u0/w_reg[2][20]  ( .D(\u0/n47 ), .CK(clk), .Q(w2[20]) );
  DFFHQX1 \u0/w_reg[0][19]  ( .D(\u0/n49 ), .CK(clk), .Q(w0[19]) );
  DFFHQX1 \u0/w_reg[1][19]  ( .D(\u0/n50 ), .CK(clk), .Q(w1[19]) );
  DFFHQX1 \u0/w_reg[2][19]  ( .D(\u0/n51 ), .CK(clk), .Q(w2[19]) );
  DFFHQX1 \u0/w_reg[0][18]  ( .D(\u0/n53 ), .CK(clk), .Q(w0[18]) );
  DFFHQX1 \u0/w_reg[1][18]  ( .D(\u0/n54 ), .CK(clk), .Q(w1[18]) );
  DFFHQX1 \u0/w_reg[2][18]  ( .D(\u0/n55 ), .CK(clk), .Q(w2[18]) );
  DFFHQX1 \u0/w_reg[0][17]  ( .D(\u0/n57 ), .CK(clk), .Q(w0[17]) );
  DFFHQX1 \u0/w_reg[1][17]  ( .D(\u0/n58 ), .CK(clk), .Q(w1[17]) );
  DFFHQX1 \u0/w_reg[2][17]  ( .D(\u0/n59 ), .CK(clk), .Q(w2[17]) );
  DFFHQX1 \u0/w_reg[0][16]  ( .D(\u0/n61 ), .CK(clk), .Q(w0[16]) );
  DFFHQX1 \u0/w_reg[1][16]  ( .D(\u0/n62 ), .CK(clk), .Q(w1[16]) );
  DFFHQX1 \u0/w_reg[2][16]  ( .D(\u0/n63 ), .CK(clk), .Q(w2[16]) );
  DFFHQX1 \u0/w_reg[0][14]  ( .D(\u0/n69 ), .CK(clk), .Q(w0[14]) );
  DFFHQX1 \u0/w_reg[1][14]  ( .D(\u0/n70 ), .CK(clk), .Q(w1[14]) );
  DFFHQX1 \u0/w_reg[2][14]  ( .D(\u0/n71 ), .CK(clk), .Q(w2[14]) );
  DFFHQX1 \u0/w_reg[0][13]  ( .D(\u0/n73 ), .CK(clk), .Q(w0[13]) );
  DFFHQX1 \u0/w_reg[1][13]  ( .D(\u0/n74 ), .CK(clk), .Q(w1[13]) );
  DFFHQX1 \u0/w_reg[2][13]  ( .D(\u0/n75 ), .CK(clk), .Q(w2[13]) );
  DFFHQX1 \u0/w_reg[0][12]  ( .D(\u0/n77 ), .CK(clk), .Q(w0[12]) );
  DFFHQX1 \u0/w_reg[1][12]  ( .D(\u0/n78 ), .CK(clk), .Q(w1[12]) );
  DFFHQX1 \u0/w_reg[2][12]  ( .D(\u0/n79 ), .CK(clk), .Q(w2[12]) );
  DFFHQX1 \u0/w_reg[0][11]  ( .D(\u0/n81 ), .CK(clk), .Q(w0[11]) );
  DFFHQX1 \u0/w_reg[1][11]  ( .D(\u0/n82 ), .CK(clk), .Q(w1[11]) );
  DFFHQX1 \u0/w_reg[2][11]  ( .D(\u0/n83 ), .CK(clk), .Q(w2[11]) );
  DFFHQX1 \u0/w_reg[0][10]  ( .D(\u0/n85 ), .CK(clk), .Q(w0[10]) );
  DFFHQX1 \u0/w_reg[1][10]  ( .D(\u0/n86 ), .CK(clk), .Q(w1[10]) );
  DFFHQX1 \u0/w_reg[2][10]  ( .D(\u0/n87 ), .CK(clk), .Q(w2[10]) );
  DFFHQX1 \u0/w_reg[0][9]  ( .D(\u0/n89 ), .CK(clk), .Q(w0[9]) );
  DFFHQX1 \u0/w_reg[1][9]  ( .D(\u0/n90 ), .CK(clk), .Q(w1[9]) );
  DFFHQX1 \u0/w_reg[2][9]  ( .D(\u0/n91 ), .CK(clk), .Q(w2[9]) );
  DFFHQX1 \u0/w_reg[0][8]  ( .D(\u0/n93 ), .CK(clk), .Q(w0[8]) );
  DFFHQX1 \u0/w_reg[1][8]  ( .D(\u0/n94 ), .CK(clk), .Q(w1[8]) );
  DFFHQX1 \u0/w_reg[2][8]  ( .D(\u0/n95 ), .CK(clk), .Q(w2[8]) );
  aes_rcon \u0/r0  ( .clk(clk), .kld(ld), .out(\u0/rcon ) );
  aes_sbox_1 \u0/u3  ( .a(w3[31:24]), .d(\u0/subword [7:0]) );
  aes_sbox_2 \u0/u2  ( .a(w3[7:0]), .d(\u0/subword [15:8]) );
  aes_sbox_3 \u0/u1  ( .a(w3[15:8]), .d(\u0/subword [23:16]) );
  aes_sbox_4 \u0/u0  ( .a(w3[23:16]), .d(\u0/subword [31:24]) );
  NAND2X1 \us00/U366  ( .A(\us00/n47 ), .B(\us00/n226 ), .Y(\us00/n189 ) );
  NOR2X1 \us00/U365  ( .A(\us00/n226 ), .B(sa00[3]), .Y(\us00/n242 ) );
  INVX1 \us00/U364  ( .A(\us00/n242 ), .Y(\us00/n205 ) );
  AND2X1 \us00/U363  ( .A(\us00/n189 ), .B(\us00/n205 ), .Y(\us00/n65 ) );
  NOR2X1 \us00/U362  ( .A(\us00/n226 ), .B(\us00/n47 ), .Y(\us00/n45 ) );
  NOR2X1 \us00/U361  ( .A(\us00/n259 ), .B(\us00/n45 ), .Y(\us00/n73 ) );
  NAND2BX1 \us00/U360  ( .AN(\us00/n73 ), .B(\us00/n6 ), .Y(\us00/n158 ) );
  NOR2X1 \us00/U359  ( .A(\us00/n226 ), .B(\us00/n159 ), .Y(\us00/n95 ) );
  INVX1 \us00/U358  ( .A(\us00/n95 ), .Y(\us00/n111 ) );
  NOR2X1 \us00/U357  ( .A(\us00/n145 ), .B(sa00[1]), .Y(\us00/n42 ) );
  INVX1 \us00/U356  ( .A(\us00/n42 ), .Y(\us00/n121 ) );
  INVX1 \us00/U355  ( .A(\us00/n47 ), .Y(\us00/n96 ) );
  OAI211X1 \us00/U354  ( .A0(\us00/n65 ), .A1(\us00/n27 ), .B0(\us00/n158 ), 
        .C0(\us00/n358 ), .Y(\us00/n355 ) );
  NOR2X1 \us00/U353  ( .A(\us00/n226 ), .B(\us00/n145 ), .Y(\us00/n59 ) );
  NOR2X1 \us00/U352  ( .A(\us00/n96 ), .B(\us00/n59 ), .Y(\us00/n271 ) );
  NOR2X1 \us00/U351  ( .A(\us00/n226 ), .B(\us00/n278 ), .Y(\us00/n217 ) );
  INVX1 \us00/U350  ( .A(\us00/n217 ), .Y(\us00/n150 ) );
  NAND2X1 \us00/U349  ( .A(\us00/n44 ), .B(\us00/n150 ), .Y(\us00/n147 ) );
  NAND2X1 \us00/U348  ( .A(sa00[4]), .B(\us00/n226 ), .Y(\us00/n101 ) );
  INVX1 \us00/U347  ( .A(\us00/n159 ), .Y(\us00/n188 ) );
  NOR2X1 \us00/U346  ( .A(\us00/n188 ), .B(\us00/n226 ), .Y(\us00/n25 ) );
  INVX1 \us00/U345  ( .A(\us00/n172 ), .Y(\us00/n107 ) );
  AOI22X1 \us00/U344  ( .A0(\us00/n33 ), .A1(\us00/n147 ), .B0(\us00/n24 ), 
        .B1(\us00/n107 ), .Y(\us00/n357 ) );
  OAI221XL \us00/U343  ( .A0(\us00/n18 ), .A1(\us00/n121 ), .B0(\us00/n271 ), 
        .B1(\us00/n20 ), .C0(\us00/n357 ), .Y(\us00/n356 ) );
  MXI2X1 \us00/U342  ( .A(\us00/n355 ), .B(\us00/n356 ), .S0(\us00/n252 ), .Y(
        \us00/n331 ) );
  INVX1 \us00/U341  ( .A(\us00/n59 ), .Y(\us00/n79 ) );
  AND2X1 \us00/U340  ( .A(\us00/n101 ), .B(\us00/n79 ), .Y(\us00/n325 ) );
  XNOR2X1 \us00/U339  ( .A(sa00[5]), .B(\us00/n226 ), .Y(\us00/n352 ) );
  NOR2X1 \us00/U338  ( .A(\us00/n226 ), .B(\us00/n136 ), .Y(\us00/n281 ) );
  INVX1 \us00/U337  ( .A(\us00/n281 ), .Y(\us00/n19 ) );
  NAND2X1 \us00/U336  ( .A(\us00/n145 ), .B(\us00/n226 ), .Y(\us00/n223 ) );
  AOI21X1 \us00/U335  ( .A0(\us00/n19 ), .A1(\us00/n223 ), .B0(\us00/n27 ), 
        .Y(\us00/n354 ) );
  AOI31X1 \us00/U334  ( .A0(\us00/n6 ), .A1(\us00/n352 ), .A2(\us00/n259 ), 
        .B0(\us00/n354 ), .Y(\us00/n353 ) );
  OAI221XL \us00/U333  ( .A0(\us00/n20 ), .A1(\us00/n34 ), .B0(\us00/n325 ), 
        .B1(\us00/n4 ), .C0(\us00/n353 ), .Y(\us00/n347 ) );
  INVX1 \us00/U332  ( .A(\us00/n352 ), .Y(\us00/n349 ) );
  NAND2X1 \us00/U331  ( .A(\us00/n278 ), .B(\us00/n6 ), .Y(\us00/n74 ) );
  OAI211X1 \us00/U330  ( .A0(\us00/n349 ), .A1(\us00/n74 ), .B0(\us00/n350 ), 
        .C0(\us00/n351 ), .Y(\us00/n348 ) );
  MXI2X1 \us00/U329  ( .A(\us00/n347 ), .B(\us00/n348 ), .S0(\us00/n252 ), .Y(
        \us00/n332 ) );
  NOR2X1 \us00/U328  ( .A(\us00/n44 ), .B(\us00/n226 ), .Y(\us00/n157 ) );
  INVX1 \us00/U327  ( .A(\us00/n157 ), .Y(\us00/n240 ) );
  NAND2X1 \us00/U326  ( .A(\us00/n240 ), .B(\us00/n189 ), .Y(\us00/n68 ) );
  NOR2X1 \us00/U325  ( .A(\us00/n20 ), .B(\us00/n159 ), .Y(\us00/n225 ) );
  NOR2X1 \us00/U324  ( .A(\us00/n225 ), .B(\us00/n40 ), .Y(\us00/n345 ) );
  INVX1 \us00/U323  ( .A(\us00/n278 ), .Y(\us00/n94 ) );
  NAND2X1 \us00/U322  ( .A(\us00/n94 ), .B(\us00/n226 ), .Y(\us00/n199 ) );
  NAND2X1 \us00/U321  ( .A(\us00/n199 ), .B(\us00/n205 ), .Y(\us00/n82 ) );
  NAND2X1 \us00/U320  ( .A(\us00/n19 ), .B(\us00/n199 ), .Y(\us00/n295 ) );
  NOR2X1 \us00/U319  ( .A(\us00/n226 ), .B(\us00/n259 ), .Y(\us00/n210 ) );
  NOR2X1 \us00/U318  ( .A(\us00/n27 ), .B(\us00/n210 ), .Y(\us00/n173 ) );
  MXI2X1 \us00/U317  ( .A(\us00/n345 ), .B(\us00/n346 ), .S0(\us00/n252 ), .Y(
        \us00/n342 ) );
  NOR2X1 \us00/U316  ( .A(sa00[1]), .B(sa00[3]), .Y(\us00/n163 ) );
  INVX1 \us00/U315  ( .A(\us00/n163 ), .Y(\us00/n37 ) );
  INVX1 \us00/U314  ( .A(\us00/n173 ), .Y(\us00/n344 ) );
  AOI21X1 \us00/U313  ( .A0(\us00/n240 ), .A1(\us00/n37 ), .B0(\us00/n344 ), 
        .Y(\us00/n343 ) );
  AOI211X1 \us00/U312  ( .A0(\us00/n5 ), .A1(\us00/n68 ), .B0(\us00/n342 ), 
        .C0(\us00/n343 ), .Y(\us00/n333 ) );
  NOR2X1 \us00/U311  ( .A(\us00/n18 ), .B(\us00/n226 ), .Y(\us00/n258 ) );
  NAND2X1 \us00/U310  ( .A(\us00/n278 ), .B(sa00[1]), .Y(\us00/n204 ) );
  NOR2X1 \us00/U309  ( .A(\us00/n188 ), .B(sa00[1]), .Y(\us00/n179 ) );
  INVX1 \us00/U308  ( .A(\us00/n179 ), .Y(\us00/n330 ) );
  NAND2X1 \us00/U307  ( .A(\us00/n204 ), .B(\us00/n330 ), .Y(\us00/n239 ) );
  NOR2X1 \us00/U306  ( .A(\us00/n136 ), .B(sa00[1]), .Y(\us00/n299 ) );
  NOR2X1 \us00/U305  ( .A(\us00/n299 ), .B(\us00/n210 ), .Y(\us00/n341 ) );
  OAI32X1 \us00/U304  ( .A0(\us00/n27 ), .A1(\us00/n278 ), .A2(\us00/n95 ), 
        .B0(\us00/n341 ), .B1(\us00/n4 ), .Y(\us00/n340 ) );
  INVX1 \us00/U303  ( .A(\us00/n45 ), .Y(\us00/n126 ) );
  NAND2X1 \us00/U302  ( .A(\us00/n126 ), .B(\us00/n101 ), .Y(\us00/n178 ) );
  NOR2X1 \us00/U301  ( .A(\us00/n18 ), .B(\us00/n136 ), .Y(\us00/n280 ) );
  OAI21XL \us00/U300  ( .A0(\us00/n4 ), .A1(\us00/n121 ), .B0(\us00/n339 ), 
        .Y(\us00/n338 ) );
  MXI2X1 \us00/U299  ( .A(\us00/n336 ), .B(\us00/n337 ), .S0(\us00/n252 ), .Y(
        \us00/n335 ) );
  NOR2X1 \us00/U298  ( .A(\us00/n258 ), .B(\us00/n335 ), .Y(\us00/n334 ) );
  MX4X1 \us00/U297  ( .A(\us00/n331 ), .B(\us00/n332 ), .C(\us00/n333 ), .D(
        \us00/n334 ), .S0(sa00[6]), .S1(\us00/n234 ), .Y(sa00_sr[0]) );
  INVX1 \us00/U296  ( .A(\us00/n299 ), .Y(\us00/n80 ) );
  NOR2X1 \us00/U295  ( .A(\us00/n111 ), .B(\us00/n18 ), .Y(\us00/n269 ) );
  INVX1 \us00/U294  ( .A(\us00/n269 ), .Y(\us00/n75 ) );
  OAI221XL \us00/U293  ( .A0(\us00/n18 ), .A1(\us00/n330 ), .B0(\us00/n20 ), 
        .B1(\us00/n80 ), .C0(\us00/n75 ), .Y(\us00/n329 ) );
  AOI221X1 \us00/U292  ( .A0(\us00/n325 ), .A1(\us00/n33 ), .B0(\us00/n24 ), 
        .B1(\us00/n303 ), .C0(\us00/n329 ), .Y(\us00/n319 ) );
  NOR2X1 \us00/U291  ( .A(\us00/n234 ), .B(sa00[5]), .Y(\us00/n14 ) );
  NOR2X1 \us00/U290  ( .A(\us00/n25 ), .B(\us00/n299 ), .Y(\us00/n313 ) );
  NAND2X1 \us00/U289  ( .A(\us00/n44 ), .B(\us00/n226 ), .Y(\us00/n300 ) );
  AND2X1 \us00/U288  ( .A(\us00/n300 ), .B(\us00/n240 ), .Y(\us00/n23 ) );
  OAI32X1 \us00/U287  ( .A0(\us00/n4 ), .A1(\us00/n145 ), .A2(\us00/n210 ), 
        .B0(\us00/n137 ), .B1(\us00/n27 ), .Y(\us00/n328 ) );
  NOR2X1 \us00/U286  ( .A(sa00[0]), .B(sa00[5]), .Y(\us00/n16 ) );
  INVX1 \us00/U285  ( .A(\us00/n16 ), .Y(\us00/n114 ) );
  INVX1 \us00/U284  ( .A(\us00/n145 ), .Y(\us00/n149 ) );
  NOR2X1 \us00/U283  ( .A(\us00/n47 ), .B(sa00[1]), .Y(\us00/n98 ) );
  INVX1 \us00/U282  ( .A(\us00/n98 ), .Y(\us00/n284 ) );
  OAI21XL \us00/U281  ( .A0(\us00/n69 ), .A1(\us00/n284 ), .B0(\us00/n27 ), 
        .Y(\us00/n327 ) );
  AOI31X1 \us00/U280  ( .A0(\us00/n111 ), .A1(\us00/n149 ), .A2(\us00/n327 ), 
        .B0(\us00/n225 ), .Y(\us00/n326 ) );
  OAI21XL \us00/U279  ( .A0(\us00/n325 ), .A1(\us00/n18 ), .B0(\us00/n326 ), 
        .Y(\us00/n322 ) );
  NAND2X1 \us00/U278  ( .A(\us00/n19 ), .B(\us00/n189 ), .Y(\us00/n71 ) );
  NOR2X1 \us00/U277  ( .A(\us00/n71 ), .B(\us00/n18 ), .Y(\us00/n135 ) );
  AOI21X1 \us00/U276  ( .A0(\us00/n40 ), .A1(sa00[4]), .B0(\us00/n135 ), .Y(
        \us00/n324 ) );
  OAI221XL \us00/U275  ( .A0(\us00/n47 ), .A1(\us00/n27 ), .B0(\us00/n65 ), 
        .B1(\us00/n20 ), .C0(\us00/n324 ), .Y(\us00/n323 ) );
  AOI22X1 \us00/U274  ( .A0(\us00/n55 ), .A1(\us00/n322 ), .B0(\us00/n89 ), 
        .B1(\us00/n323 ), .Y(\us00/n321 ) );
  OAI221XL \us00/U273  ( .A0(\us00/n319 ), .A1(\us00/n52 ), .B0(\us00/n320 ), 
        .B1(\us00/n114 ), .C0(\us00/n321 ), .Y(\us00/n304 ) );
  NOR2X1 \us00/U272  ( .A(\us00/n226 ), .B(\us00/n58 ), .Y(\us00/n290 ) );
  INVX1 \us00/U271  ( .A(\us00/n290 ), .Y(\us00/n200 ) );
  NAND2X1 \us00/U270  ( .A(\us00/n34 ), .B(\us00/n200 ), .Y(\us00/n120 ) );
  INVX1 \us00/U269  ( .A(\us00/n210 ), .Y(\us00/n100 ) );
  OAI221XL \us00/U268  ( .A0(\us00/n20 ), .A1(\us00/n100 ), .B0(sa00[3]), .B1(
        \us00/n4 ), .C0(\us00/n262 ), .Y(\us00/n317 ) );
  INVX1 \us00/U267  ( .A(\us00/n258 ), .Y(\us00/n182 ) );
  AOI211X1 \us00/U266  ( .A0(\us00/n33 ), .A1(\us00/n120 ), .B0(\us00/n317 ), 
        .C0(\us00/n318 ), .Y(\us00/n306 ) );
  NAND2X1 \us00/U265  ( .A(\us00/n100 ), .B(\us00/n199 ), .Y(\us00/n151 ) );
  INVX1 \us00/U264  ( .A(\us00/n151 ), .Y(\us00/n314 ) );
  NOR2X1 \us00/U263  ( .A(\us00/n45 ), .B(\us00/n163 ), .Y(\us00/n160 ) );
  INVX1 \us00/U262  ( .A(\us00/n295 ), .Y(\us00/n92 ) );
  AOI21X1 \us00/U261  ( .A0(sa00[1]), .A1(\us00/n58 ), .B0(\us00/n98 ), .Y(
        \us00/n316 ) );
  OAI22X1 \us00/U260  ( .A0(\us00/n92 ), .A1(\us00/n18 ), .B0(\us00/n316 ), 
        .B1(\us00/n27 ), .Y(\us00/n315 ) );
  NOR2X1 \us00/U259  ( .A(\us00/n149 ), .B(\us00/n226 ), .Y(\us00/n41 ) );
  INVX1 \us00/U258  ( .A(\us00/n41 ), .Y(\us00/n105 ) );
  NAND2X1 \us00/U257  ( .A(\us00/n284 ), .B(\us00/n105 ), .Y(\us00/n227 ) );
  AOI21X1 \us00/U256  ( .A0(\us00/n313 ), .A1(\us00/n33 ), .B0(\us00/n269 ), 
        .Y(\us00/n312 ) );
  OAI221XL \us00/U255  ( .A0(\us00/n149 ), .A1(\us00/n20 ), .B0(\us00/n4 ), 
        .B1(\us00/n227 ), .C0(\us00/n312 ), .Y(\us00/n309 ) );
  AOI21X1 \us00/U254  ( .A0(\us00/n226 ), .A1(\us00/n188 ), .B0(\us00/n242 ), 
        .Y(\us00/n185 ) );
  INVX1 \us00/U253  ( .A(\us00/n185 ), .Y(\us00/n48 ) );
  AND2X1 \us00/U252  ( .A(\us00/n223 ), .B(\us00/n240 ), .Y(\us00/n28 ) );
  OAI221XL \us00/U251  ( .A0(\us00/n27 ), .A1(\us00/n44 ), .B0(\us00/n4 ), 
        .B1(\us00/n48 ), .C0(\us00/n311 ), .Y(\us00/n310 ) );
  AOI22X1 \us00/U250  ( .A0(\us00/n89 ), .A1(\us00/n309 ), .B0(\us00/n55 ), 
        .B1(\us00/n310 ), .Y(\us00/n308 ) );
  OAI221XL \us00/U249  ( .A0(\us00/n306 ), .A1(\us00/n52 ), .B0(\us00/n307 ), 
        .B1(\us00/n114 ), .C0(\us00/n308 ), .Y(\us00/n305 ) );
  MX2X1 \us00/U248  ( .A(\us00/n304 ), .B(\us00/n305 ), .S0(sa00[6]), .Y(
        sa00_sr[1]) );
  INVX1 \us00/U247  ( .A(\us00/n187 ), .Y(\us00/n61 ) );
  MXI2X1 \us00/U246  ( .A(\us00/n303 ), .B(\us00/n61 ), .S0(\us00/n69 ), .Y(
        \us00/n301 ) );
  MXI2X1 \us00/U245  ( .A(\us00/n301 ), .B(\us00/n147 ), .S0(\us00/n302 ), .Y(
        \us00/n285 ) );
  NAND2X1 \us00/U244  ( .A(\us00/n200 ), .B(\us00/n300 ), .Y(\us00/n99 ) );
  INVX1 \us00/U243  ( .A(\us00/n99 ), .Y(\us00/n296 ) );
  NOR2X1 \us00/U242  ( .A(\us00/n299 ), .B(\us00/n242 ), .Y(\us00/n298 ) );
  NAND2X1 \us00/U241  ( .A(sa00[1]), .B(\us00/n47 ), .Y(\us00/n122 ) );
  NOR2X1 \us00/U240  ( .A(\us00/n159 ), .B(\us00/n217 ), .Y(\us00/n198 ) );
  OAI221XL \us00/U239  ( .A0(\us00/n298 ), .A1(\us00/n27 ), .B0(\us00/n20 ), 
        .B1(\us00/n122 ), .C0(\us00/n132 ), .Y(\us00/n297 ) );
  AOI221X1 \us00/U238  ( .A0(\us00/n225 ), .A1(\us00/n226 ), .B0(\us00/n296 ), 
        .B1(\us00/n6 ), .C0(\us00/n297 ), .Y(\us00/n291 ) );
  OAI2BB2X1 \us00/U237  ( .B0(\us00/n27 ), .B1(\us00/n295 ), .A0N(\us00/n34 ), 
        .A1N(\us00/n24 ), .Y(\us00/n293 ) );
  AOI21X1 \us00/U236  ( .A0(\us00/n101 ), .A1(\us00/n150 ), .B0(\us00/n20 ), 
        .Y(\us00/n294 ) );
  AOI211X1 \us00/U235  ( .A0(\us00/n5 ), .A1(\us00/n79 ), .B0(\us00/n293 ), 
        .C0(\us00/n294 ), .Y(\us00/n292 ) );
  INVX1 \us00/U234  ( .A(\us00/n89 ), .Y(\us00/n10 ) );
  OAI22X1 \us00/U233  ( .A0(\us00/n291 ), .A1(\us00/n114 ), .B0(\us00/n292 ), 
        .B1(\us00/n10 ), .Y(\us00/n286 ) );
  INVX1 \us00/U232  ( .A(\us00/n225 ), .Y(\us00/n288 ) );
  NAND2X1 \us00/U231  ( .A(\us00/n200 ), .B(\us00/n284 ), .Y(\us00/n102 ) );
  NOR2X1 \us00/U230  ( .A(\us00/n290 ), .B(\us00/n163 ), .Y(\us00/n184 ) );
  AOI22X1 \us00/U229  ( .A0(\us00/n102 ), .A1(\us00/n69 ), .B0(\us00/n184 ), 
        .B1(\us00/n33 ), .Y(\us00/n289 ) );
  AOI31X1 \us00/U228  ( .A0(\us00/n132 ), .A1(\us00/n288 ), .A2(\us00/n289 ), 
        .B0(\us00/n52 ), .Y(\us00/n287 ) );
  AOI211X1 \us00/U227  ( .A0(\us00/n285 ), .A1(\us00/n55 ), .B0(\us00/n286 ), 
        .C0(\us00/n287 ), .Y(\us00/n263 ) );
  NAND2X1 \us00/U226  ( .A(\us00/n284 ), .B(\us00/n122 ), .Y(\us00/n125 ) );
  NOR2X1 \us00/U225  ( .A(\us00/n199 ), .B(\us00/n4 ), .Y(\us00/n50 ) );
  AOI21X1 \us00/U224  ( .A0(\us00/n200 ), .A1(\us00/n223 ), .B0(\us00/n20 ), 
        .Y(\us00/n283 ) );
  AOI211X1 \us00/U223  ( .A0(\us00/n5 ), .A1(\us00/n125 ), .B0(\us00/n50 ), 
        .C0(\us00/n283 ), .Y(\us00/n282 ) );
  OAI221XL \us00/U222  ( .A0(\us00/n281 ), .A1(\us00/n27 ), .B0(\us00/n4 ), 
        .B1(\us00/n111 ), .C0(\us00/n282 ), .Y(\us00/n265 ) );
  INVX1 \us00/U221  ( .A(\us00/n280 ), .Y(\us00/n247 ) );
  NAND2X1 \us00/U220  ( .A(\us00/n41 ), .B(\us00/n33 ), .Y(\us00/n272 ) );
  OAI221XL \us00/U219  ( .A0(sa00[1]), .A1(\us00/n247 ), .B0(\us00/n4 ), .B1(
        \us00/n189 ), .C0(\us00/n272 ), .Y(\us00/n279 ) );
  NAND2X1 \us00/U218  ( .A(sa00[2]), .B(\us00/n149 ), .Y(\us00/n276 ) );
  XNOR2X1 \us00/U217  ( .A(\us00/n129 ), .B(sa00[1]), .Y(\us00/n155 ) );
  MXI2X1 \us00/U216  ( .A(\us00/n276 ), .B(\us00/n277 ), .S0(\us00/n155 ), .Y(
        \us00/n275 ) );
  OAI22X1 \us00/U215  ( .A0(\us00/n273 ), .A1(\us00/n10 ), .B0(\us00/n274 ), 
        .B1(\us00/n52 ), .Y(\us00/n266 ) );
  NOR2X1 \us00/U214  ( .A(\us00/n20 ), .B(\us00/n226 ), .Y(\us00/n176 ) );
  OAI21XL \us00/U213  ( .A0(\us00/n4 ), .A1(\us00/n271 ), .B0(\us00/n272 ), 
        .Y(\us00/n270 ) );
  OAI31X1 \us00/U212  ( .A0(\us00/n176 ), .A1(\us00/n269 ), .A2(\us00/n270 ), 
        .B0(\us00/n16 ), .Y(\us00/n268 ) );
  INVX1 \us00/U211  ( .A(\us00/n268 ), .Y(\us00/n267 ) );
  AOI211X1 \us00/U210  ( .A0(\us00/n55 ), .A1(\us00/n265 ), .B0(\us00/n266 ), 
        .C0(\us00/n267 ), .Y(\us00/n264 ) );
  MXI2X1 \us00/U209  ( .A(\us00/n263 ), .B(\us00/n264 ), .S0(sa00[6]), .Y(
        sa00_sr[2]) );
  NOR2X1 \us00/U208  ( .A(\us00/n94 ), .B(sa00[1]), .Y(\us00/n211 ) );
  INVX1 \us00/U207  ( .A(\us00/n262 ), .Y(\us00/n261 ) );
  AOI211X1 \us00/U206  ( .A0(\us00/n259 ), .A1(\us00/n24 ), .B0(\us00/n260 ), 
        .C0(\us00/n261 ), .Y(\us00/n255 ) );
  OAI22X1 \us00/U205  ( .A0(\us00/n20 ), .A1(\us00/n68 ), .B0(\us00/n27 ), 
        .B1(\us00/n37 ), .Y(\us00/n257 ) );
  NOR3X1 \us00/U204  ( .A(\us00/n257 ), .B(\us00/n258 ), .C(\us00/n50 ), .Y(
        \us00/n256 ) );
  MXI2X1 \us00/U203  ( .A(\us00/n255 ), .B(\us00/n256 ), .S0(\us00/n252 ), .Y(
        \us00/n254 ) );
  AOI221X1 \us00/U202  ( .A0(\us00/n211 ), .A1(\us00/n5 ), .B0(\us00/n40 ), 
        .B1(sa00[4]), .C0(\us00/n254 ), .Y(\us00/n248 ) );
  INVX1 \us00/U201  ( .A(\us00/n211 ), .Y(\us00/n106 ) );
  NAND2X1 \us00/U200  ( .A(\us00/n200 ), .B(\us00/n106 ), .Y(\us00/n83 ) );
  NAND2X1 \us00/U199  ( .A(\us00/n199 ), .B(\us00/n204 ), .Y(\us00/n169 ) );
  AOI2BB2X1 \us00/U198  ( .B0(\us00/n65 ), .B1(\us00/n24 ), .A0N(\us00/n169 ), 
        .A1N(\us00/n20 ), .Y(\us00/n253 ) );
  OAI221XL \us00/U197  ( .A0(\us00/n172 ), .A1(\us00/n18 ), .B0(\us00/n27 ), 
        .B1(\us00/n83 ), .C0(\us00/n253 ), .Y(\us00/n251 ) );
  MXI2X1 \us00/U196  ( .A(\us00/n250 ), .B(\us00/n251 ), .S0(\us00/n252 ), .Y(
        \us00/n249 ) );
  MXI2X1 \us00/U195  ( .A(\us00/n248 ), .B(\us00/n249 ), .S0(\us00/n234 ), .Y(
        \us00/n228 ) );
  OAI21XL \us00/U194  ( .A0(\us00/n58 ), .A1(\us00/n27 ), .B0(\us00/n247 ), 
        .Y(\us00/n245 ) );
  NOR2X1 \us00/U193  ( .A(sa00[7]), .B(\us00/n145 ), .Y(\us00/n246 ) );
  XNOR2X1 \us00/U192  ( .A(\us00/n69 ), .B(sa00[1]), .Y(\us00/n130 ) );
  MXI2X1 \us00/U191  ( .A(\us00/n245 ), .B(\us00/n246 ), .S0(\us00/n130 ), .Y(
        \us00/n243 ) );
  OAI211X1 \us00/U190  ( .A0(\us00/n4 ), .A1(\us00/n149 ), .B0(\us00/n243 ), 
        .C0(\us00/n244 ), .Y(\us00/n230 ) );
  NOR2X1 \us00/U189  ( .A(\us00/n242 ), .B(\us00/n137 ), .Y(\us00/n70 ) );
  OAI221XL \us00/U188  ( .A0(\us00/n159 ), .A1(\us00/n27 ), .B0(\us00/n20 ), 
        .B1(\us00/n34 ), .C0(\us00/n241 ), .Y(\us00/n231 ) );
  NAND2X1 \us00/U187  ( .A(\us00/n101 ), .B(\us00/n240 ), .Y(\us00/n76 ) );
  AOI21X1 \us00/U186  ( .A0(\us00/n122 ), .A1(\us00/n106 ), .B0(\us00/n129 ), 
        .Y(\us00/n237 ) );
  INVX1 \us00/U185  ( .A(\us00/n239 ), .Y(\us00/n238 ) );
  OAI21XL \us00/U184  ( .A0(\us00/n237 ), .A1(\us00/n43 ), .B0(\us00/n238 ), 
        .Y(\us00/n236 ) );
  OAI221XL \us00/U183  ( .A0(\us00/n18 ), .A1(\us00/n76 ), .B0(\us00/n59 ), 
        .B1(\us00/n27 ), .C0(\us00/n236 ), .Y(\us00/n232 ) );
  AOI2BB2X1 \us00/U182  ( .B0(\us00/n24 ), .B1(\us00/n187 ), .A0N(\us00/n227 ), 
        .A1N(\us00/n20 ), .Y(\us00/n235 ) );
  OAI211X1 \us00/U181  ( .A0(\us00/n27 ), .A1(\us00/n122 ), .B0(\us00/n158 ), 
        .C0(\us00/n235 ), .Y(\us00/n233 ) );
  MX4X1 \us00/U180  ( .A(\us00/n230 ), .B(\us00/n231 ), .C(\us00/n232 ), .D(
        \us00/n233 ), .S0(\us00/n234 ), .S1(sa00[5]), .Y(\us00/n229 ) );
  MX2X1 \us00/U179  ( .A(\us00/n228 ), .B(\us00/n229 ), .S0(sa00[6]), .Y(
        sa00_sr[3]) );
  NOR2BX1 \us00/U178  ( .AN(\us00/n204 ), .B(\us00/n137 ), .Y(\us00/n110 ) );
  INVX1 \us00/U177  ( .A(\us00/n110 ), .Y(\us00/n64 ) );
  AOI22X1 \us00/U176  ( .A0(\us00/n225 ), .A1(\us00/n226 ), .B0(\us00/n6 ), 
        .B1(\us00/n227 ), .Y(\us00/n224 ) );
  OAI221XL \us00/U175  ( .A0(\us00/n27 ), .A1(\us00/n64 ), .B0(\us00/n4 ), 
        .B1(\us00/n83 ), .C0(\us00/n224 ), .Y(\us00/n212 ) );
  NAND2X1 \us00/U174  ( .A(\us00/n34 ), .B(\us00/n204 ), .Y(\us00/n221 ) );
  OAI21XL \us00/U173  ( .A0(\us00/n69 ), .A1(\us00/n223 ), .B0(\us00/n27 ), 
        .Y(\us00/n222 ) );
  NOR2X1 \us00/U172  ( .A(\us00/n217 ), .B(\us00/n42 ), .Y(\us00/n208 ) );
  AOI211X1 \us00/U171  ( .A0(\us00/n208 ), .A1(\us00/n5 ), .B0(\us00/n220 ), 
        .C0(\us00/n173 ), .Y(\us00/n219 ) );
  OAI22X1 \us00/U170  ( .A0(\us00/n218 ), .A1(\us00/n10 ), .B0(\us00/n219 ), 
        .B1(\us00/n114 ), .Y(\us00/n213 ) );
  INVX1 \us00/U169  ( .A(\us00/n135 ), .Y(\us00/n215 ) );
  NOR2X1 \us00/U168  ( .A(\us00/n4 ), .B(\us00/n159 ), .Y(\us00/n31 ) );
  INVX1 \us00/U167  ( .A(\us00/n31 ), .Y(\us00/n196 ) );
  AOI31X1 \us00/U166  ( .A0(\us00/n215 ), .A1(\us00/n196 ), .A2(\us00/n216 ), 
        .B0(\us00/n52 ), .Y(\us00/n214 ) );
  AOI211X1 \us00/U165  ( .A0(\us00/n55 ), .A1(\us00/n212 ), .B0(\us00/n213 ), 
        .C0(\us00/n214 ), .Y(\us00/n190 ) );
  INVX1 \us00/U164  ( .A(\us00/n207 ), .Y(\us00/n192 ) );
  NOR2X1 \us00/U163  ( .A(\us00/n25 ), .B(\us00/n98 ), .Y(\us00/n32 ) );
  OAI22X1 \us00/U162  ( .A0(\us00/n28 ), .A1(\us00/n4 ), .B0(\us00/n188 ), 
        .B1(\us00/n27 ), .Y(\us00/n206 ) );
  NAND2X1 \us00/U161  ( .A(\us00/n204 ), .B(\us00/n80 ), .Y(\us00/n118 ) );
  INVX1 \us00/U160  ( .A(\us00/n118 ), .Y(\us00/n123 ) );
  NAND2X1 \us00/U159  ( .A(\us00/n94 ), .B(\us00/n79 ), .Y(\us00/n203 ) );
  OAI2BB1X1 \us00/U158  ( .A0N(\us00/n199 ), .A1N(\us00/n200 ), .B0(\us00/n33 ), .Y(\us00/n195 ) );
  INVX1 \us00/U157  ( .A(\us00/n55 ), .Y(\us00/n12 ) );
  AOI31X1 \us00/U156  ( .A0(\us00/n195 ), .A1(\us00/n196 ), .A2(\us00/n197 ), 
        .B0(\us00/n12 ), .Y(\us00/n194 ) );
  AOI211X1 \us00/U155  ( .A0(\us00/n89 ), .A1(\us00/n192 ), .B0(\us00/n193 ), 
        .C0(\us00/n194 ), .Y(\us00/n191 ) );
  MXI2X1 \us00/U154  ( .A(\us00/n190 ), .B(\us00/n191 ), .S0(sa00[6]), .Y(
        sa00_sr[4]) );
  OAI21XL \us00/U153  ( .A0(\us00/n69 ), .A1(\us00/n189 ), .B0(\us00/n27 ), 
        .Y(\us00/n186 ) );
  INVX1 \us00/U152  ( .A(\us00/n183 ), .Y(\us00/n180 ) );
  NAND2X1 \us00/U151  ( .A(\us00/n74 ), .B(\us00/n182 ), .Y(\us00/n181 ) );
  AOI211X1 \us00/U150  ( .A0(\us00/n179 ), .A1(\us00/n24 ), .B0(\us00/n180 ), 
        .C0(\us00/n181 ), .Y(\us00/n165 ) );
  INVX1 \us00/U149  ( .A(\us00/n178 ), .Y(\us00/n175 ) );
  AOI211X1 \us00/U148  ( .A0(\us00/n175 ), .A1(\us00/n5 ), .B0(\us00/n176 ), 
        .C0(\us00/n177 ), .Y(\us00/n174 ) );
  OAI221XL \us00/U147  ( .A0(\us00/n159 ), .A1(\us00/n27 ), .B0(\us00/n145 ), 
        .B1(\us00/n20 ), .C0(\us00/n174 ), .Y(\us00/n167 ) );
  MXI2X1 \us00/U146  ( .A(\us00/n40 ), .B(\us00/n173 ), .S0(\us00/n96 ), .Y(
        \us00/n170 ) );
  AOI22X1 \us00/U145  ( .A0(\us00/n137 ), .A1(\us00/n24 ), .B0(\us00/n172 ), 
        .B1(\us00/n6 ), .Y(\us00/n171 ) );
  OAI211X1 \us00/U144  ( .A0(\us00/n20 ), .A1(\us00/n169 ), .B0(\us00/n170 ), 
        .C0(\us00/n171 ), .Y(\us00/n168 ) );
  AOI22X1 \us00/U143  ( .A0(\us00/n89 ), .A1(\us00/n167 ), .B0(\us00/n55 ), 
        .B1(\us00/n168 ), .Y(\us00/n166 ) );
  OAI221XL \us00/U142  ( .A0(\us00/n164 ), .A1(\us00/n114 ), .B0(\us00/n165 ), 
        .B1(\us00/n52 ), .C0(\us00/n166 ), .Y(\us00/n138 ) );
  OAI21XL \us00/U141  ( .A0(\us00/n41 ), .A1(\us00/n163 ), .B0(\us00/n69 ), 
        .Y(\us00/n162 ) );
  AOI221X1 \us00/U140  ( .A0(\us00/n159 ), .A1(\us00/n24 ), .B0(\us00/n160 ), 
        .B1(\us00/n33 ), .C0(\us00/n161 ), .Y(\us00/n140 ) );
  OAI21XL \us00/U139  ( .A0(\us00/n157 ), .A1(\us00/n20 ), .B0(\us00/n158 ), 
        .Y(\us00/n156 ) );
  NOR2X1 \us00/U138  ( .A(\us00/n4 ), .B(\us00/n136 ), .Y(\us00/n153 ) );
  NOR2X1 \us00/U137  ( .A(\us00/n145 ), .B(\us00/n69 ), .Y(\us00/n154 ) );
  MXI2X1 \us00/U136  ( .A(\us00/n153 ), .B(\us00/n154 ), .S0(\us00/n155 ), .Y(
        \us00/n152 ) );
  OAI221XL \us00/U135  ( .A0(\us00/n110 ), .A1(\us00/n18 ), .B0(\us00/n20 ), 
        .B1(\us00/n151 ), .C0(\us00/n152 ), .Y(\us00/n143 ) );
  AOI21X1 \us00/U134  ( .A0(\us00/n149 ), .A1(\us00/n150 ), .B0(\us00/n18 ), 
        .Y(\us00/n148 ) );
  AOI2BB1X1 \us00/U133  ( .A0N(\us00/n147 ), .A1N(\us00/n27 ), .B0(\us00/n148 ), .Y(\us00/n146 ) );
  OAI221XL \us00/U132  ( .A0(\us00/n145 ), .A1(\us00/n20 ), .B0(\us00/n4 ), 
        .B1(\us00/n34 ), .C0(\us00/n146 ), .Y(\us00/n144 ) );
  AOI22X1 \us00/U131  ( .A0(\us00/n89 ), .A1(\us00/n143 ), .B0(\us00/n14 ), 
        .B1(\us00/n144 ), .Y(\us00/n142 ) );
  OAI221XL \us00/U130  ( .A0(\us00/n140 ), .A1(\us00/n12 ), .B0(\us00/n141 ), 
        .B1(\us00/n114 ), .C0(\us00/n142 ), .Y(\us00/n139 ) );
  MX2X1 \us00/U129  ( .A(\us00/n138 ), .B(\us00/n139 ), .S0(sa00[6]), .Y(
        sa00_sr[5]) );
  INVX1 \us00/U128  ( .A(\us00/n70 ), .Y(\us00/n133 ) );
  OAI22X1 \us00/U127  ( .A0(\us00/n4 ), .A1(\us00/n136 ), .B0(\us00/n137 ), 
        .B1(\us00/n27 ), .Y(\us00/n134 ) );
  AOI211X1 \us00/U126  ( .A0(\us00/n133 ), .A1(\us00/n69 ), .B0(\us00/n134 ), 
        .C0(\us00/n135 ), .Y(\us00/n112 ) );
  INVX1 \us00/U125  ( .A(\us00/n132 ), .Y(\us00/n131 ) );
  OAI21XL \us00/U124  ( .A0(\us00/n18 ), .A1(\us00/n37 ), .B0(\us00/n128 ), 
        .Y(\us00/n127 ) );
  OAI221XL \us00/U123  ( .A0(\us00/n18 ), .A1(\us00/n105 ), .B0(\us00/n123 ), 
        .B1(\us00/n27 ), .C0(\us00/n124 ), .Y(\us00/n116 ) );
  NAND2X1 \us00/U122  ( .A(\us00/n121 ), .B(\us00/n122 ), .Y(\us00/n30 ) );
  OAI221XL \us00/U121  ( .A0(\us00/n18 ), .A1(\us00/n118 ), .B0(\us00/n27 ), 
        .B1(\us00/n30 ), .C0(\us00/n119 ), .Y(\us00/n117 ) );
  AOI22X1 \us00/U120  ( .A0(\us00/n89 ), .A1(\us00/n116 ), .B0(\us00/n55 ), 
        .B1(\us00/n117 ), .Y(\us00/n115 ) );
  OAI221XL \us00/U119  ( .A0(\us00/n112 ), .A1(\us00/n52 ), .B0(\us00/n113 ), 
        .B1(\us00/n114 ), .C0(\us00/n115 ), .Y(\us00/n84 ) );
  OAI22X1 \us00/U118  ( .A0(\us00/n110 ), .A1(\us00/n4 ), .B0(\us00/n20 ), 
        .B1(\us00/n21 ), .Y(\us00/n108 ) );
  AOI21X1 \us00/U117  ( .A0(sa00[1]), .A1(\us00/n58 ), .B0(\us00/n27 ), .Y(
        \us00/n109 ) );
  AOI211X1 \us00/U116  ( .A0(\us00/n5 ), .A1(\us00/n107 ), .B0(\us00/n108 ), 
        .C0(\us00/n109 ), .Y(\us00/n86 ) );
  OAI22X1 \us00/U115  ( .A0(\us00/n45 ), .A1(\us00/n4 ), .B0(sa00[4]), .B1(
        \us00/n18 ), .Y(\us00/n103 ) );
  AOI21X1 \us00/U114  ( .A0(\us00/n105 ), .A1(\us00/n106 ), .B0(\us00/n20 ), 
        .Y(\us00/n104 ) );
  AOI211X1 \us00/U113  ( .A0(\us00/n33 ), .A1(\us00/n102 ), .B0(\us00/n103 ), 
        .C0(\us00/n104 ), .Y(\us00/n87 ) );
  NAND2X1 \us00/U112  ( .A(\us00/n100 ), .B(\us00/n101 ), .Y(\us00/n62 ) );
  OAI221XL \us00/U111  ( .A0(\us00/n27 ), .A1(\us00/n62 ), .B0(\us00/n4 ), 
        .B1(\us00/n21 ), .C0(\us00/n97 ), .Y(\us00/n90 ) );
  NOR3X1 \us00/U110  ( .A(\us00/n4 ), .B(\us00/n95 ), .C(\us00/n96 ), .Y(
        \us00/n67 ) );
  AOI31X1 \us00/U109  ( .A0(\us00/n79 ), .A1(\us00/n94 ), .A2(\us00/n6 ), .B0(
        \us00/n67 ), .Y(\us00/n93 ) );
  OAI221XL \us00/U108  ( .A0(\us00/n73 ), .A1(\us00/n27 ), .B0(\us00/n92 ), 
        .B1(\us00/n20 ), .C0(\us00/n93 ), .Y(\us00/n91 ) );
  AOI22X1 \us00/U107  ( .A0(\us00/n89 ), .A1(\us00/n90 ), .B0(\us00/n16 ), 
        .B1(\us00/n91 ), .Y(\us00/n88 ) );
  OAI221XL \us00/U106  ( .A0(\us00/n86 ), .A1(\us00/n52 ), .B0(\us00/n87 ), 
        .B1(\us00/n12 ), .C0(\us00/n88 ), .Y(\us00/n85 ) );
  MX2X1 \us00/U105  ( .A(\us00/n84 ), .B(\us00/n85 ), .S0(sa00[6]), .Y(
        sa00_sr[6]) );
  INVX1 \us00/U104  ( .A(\us00/n81 ), .Y(\us00/n77 ) );
  AOI21X1 \us00/U103  ( .A0(\us00/n79 ), .A1(\us00/n80 ), .B0(\us00/n27 ), .Y(
        \us00/n78 ) );
  AOI211X1 \us00/U102  ( .A0(\us00/n5 ), .A1(\us00/n76 ), .B0(\us00/n77 ), 
        .C0(\us00/n78 ), .Y(\us00/n51 ) );
  OAI211X1 \us00/U101  ( .A0(\us00/n73 ), .A1(\us00/n27 ), .B0(\us00/n74 ), 
        .C0(\us00/n75 ), .Y(\us00/n72 ) );
  AOI21X1 \us00/U100  ( .A0(\us00/n68 ), .A1(\us00/n69 ), .B0(\us00/n6 ), .Y(
        \us00/n63 ) );
  INVX1 \us00/U99  ( .A(\us00/n67 ), .Y(\us00/n66 ) );
  OAI221XL \us00/U98  ( .A0(\us00/n63 ), .A1(\us00/n64 ), .B0(\us00/n65 ), 
        .B1(\us00/n27 ), .C0(\us00/n66 ), .Y(\us00/n56 ) );
  AOI2BB2X1 \us00/U97  ( .B0(\us00/n61 ), .B1(\us00/n24 ), .A0N(\us00/n62 ), 
        .A1N(\us00/n20 ), .Y(\us00/n60 ) );
  OAI221XL \us00/U96  ( .A0(\us00/n58 ), .A1(\us00/n18 ), .B0(\us00/n59 ), 
        .B1(\us00/n27 ), .C0(\us00/n60 ), .Y(\us00/n57 ) );
  AOI22X1 \us00/U95  ( .A0(\us00/n55 ), .A1(\us00/n56 ), .B0(\us00/n16 ), .B1(
        \us00/n57 ), .Y(\us00/n54 ) );
  OAI221XL \us00/U94  ( .A0(\us00/n51 ), .A1(\us00/n52 ), .B0(\us00/n53 ), 
        .B1(\us00/n10 ), .C0(\us00/n54 ), .Y(\us00/n7 ) );
  INVX1 \us00/U93  ( .A(\us00/n50 ), .Y(\us00/n49 ) );
  OAI221XL \us00/U92  ( .A0(\us00/n47 ), .A1(\us00/n18 ), .B0(\us00/n27 ), 
        .B1(\us00/n48 ), .C0(\us00/n49 ), .Y(\us00/n46 ) );
  NOR2X1 \us00/U91  ( .A(\us00/n41 ), .B(\us00/n42 ), .Y(\us00/n38 ) );
  INVX1 \us00/U90  ( .A(\us00/n40 ), .Y(\us00/n39 ) );
  INVX1 \us00/U89  ( .A(\us00/n32 ), .Y(\us00/n26 ) );
  AOI21X1 \us00/U88  ( .A0(\us00/n5 ), .A1(\us00/n30 ), .B0(\us00/n31 ), .Y(
        \us00/n29 ) );
  OAI221XL \us00/U87  ( .A0(\us00/n26 ), .A1(\us00/n27 ), .B0(\us00/n28 ), 
        .B1(\us00/n20 ), .C0(\us00/n29 ), .Y(\us00/n15 ) );
  OAI221XL \us00/U86  ( .A0(\us00/n18 ), .A1(\us00/n19 ), .B0(\us00/n20 ), 
        .B1(\us00/n21 ), .C0(\us00/n22 ), .Y(\us00/n17 ) );
  AOI22X1 \us00/U85  ( .A0(\us00/n14 ), .A1(\us00/n15 ), .B0(\us00/n16 ), .B1(
        \us00/n17 ), .Y(\us00/n13 ) );
  OAI221XL \us00/U84  ( .A0(\us00/n9 ), .A1(\us00/n10 ), .B0(\us00/n11 ), .B1(
        \us00/n12 ), .C0(\us00/n13 ), .Y(\us00/n8 ) );
  MX2X1 \us00/U83  ( .A(\us00/n7 ), .B(\us00/n8 ), .S0(sa00[6]), .Y(sa00_sr[7]) );
  NOR2X4 \us00/U82  ( .A(\us00/n129 ), .B(sa00[2]), .Y(\us00/n43 ) );
  CLKINVX3 \us00/U81  ( .A(\us00/n14 ), .Y(\us00/n52 ) );
  OAI22XL \us00/U80  ( .A0(\us00/n201 ), .A1(\us00/n52 ), .B0(\us00/n202 ), 
        .B1(\us00/n114 ), .Y(\us00/n193 ) );
  CLKINVX3 \us00/U79  ( .A(sa00[5]), .Y(\us00/n252 ) );
  NOR2X2 \us00/U78  ( .A(\us00/n252 ), .B(\us00/n234 ), .Y(\us00/n55 ) );
  CLKINVX3 \us00/U77  ( .A(sa00[7]), .Y(\us00/n129 ) );
  NOR2X4 \us00/U76  ( .A(\us00/n129 ), .B(\us00/n69 ), .Y(\us00/n24 ) );
  AOI22XL \us00/U75  ( .A0(\us00/n70 ), .A1(\us00/n24 ), .B0(\us00/n96 ), .B1(
        \us00/n129 ), .Y(\us00/n241 ) );
  NOR2X2 \us00/U74  ( .A(\us00/n252 ), .B(sa00[0]), .Y(\us00/n89 ) );
  CLKINVX3 \us00/U73  ( .A(sa00[0]), .Y(\us00/n234 ) );
  NOR2X4 \us00/U72  ( .A(\us00/n69 ), .B(sa00[7]), .Y(\us00/n33 ) );
  INVX12 \us00/U71  ( .A(\us00/n33 ), .Y(\us00/n27 ) );
  CLKINVX3 \us00/U70  ( .A(\us00/n1 ), .Y(\us00/n6 ) );
  CLKINVX3 \us00/U69  ( .A(\us00/n1 ), .Y(\us00/n5 ) );
  INVXL \us00/U68  ( .A(\us00/n24 ), .Y(\us00/n36 ) );
  INVX4 \us00/U67  ( .A(\us00/n3 ), .Y(\us00/n4 ) );
  INVXL \us00/U66  ( .A(\us00/n36 ), .Y(\us00/n3 ) );
  INVX4 \us00/U65  ( .A(sa00[1]), .Y(\us00/n226 ) );
  INVX4 \us00/U64  ( .A(\us00/n43 ), .Y(\us00/n20 ) );
  AOI221X4 \us00/U63  ( .A0(\us00/n24 ), .A1(\us00/n82 ), .B0(\us00/n43 ), 
        .B1(\us00/n295 ), .C0(\us00/n173 ), .Y(\us00/n346 ) );
  AOI221X4 \us00/U62  ( .A0(\us00/n5 ), .A1(\us00/n96 ), .B0(\us00/n43 ), .B1(
        \us00/n239 ), .C0(\us00/n340 ), .Y(\us00/n336 ) );
  AOI222X4 \us00/U61  ( .A0(\us00/n59 ), .A1(\us00/n43 ), .B0(\us00/n6 ), .B1(
        \us00/n221 ), .C0(\us00/n222 ), .C1(\us00/n187 ), .Y(\us00/n218 ) );
  AOI222X4 \us00/U60  ( .A0(\us00/n123 ), .A1(\us00/n43 ), .B0(sa00[2]), .B1(
        \us00/n203 ), .C0(\us00/n6 ), .C1(\us00/n71 ), .Y(\us00/n202 ) );
  AOI221X4 \us00/U59  ( .A0(\us00/n314 ), .A1(\us00/n43 ), .B0(\us00/n160 ), 
        .B1(\us00/n24 ), .C0(\us00/n315 ), .Y(\us00/n307 ) );
  AOI221X4 \us00/U58  ( .A0(\us00/n43 ), .A1(\us00/n208 ), .B0(\us00/n76 ), 
        .B1(\us00/n24 ), .C0(\us00/n209 ), .Y(\us00/n207 ) );
  AOI221X4 \us00/U57  ( .A0(\us00/n43 ), .A1(\us00/n205 ), .B0(\us00/n32 ), 
        .B1(\us00/n6 ), .C0(\us00/n206 ), .Y(\us00/n201 ) );
  AOI221X4 \us00/U56  ( .A0(\us00/n43 ), .A1(\us00/n44 ), .B0(\us00/n45 ), 
        .B1(\us00/n24 ), .C0(\us00/n46 ), .Y(\us00/n9 ) );
  AOI22XL \us00/U55  ( .A0(\us00/n217 ), .A1(\us00/n43 ), .B0(\us00/n33 ), 
        .B1(\us00/n47 ), .Y(\us00/n216 ) );
  AOI22XL \us00/U54  ( .A0(\us00/n98 ), .A1(\us00/n43 ), .B0(\us00/n6 ), .B1(
        \us00/n99 ), .Y(\us00/n97 ) );
  AOI22XL \us00/U53  ( .A0(\us00/n82 ), .A1(\us00/n43 ), .B0(\us00/n83 ), .B1(
        \us00/n24 ), .Y(\us00/n81 ) );
  AOI2BB2XL \us00/U52  ( .B0(\us00/n43 ), .B1(\us00/n94 ), .A0N(\us00/n120 ), 
        .A1N(\us00/n4 ), .Y(\us00/n119 ) );
  AOI222X4 \us00/U51  ( .A0(\us00/n125 ), .A1(\us00/n33 ), .B0(\us00/n145 ), 
        .B1(\us00/n40 ), .C0(\us00/n43 ), .C1(\us00/n184 ), .Y(\us00/n183 ) );
  AOI22XL \us00/U50  ( .A0(\us00/n43 ), .A1(\us00/n303 ), .B0(\us00/n24 ), 
        .B1(\us00/n96 ), .Y(\us00/n358 ) );
  AOI22XL \us00/U49  ( .A0(\us00/n43 ), .A1(\us00/n100 ), .B0(\us00/n24 ), 
        .B1(\us00/n125 ), .Y(\us00/n124 ) );
  AOI21XL \us00/U48  ( .A0(\us00/n159 ), .A1(\us00/n43 ), .B0(\us00/n40 ), .Y(
        \us00/n262 ) );
  AOI22XL \us00/U47  ( .A0(\us00/n40 ), .A1(\us00/n94 ), .B0(\us00/n43 ), .B1(
        \us00/n187 ), .Y(\us00/n244 ) );
  AOI22XL \us00/U46  ( .A0(\us00/n184 ), .A1(\us00/n5 ), .B0(\us00/n198 ), 
        .B1(\us00/n43 ), .Y(\us00/n197 ) );
  NOR2XL \us00/U45  ( .A(\us00/n33 ), .B(\us00/n2 ), .Y(\us00/n302 ) );
  MXI2XL \us00/U44  ( .A(\us00/n2 ), .B(\us00/n6 ), .S0(\us00/n28 ), .Y(
        \us00/n311 ) );
  INVXL \us00/U43  ( .A(\us00/n20 ), .Y(\us00/n2 ) );
  INVX4 \us00/U42  ( .A(\us00/n6 ), .Y(\us00/n18 ) );
  AOI21XL \us00/U41  ( .A0(\us00/n18 ), .A1(\us00/n162 ), .B0(\us00/n25 ), .Y(
        \us00/n161 ) );
  INVX4 \us00/U40  ( .A(sa00[2]), .Y(\us00/n69 ) );
  NOR2X4 \us00/U39  ( .A(\us00/n226 ), .B(\us00/n4 ), .Y(\us00/n40 ) );
  CLKINVX3 \us00/U38  ( .A(sa00[3]), .Y(\us00/n136 ) );
  NOR2X2 \us00/U37  ( .A(\us00/n136 ), .B(sa00[4]), .Y(\us00/n145 ) );
  CLKINVX3 \us00/U36  ( .A(sa00[4]), .Y(\us00/n58 ) );
  NOR2X2 \us00/U35  ( .A(\us00/n58 ), .B(sa00[3]), .Y(\us00/n159 ) );
  NOR2X2 \us00/U34  ( .A(\us00/n136 ), .B(\us00/n58 ), .Y(\us00/n259 ) );
  NOR2X2 \us00/U33  ( .A(sa00[4]), .B(sa00[3]), .Y(\us00/n278 ) );
  NOR2X2 \us00/U32  ( .A(\us00/n259 ), .B(\us00/n278 ), .Y(\us00/n47 ) );
  CLKINVX3 \us00/U31  ( .A(\us00/n259 ), .Y(\us00/n44 ) );
  NOR2X2 \us00/U30  ( .A(\us00/n44 ), .B(sa00[1]), .Y(\us00/n137 ) );
  AOI21XL \us00/U29  ( .A0(\us00/n44 ), .A1(\us00/n111 ), .B0(\us00/n4 ), .Y(
        \us00/n177 ) );
  AOI22XL \us00/U28  ( .A0(\us00/n23 ), .A1(\us00/n24 ), .B0(\us00/n25 ), .B1(
        sa00[2]), .Y(\us00/n22 ) );
  AOI22XL \us00/U27  ( .A0(\us00/n33 ), .A1(sa00[3]), .B0(\us00/n24 ), .B1(
        \us00/n58 ), .Y(\us00/n277 ) );
  NAND2XL \us00/U26  ( .A(\us00/n198 ), .B(\us00/n24 ), .Y(\us00/n132 ) );
  OAI2BB2XL \us00/U25  ( .B0(\us00/n20 ), .B1(\us00/n111 ), .A0N(\us00/n125 ), 
        .A1N(\us00/n24 ), .Y(\us00/n220 ) );
  NAND2XL \us00/U24  ( .A(\us00/n111 ), .B(\us00/n101 ), .Y(\us00/n21 ) );
  NAND2XL \us00/U23  ( .A(\us00/n111 ), .B(\us00/n300 ), .Y(\us00/n187 ) );
  NAND2XL \us00/U22  ( .A(\us00/n111 ), .B(\us00/n121 ), .Y(\us00/n303 ) );
  AOI221XL \us00/U21  ( .A0(\us00/n43 ), .A1(\us00/n151 ), .B0(\us00/n25 ), 
        .B1(\us00/n69 ), .C0(\us00/n275 ), .Y(\us00/n274 ) );
  NOR2BXL \us00/U20  ( .AN(\us00/n101 ), .B(\us00/n25 ), .Y(\us00/n172 ) );
  NAND2X2 \us00/U19  ( .A(\us00/n58 ), .B(\us00/n226 ), .Y(\us00/n34 ) );
  OAI222X1 \us00/U18  ( .A0(\us00/n27 ), .A1(\us00/n34 ), .B0(\us00/n69 ), 
        .B1(\us00/n205 ), .C0(\us00/n20 ), .C1(\us00/n79 ), .Y(\us00/n260 ) );
  OAI222X1 \us00/U17  ( .A0(\us00/n20 ), .A1(\us00/n99 ), .B0(\us00/n27 ), 
        .B1(\us00/n101 ), .C0(\us00/n184 ), .C1(\us00/n4 ), .Y(\us00/n250 ) );
  OAI222X1 \us00/U16  ( .A0(\us00/n4 ), .A1(\us00/n37 ), .B0(\us00/n38 ), .B1(
        \us00/n20 ), .C0(sa00[4]), .C1(\us00/n39 ), .Y(\us00/n35 ) );
  AOI221X1 \us00/U15  ( .A0(\us00/n5 ), .A1(\us00/n19 ), .B0(\us00/n33 ), .B1(
        \us00/n34 ), .C0(\us00/n35 ), .Y(\us00/n11 ) );
  OR2X2 \us00/U14  ( .A(sa00[2]), .B(sa00[7]), .Y(\us00/n1 ) );
  AOI221XL \us00/U13  ( .A0(\us00/n70 ), .A1(\us00/n43 ), .B0(\us00/n24 ), 
        .B1(\us00/n71 ), .C0(\us00/n72 ), .Y(\us00/n53 ) );
  AOI221XL \us00/U12  ( .A0(\us00/n59 ), .A1(\us00/n33 ), .B0(\us00/n43 ), 
        .B1(\us00/n126 ), .C0(\us00/n127 ), .Y(\us00/n113 ) );
  AOI222XL \us00/U11  ( .A0(\us00/n185 ), .A1(\us00/n43 ), .B0(\us00/n186 ), 
        .B1(\us00/n187 ), .C0(\us00/n6 ), .C1(\us00/n188 ), .Y(\us00/n164 ) );
  AOI221X1 \us00/U10  ( .A0(\us00/n313 ), .A1(\us00/n5 ), .B0(\us00/n23 ), 
        .B1(\us00/n2 ), .C0(\us00/n328 ), .Y(\us00/n320 ) );
  AOI221X1 \us00/U9  ( .A0(\us00/n40 ), .A1(\us00/n136 ), .B0(\us00/n33 ), 
        .B1(\us00/n178 ), .C0(\us00/n338 ), .Y(\us00/n337 ) );
  AOI222XL \us00/U8  ( .A0(\us00/n278 ), .A1(\us00/n24 ), .B0(\us00/n42 ), 
        .B1(\us00/n33 ), .C0(\us00/n43 ), .C1(\us00/n136 ), .Y(\us00/n351 ) );
  AOI31X1 \us00/U7  ( .A0(sa00[2]), .A1(\us00/n58 ), .A2(sa00[1]), .B0(
        \us00/n40 ), .Y(\us00/n350 ) );
  AOI31X1 \us00/U6  ( .A0(\us00/n44 ), .A1(\us00/n129 ), .A2(\us00/n130 ), 
        .B0(\us00/n131 ), .Y(\us00/n128 ) );
  AOI221X1 \us00/U5  ( .A0(\us00/n40 ), .A1(\us00/n136 ), .B0(\us00/n33 ), 
        .B1(\us00/n47 ), .C0(\us00/n156 ), .Y(\us00/n141 ) );
  OAI32X1 \us00/U4  ( .A0(\us00/n210 ), .A1(\us00/n145 ), .A2(\us00/n18 ), 
        .B0(\us00/n27 ), .B1(\us00/n211 ), .Y(\us00/n209 ) );
  AOI221X1 \us00/U3  ( .A0(\us00/n278 ), .A1(\us00/n40 ), .B0(\us00/n185 ), 
        .B1(\us00/n2 ), .C0(\us00/n279 ), .Y(\us00/n273 ) );
  OAI32X1 \us00/U2  ( .A0(\us00/n18 ), .A1(sa00[1]), .A2(\us00/n159 ), .B0(
        sa00[4]), .B1(\us00/n182 ), .Y(\us00/n318 ) );
  AOI31XL \us00/U1  ( .A0(\us00/n79 ), .A1(\us00/n44 ), .A2(\us00/n2 ), .B0(
        \us00/n280 ), .Y(\us00/n339 ) );
  NAND2X1 \us01/U366  ( .A(\us01/n47 ), .B(\us01/n226 ), .Y(\us01/n189 ) );
  NOR2X1 \us01/U365  ( .A(\us01/n226 ), .B(sa01[3]), .Y(\us01/n242 ) );
  INVX1 \us01/U364  ( .A(\us01/n242 ), .Y(\us01/n205 ) );
  AND2X1 \us01/U363  ( .A(\us01/n189 ), .B(\us01/n205 ), .Y(\us01/n65 ) );
  NOR2X1 \us01/U362  ( .A(\us01/n226 ), .B(\us01/n47 ), .Y(\us01/n45 ) );
  NOR2X1 \us01/U361  ( .A(\us01/n259 ), .B(\us01/n45 ), .Y(\us01/n73 ) );
  NAND2BX1 \us01/U360  ( .AN(\us01/n73 ), .B(\us01/n6 ), .Y(\us01/n158 ) );
  NOR2X1 \us01/U359  ( .A(\us01/n226 ), .B(\us01/n159 ), .Y(\us01/n95 ) );
  INVX1 \us01/U358  ( .A(\us01/n95 ), .Y(\us01/n111 ) );
  NOR2X1 \us01/U357  ( .A(\us01/n145 ), .B(sa01[1]), .Y(\us01/n42 ) );
  INVX1 \us01/U356  ( .A(\us01/n42 ), .Y(\us01/n121 ) );
  INVX1 \us01/U355  ( .A(\us01/n47 ), .Y(\us01/n96 ) );
  OAI211X1 \us01/U354  ( .A0(\us01/n65 ), .A1(\us01/n27 ), .B0(\us01/n158 ), 
        .C0(\us01/n358 ), .Y(\us01/n355 ) );
  NOR2X1 \us01/U353  ( .A(\us01/n226 ), .B(\us01/n145 ), .Y(\us01/n59 ) );
  NOR2X1 \us01/U352  ( .A(\us01/n96 ), .B(\us01/n59 ), .Y(\us01/n271 ) );
  NOR2X1 \us01/U351  ( .A(\us01/n226 ), .B(\us01/n278 ), .Y(\us01/n217 ) );
  INVX1 \us01/U350  ( .A(\us01/n217 ), .Y(\us01/n150 ) );
  NAND2X1 \us01/U349  ( .A(\us01/n44 ), .B(\us01/n150 ), .Y(\us01/n147 ) );
  NAND2X1 \us01/U348  ( .A(sa01[4]), .B(\us01/n226 ), .Y(\us01/n101 ) );
  INVX1 \us01/U347  ( .A(\us01/n159 ), .Y(\us01/n188 ) );
  NOR2X1 \us01/U346  ( .A(\us01/n188 ), .B(\us01/n226 ), .Y(\us01/n25 ) );
  INVX1 \us01/U345  ( .A(\us01/n172 ), .Y(\us01/n107 ) );
  AOI22X1 \us01/U344  ( .A0(\us01/n33 ), .A1(\us01/n147 ), .B0(\us01/n24 ), 
        .B1(\us01/n107 ), .Y(\us01/n357 ) );
  OAI221XL \us01/U343  ( .A0(\us01/n18 ), .A1(\us01/n121 ), .B0(\us01/n271 ), 
        .B1(\us01/n20 ), .C0(\us01/n357 ), .Y(\us01/n356 ) );
  MXI2X1 \us01/U342  ( .A(\us01/n355 ), .B(\us01/n356 ), .S0(\us01/n252 ), .Y(
        \us01/n331 ) );
  INVX1 \us01/U341  ( .A(\us01/n59 ), .Y(\us01/n79 ) );
  AND2X1 \us01/U340  ( .A(\us01/n101 ), .B(\us01/n79 ), .Y(\us01/n325 ) );
  XNOR2X1 \us01/U339  ( .A(sa01[5]), .B(\us01/n226 ), .Y(\us01/n352 ) );
  NOR2X1 \us01/U338  ( .A(\us01/n226 ), .B(\us01/n136 ), .Y(\us01/n281 ) );
  INVX1 \us01/U337  ( .A(\us01/n281 ), .Y(\us01/n19 ) );
  NAND2X1 \us01/U336  ( .A(\us01/n145 ), .B(\us01/n226 ), .Y(\us01/n223 ) );
  AOI21X1 \us01/U335  ( .A0(\us01/n19 ), .A1(\us01/n223 ), .B0(\us01/n27 ), 
        .Y(\us01/n354 ) );
  AOI31X1 \us01/U334  ( .A0(\us01/n6 ), .A1(\us01/n352 ), .A2(\us01/n259 ), 
        .B0(\us01/n354 ), .Y(\us01/n353 ) );
  OAI221XL \us01/U333  ( .A0(\us01/n20 ), .A1(\us01/n34 ), .B0(\us01/n325 ), 
        .B1(\us01/n4 ), .C0(\us01/n353 ), .Y(\us01/n347 ) );
  INVX1 \us01/U332  ( .A(\us01/n352 ), .Y(\us01/n349 ) );
  NAND2X1 \us01/U331  ( .A(\us01/n278 ), .B(\us01/n6 ), .Y(\us01/n74 ) );
  OAI211X1 \us01/U330  ( .A0(\us01/n349 ), .A1(\us01/n74 ), .B0(\us01/n350 ), 
        .C0(\us01/n351 ), .Y(\us01/n348 ) );
  MXI2X1 \us01/U329  ( .A(\us01/n347 ), .B(\us01/n348 ), .S0(\us01/n252 ), .Y(
        \us01/n332 ) );
  NOR2X1 \us01/U328  ( .A(\us01/n44 ), .B(\us01/n226 ), .Y(\us01/n157 ) );
  INVX1 \us01/U327  ( .A(\us01/n157 ), .Y(\us01/n240 ) );
  NAND2X1 \us01/U326  ( .A(\us01/n240 ), .B(\us01/n189 ), .Y(\us01/n68 ) );
  NOR2X1 \us01/U325  ( .A(\us01/n20 ), .B(\us01/n159 ), .Y(\us01/n225 ) );
  NOR2X1 \us01/U324  ( .A(\us01/n225 ), .B(\us01/n40 ), .Y(\us01/n345 ) );
  INVX1 \us01/U323  ( .A(\us01/n278 ), .Y(\us01/n94 ) );
  NAND2X1 \us01/U322  ( .A(\us01/n94 ), .B(\us01/n226 ), .Y(\us01/n199 ) );
  NAND2X1 \us01/U321  ( .A(\us01/n199 ), .B(\us01/n205 ), .Y(\us01/n82 ) );
  NAND2X1 \us01/U320  ( .A(\us01/n19 ), .B(\us01/n199 ), .Y(\us01/n295 ) );
  NOR2X1 \us01/U319  ( .A(\us01/n226 ), .B(\us01/n259 ), .Y(\us01/n210 ) );
  NOR2X1 \us01/U318  ( .A(\us01/n27 ), .B(\us01/n210 ), .Y(\us01/n173 ) );
  MXI2X1 \us01/U317  ( .A(\us01/n345 ), .B(\us01/n346 ), .S0(\us01/n252 ), .Y(
        \us01/n342 ) );
  NOR2X1 \us01/U316  ( .A(sa01[1]), .B(sa01[3]), .Y(\us01/n163 ) );
  INVX1 \us01/U315  ( .A(\us01/n163 ), .Y(\us01/n37 ) );
  INVX1 \us01/U314  ( .A(\us01/n173 ), .Y(\us01/n344 ) );
  AOI21X1 \us01/U313  ( .A0(\us01/n240 ), .A1(\us01/n37 ), .B0(\us01/n344 ), 
        .Y(\us01/n343 ) );
  AOI211X1 \us01/U312  ( .A0(\us01/n5 ), .A1(\us01/n68 ), .B0(\us01/n342 ), 
        .C0(\us01/n343 ), .Y(\us01/n333 ) );
  NOR2X1 \us01/U311  ( .A(\us01/n18 ), .B(\us01/n226 ), .Y(\us01/n258 ) );
  NAND2X1 \us01/U310  ( .A(\us01/n278 ), .B(sa01[1]), .Y(\us01/n204 ) );
  NOR2X1 \us01/U309  ( .A(\us01/n188 ), .B(sa01[1]), .Y(\us01/n179 ) );
  INVX1 \us01/U308  ( .A(\us01/n179 ), .Y(\us01/n330 ) );
  NAND2X1 \us01/U307  ( .A(\us01/n204 ), .B(\us01/n330 ), .Y(\us01/n239 ) );
  NOR2X1 \us01/U306  ( .A(\us01/n136 ), .B(sa01[1]), .Y(\us01/n299 ) );
  NOR2X1 \us01/U305  ( .A(\us01/n299 ), .B(\us01/n210 ), .Y(\us01/n341 ) );
  OAI32X1 \us01/U304  ( .A0(\us01/n27 ), .A1(\us01/n278 ), .A2(\us01/n95 ), 
        .B0(\us01/n341 ), .B1(\us01/n4 ), .Y(\us01/n340 ) );
  INVX1 \us01/U303  ( .A(\us01/n45 ), .Y(\us01/n126 ) );
  NAND2X1 \us01/U302  ( .A(\us01/n126 ), .B(\us01/n101 ), .Y(\us01/n178 ) );
  NOR2X1 \us01/U301  ( .A(\us01/n18 ), .B(\us01/n136 ), .Y(\us01/n280 ) );
  OAI21XL \us01/U300  ( .A0(\us01/n4 ), .A1(\us01/n121 ), .B0(\us01/n339 ), 
        .Y(\us01/n338 ) );
  MXI2X1 \us01/U299  ( .A(\us01/n336 ), .B(\us01/n337 ), .S0(\us01/n252 ), .Y(
        \us01/n335 ) );
  NOR2X1 \us01/U298  ( .A(\us01/n258 ), .B(\us01/n335 ), .Y(\us01/n334 ) );
  MX4X1 \us01/U297  ( .A(\us01/n331 ), .B(\us01/n332 ), .C(\us01/n333 ), .D(
        \us01/n334 ), .S0(sa01[6]), .S1(\us01/n234 ), .Y(sa01_sr[0]) );
  INVX1 \us01/U296  ( .A(\us01/n299 ), .Y(\us01/n80 ) );
  NOR2X1 \us01/U295  ( .A(\us01/n111 ), .B(\us01/n18 ), .Y(\us01/n269 ) );
  INVX1 \us01/U294  ( .A(\us01/n269 ), .Y(\us01/n75 ) );
  OAI221XL \us01/U293  ( .A0(\us01/n18 ), .A1(\us01/n330 ), .B0(\us01/n20 ), 
        .B1(\us01/n80 ), .C0(\us01/n75 ), .Y(\us01/n329 ) );
  AOI221X1 \us01/U292  ( .A0(\us01/n325 ), .A1(\us01/n33 ), .B0(\us01/n24 ), 
        .B1(\us01/n303 ), .C0(\us01/n329 ), .Y(\us01/n319 ) );
  NOR2X1 \us01/U291  ( .A(\us01/n234 ), .B(sa01[5]), .Y(\us01/n14 ) );
  NOR2X1 \us01/U290  ( .A(\us01/n25 ), .B(\us01/n299 ), .Y(\us01/n313 ) );
  NAND2X1 \us01/U289  ( .A(\us01/n44 ), .B(\us01/n226 ), .Y(\us01/n300 ) );
  AND2X1 \us01/U288  ( .A(\us01/n300 ), .B(\us01/n240 ), .Y(\us01/n23 ) );
  OAI32X1 \us01/U287  ( .A0(\us01/n4 ), .A1(\us01/n145 ), .A2(\us01/n210 ), 
        .B0(\us01/n137 ), .B1(\us01/n27 ), .Y(\us01/n328 ) );
  NOR2X1 \us01/U286  ( .A(sa01[0]), .B(sa01[5]), .Y(\us01/n16 ) );
  INVX1 \us01/U285  ( .A(\us01/n16 ), .Y(\us01/n114 ) );
  INVX1 \us01/U284  ( .A(\us01/n145 ), .Y(\us01/n149 ) );
  NOR2X1 \us01/U283  ( .A(\us01/n47 ), .B(sa01[1]), .Y(\us01/n98 ) );
  INVX1 \us01/U282  ( .A(\us01/n98 ), .Y(\us01/n284 ) );
  OAI21XL \us01/U281  ( .A0(\us01/n69 ), .A1(\us01/n284 ), .B0(\us01/n27 ), 
        .Y(\us01/n327 ) );
  AOI31X1 \us01/U280  ( .A0(\us01/n111 ), .A1(\us01/n149 ), .A2(\us01/n327 ), 
        .B0(\us01/n225 ), .Y(\us01/n326 ) );
  OAI21XL \us01/U279  ( .A0(\us01/n325 ), .A1(\us01/n18 ), .B0(\us01/n326 ), 
        .Y(\us01/n322 ) );
  NAND2X1 \us01/U278  ( .A(\us01/n19 ), .B(\us01/n189 ), .Y(\us01/n71 ) );
  NOR2X1 \us01/U277  ( .A(\us01/n71 ), .B(\us01/n18 ), .Y(\us01/n135 ) );
  AOI21X1 \us01/U276  ( .A0(\us01/n40 ), .A1(sa01[4]), .B0(\us01/n135 ), .Y(
        \us01/n324 ) );
  OAI221XL \us01/U275  ( .A0(\us01/n47 ), .A1(\us01/n27 ), .B0(\us01/n65 ), 
        .B1(\us01/n20 ), .C0(\us01/n324 ), .Y(\us01/n323 ) );
  AOI22X1 \us01/U274  ( .A0(\us01/n55 ), .A1(\us01/n322 ), .B0(\us01/n89 ), 
        .B1(\us01/n323 ), .Y(\us01/n321 ) );
  OAI221XL \us01/U273  ( .A0(\us01/n319 ), .A1(\us01/n52 ), .B0(\us01/n320 ), 
        .B1(\us01/n114 ), .C0(\us01/n321 ), .Y(\us01/n304 ) );
  NOR2X1 \us01/U272  ( .A(\us01/n226 ), .B(\us01/n58 ), .Y(\us01/n290 ) );
  INVX1 \us01/U271  ( .A(\us01/n290 ), .Y(\us01/n200 ) );
  NAND2X1 \us01/U270  ( .A(\us01/n34 ), .B(\us01/n200 ), .Y(\us01/n120 ) );
  INVX1 \us01/U269  ( .A(\us01/n210 ), .Y(\us01/n100 ) );
  OAI221XL \us01/U268  ( .A0(\us01/n20 ), .A1(\us01/n100 ), .B0(sa01[3]), .B1(
        \us01/n4 ), .C0(\us01/n262 ), .Y(\us01/n317 ) );
  INVX1 \us01/U267  ( .A(\us01/n258 ), .Y(\us01/n182 ) );
  AOI211X1 \us01/U266  ( .A0(\us01/n33 ), .A1(\us01/n120 ), .B0(\us01/n317 ), 
        .C0(\us01/n318 ), .Y(\us01/n306 ) );
  NAND2X1 \us01/U265  ( .A(\us01/n100 ), .B(\us01/n199 ), .Y(\us01/n151 ) );
  INVX1 \us01/U264  ( .A(\us01/n151 ), .Y(\us01/n314 ) );
  NOR2X1 \us01/U263  ( .A(\us01/n45 ), .B(\us01/n163 ), .Y(\us01/n160 ) );
  INVX1 \us01/U262  ( .A(\us01/n295 ), .Y(\us01/n92 ) );
  AOI21X1 \us01/U261  ( .A0(sa01[1]), .A1(\us01/n58 ), .B0(\us01/n98 ), .Y(
        \us01/n316 ) );
  OAI22X1 \us01/U260  ( .A0(\us01/n92 ), .A1(\us01/n18 ), .B0(\us01/n316 ), 
        .B1(\us01/n27 ), .Y(\us01/n315 ) );
  NOR2X1 \us01/U259  ( .A(\us01/n149 ), .B(\us01/n226 ), .Y(\us01/n41 ) );
  INVX1 \us01/U258  ( .A(\us01/n41 ), .Y(\us01/n105 ) );
  NAND2X1 \us01/U257  ( .A(\us01/n284 ), .B(\us01/n105 ), .Y(\us01/n227 ) );
  AOI21X1 \us01/U256  ( .A0(\us01/n313 ), .A1(\us01/n33 ), .B0(\us01/n269 ), 
        .Y(\us01/n312 ) );
  OAI221XL \us01/U255  ( .A0(\us01/n149 ), .A1(\us01/n20 ), .B0(\us01/n4 ), 
        .B1(\us01/n227 ), .C0(\us01/n312 ), .Y(\us01/n309 ) );
  AOI21X1 \us01/U254  ( .A0(\us01/n226 ), .A1(\us01/n188 ), .B0(\us01/n242 ), 
        .Y(\us01/n185 ) );
  INVX1 \us01/U253  ( .A(\us01/n185 ), .Y(\us01/n48 ) );
  AND2X1 \us01/U252  ( .A(\us01/n223 ), .B(\us01/n240 ), .Y(\us01/n28 ) );
  OAI221XL \us01/U251  ( .A0(\us01/n27 ), .A1(\us01/n44 ), .B0(\us01/n4 ), 
        .B1(\us01/n48 ), .C0(\us01/n311 ), .Y(\us01/n310 ) );
  AOI22X1 \us01/U250  ( .A0(\us01/n89 ), .A1(\us01/n309 ), .B0(\us01/n55 ), 
        .B1(\us01/n310 ), .Y(\us01/n308 ) );
  OAI221XL \us01/U249  ( .A0(\us01/n306 ), .A1(\us01/n52 ), .B0(\us01/n307 ), 
        .B1(\us01/n114 ), .C0(\us01/n308 ), .Y(\us01/n305 ) );
  MX2X1 \us01/U248  ( .A(\us01/n304 ), .B(\us01/n305 ), .S0(sa01[6]), .Y(
        sa01_sr[1]) );
  INVX1 \us01/U247  ( .A(\us01/n187 ), .Y(\us01/n61 ) );
  MXI2X1 \us01/U246  ( .A(\us01/n303 ), .B(\us01/n61 ), .S0(\us01/n69 ), .Y(
        \us01/n301 ) );
  MXI2X1 \us01/U245  ( .A(\us01/n301 ), .B(\us01/n147 ), .S0(\us01/n302 ), .Y(
        \us01/n285 ) );
  NAND2X1 \us01/U244  ( .A(\us01/n200 ), .B(\us01/n300 ), .Y(\us01/n99 ) );
  INVX1 \us01/U243  ( .A(\us01/n99 ), .Y(\us01/n296 ) );
  NOR2X1 \us01/U242  ( .A(\us01/n299 ), .B(\us01/n242 ), .Y(\us01/n298 ) );
  NAND2X1 \us01/U241  ( .A(sa01[1]), .B(\us01/n47 ), .Y(\us01/n122 ) );
  NOR2X1 \us01/U240  ( .A(\us01/n159 ), .B(\us01/n217 ), .Y(\us01/n198 ) );
  OAI221XL \us01/U239  ( .A0(\us01/n298 ), .A1(\us01/n27 ), .B0(\us01/n20 ), 
        .B1(\us01/n122 ), .C0(\us01/n132 ), .Y(\us01/n297 ) );
  AOI221X1 \us01/U238  ( .A0(\us01/n225 ), .A1(\us01/n226 ), .B0(\us01/n296 ), 
        .B1(\us01/n6 ), .C0(\us01/n297 ), .Y(\us01/n291 ) );
  OAI2BB2X1 \us01/U237  ( .B0(\us01/n27 ), .B1(\us01/n295 ), .A0N(\us01/n34 ), 
        .A1N(\us01/n24 ), .Y(\us01/n293 ) );
  AOI21X1 \us01/U236  ( .A0(\us01/n101 ), .A1(\us01/n150 ), .B0(\us01/n20 ), 
        .Y(\us01/n294 ) );
  AOI211X1 \us01/U235  ( .A0(\us01/n5 ), .A1(\us01/n79 ), .B0(\us01/n293 ), 
        .C0(\us01/n294 ), .Y(\us01/n292 ) );
  INVX1 \us01/U234  ( .A(\us01/n89 ), .Y(\us01/n10 ) );
  OAI22X1 \us01/U233  ( .A0(\us01/n291 ), .A1(\us01/n114 ), .B0(\us01/n292 ), 
        .B1(\us01/n10 ), .Y(\us01/n286 ) );
  INVX1 \us01/U232  ( .A(\us01/n225 ), .Y(\us01/n288 ) );
  NAND2X1 \us01/U231  ( .A(\us01/n200 ), .B(\us01/n284 ), .Y(\us01/n102 ) );
  NOR2X1 \us01/U230  ( .A(\us01/n290 ), .B(\us01/n163 ), .Y(\us01/n184 ) );
  AOI22X1 \us01/U229  ( .A0(\us01/n102 ), .A1(\us01/n69 ), .B0(\us01/n184 ), 
        .B1(\us01/n33 ), .Y(\us01/n289 ) );
  AOI31X1 \us01/U228  ( .A0(\us01/n132 ), .A1(\us01/n288 ), .A2(\us01/n289 ), 
        .B0(\us01/n52 ), .Y(\us01/n287 ) );
  AOI211X1 \us01/U227  ( .A0(\us01/n285 ), .A1(\us01/n55 ), .B0(\us01/n286 ), 
        .C0(\us01/n287 ), .Y(\us01/n263 ) );
  NAND2X1 \us01/U226  ( .A(\us01/n284 ), .B(\us01/n122 ), .Y(\us01/n125 ) );
  NOR2X1 \us01/U225  ( .A(\us01/n199 ), .B(\us01/n4 ), .Y(\us01/n50 ) );
  AOI21X1 \us01/U224  ( .A0(\us01/n200 ), .A1(\us01/n223 ), .B0(\us01/n20 ), 
        .Y(\us01/n283 ) );
  AOI211X1 \us01/U223  ( .A0(\us01/n5 ), .A1(\us01/n125 ), .B0(\us01/n50 ), 
        .C0(\us01/n283 ), .Y(\us01/n282 ) );
  OAI221XL \us01/U222  ( .A0(\us01/n281 ), .A1(\us01/n27 ), .B0(\us01/n4 ), 
        .B1(\us01/n111 ), .C0(\us01/n282 ), .Y(\us01/n265 ) );
  INVX1 \us01/U221  ( .A(\us01/n280 ), .Y(\us01/n247 ) );
  NAND2X1 \us01/U220  ( .A(\us01/n41 ), .B(\us01/n33 ), .Y(\us01/n272 ) );
  OAI221XL \us01/U219  ( .A0(sa01[1]), .A1(\us01/n247 ), .B0(\us01/n4 ), .B1(
        \us01/n189 ), .C0(\us01/n272 ), .Y(\us01/n279 ) );
  NAND2X1 \us01/U218  ( .A(sa01[2]), .B(\us01/n149 ), .Y(\us01/n276 ) );
  XNOR2X1 \us01/U217  ( .A(\us01/n129 ), .B(sa01[1]), .Y(\us01/n155 ) );
  MXI2X1 \us01/U216  ( .A(\us01/n276 ), .B(\us01/n277 ), .S0(\us01/n155 ), .Y(
        \us01/n275 ) );
  OAI22X1 \us01/U215  ( .A0(\us01/n273 ), .A1(\us01/n10 ), .B0(\us01/n274 ), 
        .B1(\us01/n52 ), .Y(\us01/n266 ) );
  NOR2X1 \us01/U214  ( .A(\us01/n20 ), .B(\us01/n226 ), .Y(\us01/n176 ) );
  OAI21XL \us01/U213  ( .A0(\us01/n4 ), .A1(\us01/n271 ), .B0(\us01/n272 ), 
        .Y(\us01/n270 ) );
  OAI31X1 \us01/U212  ( .A0(\us01/n176 ), .A1(\us01/n269 ), .A2(\us01/n270 ), 
        .B0(\us01/n16 ), .Y(\us01/n268 ) );
  INVX1 \us01/U211  ( .A(\us01/n268 ), .Y(\us01/n267 ) );
  AOI211X1 \us01/U210  ( .A0(\us01/n55 ), .A1(\us01/n265 ), .B0(\us01/n266 ), 
        .C0(\us01/n267 ), .Y(\us01/n264 ) );
  MXI2X1 \us01/U209  ( .A(\us01/n263 ), .B(\us01/n264 ), .S0(sa01[6]), .Y(
        sa01_sr[2]) );
  NOR2X1 \us01/U208  ( .A(\us01/n94 ), .B(sa01[1]), .Y(\us01/n211 ) );
  INVX1 \us01/U207  ( .A(\us01/n262 ), .Y(\us01/n261 ) );
  AOI211X1 \us01/U206  ( .A0(\us01/n259 ), .A1(\us01/n24 ), .B0(\us01/n260 ), 
        .C0(\us01/n261 ), .Y(\us01/n255 ) );
  OAI22X1 \us01/U205  ( .A0(\us01/n20 ), .A1(\us01/n68 ), .B0(\us01/n27 ), 
        .B1(\us01/n37 ), .Y(\us01/n257 ) );
  NOR3X1 \us01/U204  ( .A(\us01/n257 ), .B(\us01/n258 ), .C(\us01/n50 ), .Y(
        \us01/n256 ) );
  MXI2X1 \us01/U203  ( .A(\us01/n255 ), .B(\us01/n256 ), .S0(\us01/n252 ), .Y(
        \us01/n254 ) );
  AOI221X1 \us01/U202  ( .A0(\us01/n211 ), .A1(\us01/n5 ), .B0(\us01/n40 ), 
        .B1(sa01[4]), .C0(\us01/n254 ), .Y(\us01/n248 ) );
  INVX1 \us01/U201  ( .A(\us01/n211 ), .Y(\us01/n106 ) );
  NAND2X1 \us01/U200  ( .A(\us01/n200 ), .B(\us01/n106 ), .Y(\us01/n83 ) );
  NAND2X1 \us01/U199  ( .A(\us01/n199 ), .B(\us01/n204 ), .Y(\us01/n169 ) );
  AOI2BB2X1 \us01/U198  ( .B0(\us01/n65 ), .B1(\us01/n24 ), .A0N(\us01/n169 ), 
        .A1N(\us01/n20 ), .Y(\us01/n253 ) );
  OAI221XL \us01/U197  ( .A0(\us01/n172 ), .A1(\us01/n18 ), .B0(\us01/n27 ), 
        .B1(\us01/n83 ), .C0(\us01/n253 ), .Y(\us01/n251 ) );
  MXI2X1 \us01/U196  ( .A(\us01/n250 ), .B(\us01/n251 ), .S0(\us01/n252 ), .Y(
        \us01/n249 ) );
  MXI2X1 \us01/U195  ( .A(\us01/n248 ), .B(\us01/n249 ), .S0(\us01/n234 ), .Y(
        \us01/n228 ) );
  OAI21XL \us01/U194  ( .A0(\us01/n58 ), .A1(\us01/n27 ), .B0(\us01/n247 ), 
        .Y(\us01/n245 ) );
  NOR2X1 \us01/U193  ( .A(sa01[7]), .B(\us01/n145 ), .Y(\us01/n246 ) );
  XNOR2X1 \us01/U192  ( .A(\us01/n69 ), .B(sa01[1]), .Y(\us01/n130 ) );
  MXI2X1 \us01/U191  ( .A(\us01/n245 ), .B(\us01/n246 ), .S0(\us01/n130 ), .Y(
        \us01/n243 ) );
  OAI211X1 \us01/U190  ( .A0(\us01/n4 ), .A1(\us01/n149 ), .B0(\us01/n243 ), 
        .C0(\us01/n244 ), .Y(\us01/n230 ) );
  NOR2X1 \us01/U189  ( .A(\us01/n242 ), .B(\us01/n137 ), .Y(\us01/n70 ) );
  OAI221XL \us01/U188  ( .A0(\us01/n159 ), .A1(\us01/n27 ), .B0(\us01/n20 ), 
        .B1(\us01/n34 ), .C0(\us01/n241 ), .Y(\us01/n231 ) );
  NAND2X1 \us01/U187  ( .A(\us01/n101 ), .B(\us01/n240 ), .Y(\us01/n76 ) );
  AOI21X1 \us01/U186  ( .A0(\us01/n122 ), .A1(\us01/n106 ), .B0(\us01/n129 ), 
        .Y(\us01/n237 ) );
  INVX1 \us01/U185  ( .A(\us01/n239 ), .Y(\us01/n238 ) );
  OAI21XL \us01/U184  ( .A0(\us01/n237 ), .A1(\us01/n43 ), .B0(\us01/n238 ), 
        .Y(\us01/n236 ) );
  OAI221XL \us01/U183  ( .A0(\us01/n18 ), .A1(\us01/n76 ), .B0(\us01/n59 ), 
        .B1(\us01/n27 ), .C0(\us01/n236 ), .Y(\us01/n232 ) );
  AOI2BB2X1 \us01/U182  ( .B0(\us01/n24 ), .B1(\us01/n187 ), .A0N(\us01/n227 ), 
        .A1N(\us01/n20 ), .Y(\us01/n235 ) );
  OAI211X1 \us01/U181  ( .A0(\us01/n27 ), .A1(\us01/n122 ), .B0(\us01/n158 ), 
        .C0(\us01/n235 ), .Y(\us01/n233 ) );
  MX4X1 \us01/U180  ( .A(\us01/n230 ), .B(\us01/n231 ), .C(\us01/n232 ), .D(
        \us01/n233 ), .S0(\us01/n234 ), .S1(sa01[5]), .Y(\us01/n229 ) );
  MX2X1 \us01/U179  ( .A(\us01/n228 ), .B(\us01/n229 ), .S0(sa01[6]), .Y(
        sa01_sr[3]) );
  NOR2BX1 \us01/U178  ( .AN(\us01/n204 ), .B(\us01/n137 ), .Y(\us01/n110 ) );
  INVX1 \us01/U177  ( .A(\us01/n110 ), .Y(\us01/n64 ) );
  AOI22X1 \us01/U176  ( .A0(\us01/n225 ), .A1(\us01/n226 ), .B0(\us01/n6 ), 
        .B1(\us01/n227 ), .Y(\us01/n224 ) );
  OAI221XL \us01/U175  ( .A0(\us01/n27 ), .A1(\us01/n64 ), .B0(\us01/n4 ), 
        .B1(\us01/n83 ), .C0(\us01/n224 ), .Y(\us01/n212 ) );
  NAND2X1 \us01/U174  ( .A(\us01/n34 ), .B(\us01/n204 ), .Y(\us01/n221 ) );
  OAI21XL \us01/U173  ( .A0(\us01/n69 ), .A1(\us01/n223 ), .B0(\us01/n27 ), 
        .Y(\us01/n222 ) );
  NOR2X1 \us01/U172  ( .A(\us01/n217 ), .B(\us01/n42 ), .Y(\us01/n208 ) );
  AOI211X1 \us01/U171  ( .A0(\us01/n208 ), .A1(\us01/n5 ), .B0(\us01/n220 ), 
        .C0(\us01/n173 ), .Y(\us01/n219 ) );
  OAI22X1 \us01/U170  ( .A0(\us01/n218 ), .A1(\us01/n10 ), .B0(\us01/n219 ), 
        .B1(\us01/n114 ), .Y(\us01/n213 ) );
  INVX1 \us01/U169  ( .A(\us01/n135 ), .Y(\us01/n215 ) );
  NOR2X1 \us01/U168  ( .A(\us01/n4 ), .B(\us01/n159 ), .Y(\us01/n31 ) );
  INVX1 \us01/U167  ( .A(\us01/n31 ), .Y(\us01/n196 ) );
  AOI31X1 \us01/U166  ( .A0(\us01/n215 ), .A1(\us01/n196 ), .A2(\us01/n216 ), 
        .B0(\us01/n52 ), .Y(\us01/n214 ) );
  AOI211X1 \us01/U165  ( .A0(\us01/n55 ), .A1(\us01/n212 ), .B0(\us01/n213 ), 
        .C0(\us01/n214 ), .Y(\us01/n190 ) );
  INVX1 \us01/U164  ( .A(\us01/n207 ), .Y(\us01/n192 ) );
  NOR2X1 \us01/U163  ( .A(\us01/n25 ), .B(\us01/n98 ), .Y(\us01/n32 ) );
  OAI22X1 \us01/U162  ( .A0(\us01/n28 ), .A1(\us01/n4 ), .B0(\us01/n188 ), 
        .B1(\us01/n27 ), .Y(\us01/n206 ) );
  NAND2X1 \us01/U161  ( .A(\us01/n204 ), .B(\us01/n80 ), .Y(\us01/n118 ) );
  INVX1 \us01/U160  ( .A(\us01/n118 ), .Y(\us01/n123 ) );
  NAND2X1 \us01/U159  ( .A(\us01/n94 ), .B(\us01/n79 ), .Y(\us01/n203 ) );
  OAI2BB1X1 \us01/U158  ( .A0N(\us01/n199 ), .A1N(\us01/n200 ), .B0(\us01/n33 ), .Y(\us01/n195 ) );
  INVX1 \us01/U157  ( .A(\us01/n55 ), .Y(\us01/n12 ) );
  AOI31X1 \us01/U156  ( .A0(\us01/n195 ), .A1(\us01/n196 ), .A2(\us01/n197 ), 
        .B0(\us01/n12 ), .Y(\us01/n194 ) );
  AOI211X1 \us01/U155  ( .A0(\us01/n89 ), .A1(\us01/n192 ), .B0(\us01/n193 ), 
        .C0(\us01/n194 ), .Y(\us01/n191 ) );
  MXI2X1 \us01/U154  ( .A(\us01/n190 ), .B(\us01/n191 ), .S0(sa01[6]), .Y(
        sa01_sr[4]) );
  OAI21XL \us01/U153  ( .A0(\us01/n69 ), .A1(\us01/n189 ), .B0(\us01/n27 ), 
        .Y(\us01/n186 ) );
  INVX1 \us01/U152  ( .A(\us01/n183 ), .Y(\us01/n180 ) );
  NAND2X1 \us01/U151  ( .A(\us01/n74 ), .B(\us01/n182 ), .Y(\us01/n181 ) );
  AOI211X1 \us01/U150  ( .A0(\us01/n179 ), .A1(\us01/n24 ), .B0(\us01/n180 ), 
        .C0(\us01/n181 ), .Y(\us01/n165 ) );
  INVX1 \us01/U149  ( .A(\us01/n178 ), .Y(\us01/n175 ) );
  AOI211X1 \us01/U148  ( .A0(\us01/n175 ), .A1(\us01/n5 ), .B0(\us01/n176 ), 
        .C0(\us01/n177 ), .Y(\us01/n174 ) );
  OAI221XL \us01/U147  ( .A0(\us01/n159 ), .A1(\us01/n27 ), .B0(\us01/n145 ), 
        .B1(\us01/n20 ), .C0(\us01/n174 ), .Y(\us01/n167 ) );
  MXI2X1 \us01/U146  ( .A(\us01/n40 ), .B(\us01/n173 ), .S0(\us01/n96 ), .Y(
        \us01/n170 ) );
  AOI22X1 \us01/U145  ( .A0(\us01/n137 ), .A1(\us01/n24 ), .B0(\us01/n172 ), 
        .B1(\us01/n6 ), .Y(\us01/n171 ) );
  OAI211X1 \us01/U144  ( .A0(\us01/n20 ), .A1(\us01/n169 ), .B0(\us01/n170 ), 
        .C0(\us01/n171 ), .Y(\us01/n168 ) );
  AOI22X1 \us01/U143  ( .A0(\us01/n89 ), .A1(\us01/n167 ), .B0(\us01/n55 ), 
        .B1(\us01/n168 ), .Y(\us01/n166 ) );
  OAI221XL \us01/U142  ( .A0(\us01/n164 ), .A1(\us01/n114 ), .B0(\us01/n165 ), 
        .B1(\us01/n52 ), .C0(\us01/n166 ), .Y(\us01/n138 ) );
  OAI21XL \us01/U141  ( .A0(\us01/n41 ), .A1(\us01/n163 ), .B0(\us01/n69 ), 
        .Y(\us01/n162 ) );
  AOI221X1 \us01/U140  ( .A0(\us01/n159 ), .A1(\us01/n24 ), .B0(\us01/n160 ), 
        .B1(\us01/n33 ), .C0(\us01/n161 ), .Y(\us01/n140 ) );
  OAI21XL \us01/U139  ( .A0(\us01/n157 ), .A1(\us01/n20 ), .B0(\us01/n158 ), 
        .Y(\us01/n156 ) );
  NOR2X1 \us01/U138  ( .A(\us01/n4 ), .B(\us01/n136 ), .Y(\us01/n153 ) );
  NOR2X1 \us01/U137  ( .A(\us01/n145 ), .B(\us01/n69 ), .Y(\us01/n154 ) );
  MXI2X1 \us01/U136  ( .A(\us01/n153 ), .B(\us01/n154 ), .S0(\us01/n155 ), .Y(
        \us01/n152 ) );
  OAI221XL \us01/U135  ( .A0(\us01/n110 ), .A1(\us01/n18 ), .B0(\us01/n20 ), 
        .B1(\us01/n151 ), .C0(\us01/n152 ), .Y(\us01/n143 ) );
  AOI21X1 \us01/U134  ( .A0(\us01/n149 ), .A1(\us01/n150 ), .B0(\us01/n18 ), 
        .Y(\us01/n148 ) );
  AOI2BB1X1 \us01/U133  ( .A0N(\us01/n147 ), .A1N(\us01/n27 ), .B0(\us01/n148 ), .Y(\us01/n146 ) );
  OAI221XL \us01/U132  ( .A0(\us01/n145 ), .A1(\us01/n20 ), .B0(\us01/n4 ), 
        .B1(\us01/n34 ), .C0(\us01/n146 ), .Y(\us01/n144 ) );
  AOI22X1 \us01/U131  ( .A0(\us01/n89 ), .A1(\us01/n143 ), .B0(\us01/n14 ), 
        .B1(\us01/n144 ), .Y(\us01/n142 ) );
  OAI221XL \us01/U130  ( .A0(\us01/n140 ), .A1(\us01/n12 ), .B0(\us01/n141 ), 
        .B1(\us01/n114 ), .C0(\us01/n142 ), .Y(\us01/n139 ) );
  MX2X1 \us01/U129  ( .A(\us01/n138 ), .B(\us01/n139 ), .S0(sa01[6]), .Y(
        sa01_sr[5]) );
  INVX1 \us01/U128  ( .A(\us01/n70 ), .Y(\us01/n133 ) );
  OAI22X1 \us01/U127  ( .A0(\us01/n4 ), .A1(\us01/n136 ), .B0(\us01/n137 ), 
        .B1(\us01/n27 ), .Y(\us01/n134 ) );
  AOI211X1 \us01/U126  ( .A0(\us01/n133 ), .A1(\us01/n69 ), .B0(\us01/n134 ), 
        .C0(\us01/n135 ), .Y(\us01/n112 ) );
  INVX1 \us01/U125  ( .A(\us01/n132 ), .Y(\us01/n131 ) );
  OAI21XL \us01/U124  ( .A0(\us01/n18 ), .A1(\us01/n37 ), .B0(\us01/n128 ), 
        .Y(\us01/n127 ) );
  OAI221XL \us01/U123  ( .A0(\us01/n18 ), .A1(\us01/n105 ), .B0(\us01/n123 ), 
        .B1(\us01/n27 ), .C0(\us01/n124 ), .Y(\us01/n116 ) );
  NAND2X1 \us01/U122  ( .A(\us01/n121 ), .B(\us01/n122 ), .Y(\us01/n30 ) );
  OAI221XL \us01/U121  ( .A0(\us01/n18 ), .A1(\us01/n118 ), .B0(\us01/n27 ), 
        .B1(\us01/n30 ), .C0(\us01/n119 ), .Y(\us01/n117 ) );
  AOI22X1 \us01/U120  ( .A0(\us01/n89 ), .A1(\us01/n116 ), .B0(\us01/n55 ), 
        .B1(\us01/n117 ), .Y(\us01/n115 ) );
  OAI221XL \us01/U119  ( .A0(\us01/n112 ), .A1(\us01/n52 ), .B0(\us01/n113 ), 
        .B1(\us01/n114 ), .C0(\us01/n115 ), .Y(\us01/n84 ) );
  OAI22X1 \us01/U118  ( .A0(\us01/n110 ), .A1(\us01/n4 ), .B0(\us01/n20 ), 
        .B1(\us01/n21 ), .Y(\us01/n108 ) );
  AOI21X1 \us01/U117  ( .A0(sa01[1]), .A1(\us01/n58 ), .B0(\us01/n27 ), .Y(
        \us01/n109 ) );
  AOI211X1 \us01/U116  ( .A0(\us01/n5 ), .A1(\us01/n107 ), .B0(\us01/n108 ), 
        .C0(\us01/n109 ), .Y(\us01/n86 ) );
  OAI22X1 \us01/U115  ( .A0(\us01/n45 ), .A1(\us01/n4 ), .B0(sa01[4]), .B1(
        \us01/n18 ), .Y(\us01/n103 ) );
  AOI21X1 \us01/U114  ( .A0(\us01/n105 ), .A1(\us01/n106 ), .B0(\us01/n20 ), 
        .Y(\us01/n104 ) );
  AOI211X1 \us01/U113  ( .A0(\us01/n33 ), .A1(\us01/n102 ), .B0(\us01/n103 ), 
        .C0(\us01/n104 ), .Y(\us01/n87 ) );
  NAND2X1 \us01/U112  ( .A(\us01/n100 ), .B(\us01/n101 ), .Y(\us01/n62 ) );
  OAI221XL \us01/U111  ( .A0(\us01/n27 ), .A1(\us01/n62 ), .B0(\us01/n4 ), 
        .B1(\us01/n21 ), .C0(\us01/n97 ), .Y(\us01/n90 ) );
  NOR3X1 \us01/U110  ( .A(\us01/n4 ), .B(\us01/n95 ), .C(\us01/n96 ), .Y(
        \us01/n67 ) );
  AOI31X1 \us01/U109  ( .A0(\us01/n79 ), .A1(\us01/n94 ), .A2(\us01/n6 ), .B0(
        \us01/n67 ), .Y(\us01/n93 ) );
  OAI221XL \us01/U108  ( .A0(\us01/n73 ), .A1(\us01/n27 ), .B0(\us01/n92 ), 
        .B1(\us01/n20 ), .C0(\us01/n93 ), .Y(\us01/n91 ) );
  AOI22X1 \us01/U107  ( .A0(\us01/n89 ), .A1(\us01/n90 ), .B0(\us01/n16 ), 
        .B1(\us01/n91 ), .Y(\us01/n88 ) );
  OAI221XL \us01/U106  ( .A0(\us01/n86 ), .A1(\us01/n52 ), .B0(\us01/n87 ), 
        .B1(\us01/n12 ), .C0(\us01/n88 ), .Y(\us01/n85 ) );
  MX2X1 \us01/U105  ( .A(\us01/n84 ), .B(\us01/n85 ), .S0(sa01[6]), .Y(
        sa01_sr[6]) );
  INVX1 \us01/U104  ( .A(\us01/n81 ), .Y(\us01/n77 ) );
  AOI21X1 \us01/U103  ( .A0(\us01/n79 ), .A1(\us01/n80 ), .B0(\us01/n27 ), .Y(
        \us01/n78 ) );
  AOI211X1 \us01/U102  ( .A0(\us01/n5 ), .A1(\us01/n76 ), .B0(\us01/n77 ), 
        .C0(\us01/n78 ), .Y(\us01/n51 ) );
  OAI211X1 \us01/U101  ( .A0(\us01/n73 ), .A1(\us01/n27 ), .B0(\us01/n74 ), 
        .C0(\us01/n75 ), .Y(\us01/n72 ) );
  AOI21X1 \us01/U100  ( .A0(\us01/n68 ), .A1(\us01/n69 ), .B0(\us01/n6 ), .Y(
        \us01/n63 ) );
  INVX1 \us01/U99  ( .A(\us01/n67 ), .Y(\us01/n66 ) );
  OAI221XL \us01/U98  ( .A0(\us01/n63 ), .A1(\us01/n64 ), .B0(\us01/n65 ), 
        .B1(\us01/n27 ), .C0(\us01/n66 ), .Y(\us01/n56 ) );
  AOI2BB2X1 \us01/U97  ( .B0(\us01/n61 ), .B1(\us01/n24 ), .A0N(\us01/n62 ), 
        .A1N(\us01/n20 ), .Y(\us01/n60 ) );
  OAI221XL \us01/U96  ( .A0(\us01/n58 ), .A1(\us01/n18 ), .B0(\us01/n59 ), 
        .B1(\us01/n27 ), .C0(\us01/n60 ), .Y(\us01/n57 ) );
  AOI22X1 \us01/U95  ( .A0(\us01/n55 ), .A1(\us01/n56 ), .B0(\us01/n16 ), .B1(
        \us01/n57 ), .Y(\us01/n54 ) );
  OAI221XL \us01/U94  ( .A0(\us01/n51 ), .A1(\us01/n52 ), .B0(\us01/n53 ), 
        .B1(\us01/n10 ), .C0(\us01/n54 ), .Y(\us01/n7 ) );
  INVX1 \us01/U93  ( .A(\us01/n50 ), .Y(\us01/n49 ) );
  OAI221XL \us01/U92  ( .A0(\us01/n47 ), .A1(\us01/n18 ), .B0(\us01/n27 ), 
        .B1(\us01/n48 ), .C0(\us01/n49 ), .Y(\us01/n46 ) );
  NOR2X1 \us01/U91  ( .A(\us01/n41 ), .B(\us01/n42 ), .Y(\us01/n38 ) );
  INVX1 \us01/U90  ( .A(\us01/n40 ), .Y(\us01/n39 ) );
  INVX1 \us01/U89  ( .A(\us01/n32 ), .Y(\us01/n26 ) );
  AOI21X1 \us01/U88  ( .A0(\us01/n5 ), .A1(\us01/n30 ), .B0(\us01/n31 ), .Y(
        \us01/n29 ) );
  OAI221XL \us01/U87  ( .A0(\us01/n26 ), .A1(\us01/n27 ), .B0(\us01/n28 ), 
        .B1(\us01/n20 ), .C0(\us01/n29 ), .Y(\us01/n15 ) );
  OAI221XL \us01/U86  ( .A0(\us01/n18 ), .A1(\us01/n19 ), .B0(\us01/n20 ), 
        .B1(\us01/n21 ), .C0(\us01/n22 ), .Y(\us01/n17 ) );
  AOI22X1 \us01/U85  ( .A0(\us01/n14 ), .A1(\us01/n15 ), .B0(\us01/n16 ), .B1(
        \us01/n17 ), .Y(\us01/n13 ) );
  OAI221XL \us01/U84  ( .A0(\us01/n9 ), .A1(\us01/n10 ), .B0(\us01/n11 ), .B1(
        \us01/n12 ), .C0(\us01/n13 ), .Y(\us01/n8 ) );
  MX2X1 \us01/U83  ( .A(\us01/n7 ), .B(\us01/n8 ), .S0(sa01[6]), .Y(sa01_sr[7]) );
  NOR2X4 \us01/U82  ( .A(\us01/n129 ), .B(sa01[2]), .Y(\us01/n43 ) );
  CLKINVX3 \us01/U81  ( .A(\us01/n14 ), .Y(\us01/n52 ) );
  OAI22XL \us01/U80  ( .A0(\us01/n201 ), .A1(\us01/n52 ), .B0(\us01/n202 ), 
        .B1(\us01/n114 ), .Y(\us01/n193 ) );
  CLKINVX3 \us01/U79  ( .A(sa01[5]), .Y(\us01/n252 ) );
  NOR2X2 \us01/U78  ( .A(\us01/n252 ), .B(\us01/n234 ), .Y(\us01/n55 ) );
  CLKINVX3 \us01/U77  ( .A(sa01[7]), .Y(\us01/n129 ) );
  NOR2X4 \us01/U76  ( .A(\us01/n129 ), .B(\us01/n69 ), .Y(\us01/n24 ) );
  AOI22XL \us01/U75  ( .A0(\us01/n70 ), .A1(\us01/n24 ), .B0(\us01/n96 ), .B1(
        \us01/n129 ), .Y(\us01/n241 ) );
  NOR2X2 \us01/U74  ( .A(\us01/n252 ), .B(sa01[0]), .Y(\us01/n89 ) );
  CLKINVX3 \us01/U73  ( .A(sa01[0]), .Y(\us01/n234 ) );
  NOR2X4 \us01/U72  ( .A(\us01/n69 ), .B(sa01[7]), .Y(\us01/n33 ) );
  INVX12 \us01/U71  ( .A(\us01/n33 ), .Y(\us01/n27 ) );
  CLKINVX3 \us01/U70  ( .A(\us01/n1 ), .Y(\us01/n6 ) );
  CLKINVX3 \us01/U69  ( .A(\us01/n1 ), .Y(\us01/n5 ) );
  INVXL \us01/U68  ( .A(\us01/n24 ), .Y(\us01/n36 ) );
  INVX4 \us01/U67  ( .A(\us01/n3 ), .Y(\us01/n4 ) );
  INVXL \us01/U66  ( .A(\us01/n36 ), .Y(\us01/n3 ) );
  INVX4 \us01/U65  ( .A(sa01[1]), .Y(\us01/n226 ) );
  INVX4 \us01/U64  ( .A(\us01/n43 ), .Y(\us01/n20 ) );
  AOI221X4 \us01/U63  ( .A0(\us01/n24 ), .A1(\us01/n82 ), .B0(\us01/n43 ), 
        .B1(\us01/n295 ), .C0(\us01/n173 ), .Y(\us01/n346 ) );
  AOI221X4 \us01/U62  ( .A0(\us01/n5 ), .A1(\us01/n96 ), .B0(\us01/n43 ), .B1(
        \us01/n239 ), .C0(\us01/n340 ), .Y(\us01/n336 ) );
  AOI222X4 \us01/U61  ( .A0(\us01/n59 ), .A1(\us01/n43 ), .B0(\us01/n6 ), .B1(
        \us01/n221 ), .C0(\us01/n222 ), .C1(\us01/n187 ), .Y(\us01/n218 ) );
  AOI222X4 \us01/U60  ( .A0(\us01/n123 ), .A1(\us01/n43 ), .B0(sa01[2]), .B1(
        \us01/n203 ), .C0(\us01/n6 ), .C1(\us01/n71 ), .Y(\us01/n202 ) );
  AOI221X4 \us01/U59  ( .A0(\us01/n314 ), .A1(\us01/n43 ), .B0(\us01/n160 ), 
        .B1(\us01/n24 ), .C0(\us01/n315 ), .Y(\us01/n307 ) );
  AOI221X4 \us01/U58  ( .A0(\us01/n43 ), .A1(\us01/n208 ), .B0(\us01/n76 ), 
        .B1(\us01/n24 ), .C0(\us01/n209 ), .Y(\us01/n207 ) );
  AOI221X4 \us01/U57  ( .A0(\us01/n43 ), .A1(\us01/n205 ), .B0(\us01/n32 ), 
        .B1(\us01/n6 ), .C0(\us01/n206 ), .Y(\us01/n201 ) );
  AOI221X4 \us01/U56  ( .A0(\us01/n43 ), .A1(\us01/n44 ), .B0(\us01/n45 ), 
        .B1(\us01/n24 ), .C0(\us01/n46 ), .Y(\us01/n9 ) );
  AOI22XL \us01/U55  ( .A0(\us01/n217 ), .A1(\us01/n43 ), .B0(\us01/n33 ), 
        .B1(\us01/n47 ), .Y(\us01/n216 ) );
  AOI22XL \us01/U54  ( .A0(\us01/n98 ), .A1(\us01/n43 ), .B0(\us01/n6 ), .B1(
        \us01/n99 ), .Y(\us01/n97 ) );
  AOI22XL \us01/U53  ( .A0(\us01/n82 ), .A1(\us01/n43 ), .B0(\us01/n83 ), .B1(
        \us01/n24 ), .Y(\us01/n81 ) );
  AOI2BB2XL \us01/U52  ( .B0(\us01/n43 ), .B1(\us01/n94 ), .A0N(\us01/n120 ), 
        .A1N(\us01/n4 ), .Y(\us01/n119 ) );
  AOI222X4 \us01/U51  ( .A0(\us01/n125 ), .A1(\us01/n33 ), .B0(\us01/n145 ), 
        .B1(\us01/n40 ), .C0(\us01/n43 ), .C1(\us01/n184 ), .Y(\us01/n183 ) );
  AOI22XL \us01/U50  ( .A0(\us01/n43 ), .A1(\us01/n303 ), .B0(\us01/n24 ), 
        .B1(\us01/n96 ), .Y(\us01/n358 ) );
  AOI22XL \us01/U49  ( .A0(\us01/n43 ), .A1(\us01/n100 ), .B0(\us01/n24 ), 
        .B1(\us01/n125 ), .Y(\us01/n124 ) );
  AOI21XL \us01/U48  ( .A0(\us01/n159 ), .A1(\us01/n43 ), .B0(\us01/n40 ), .Y(
        \us01/n262 ) );
  AOI22XL \us01/U47  ( .A0(\us01/n40 ), .A1(\us01/n94 ), .B0(\us01/n43 ), .B1(
        \us01/n187 ), .Y(\us01/n244 ) );
  AOI22XL \us01/U46  ( .A0(\us01/n184 ), .A1(\us01/n5 ), .B0(\us01/n198 ), 
        .B1(\us01/n43 ), .Y(\us01/n197 ) );
  NOR2XL \us01/U45  ( .A(\us01/n33 ), .B(\us01/n2 ), .Y(\us01/n302 ) );
  MXI2XL \us01/U44  ( .A(\us01/n2 ), .B(\us01/n6 ), .S0(\us01/n28 ), .Y(
        \us01/n311 ) );
  INVXL \us01/U43  ( .A(\us01/n20 ), .Y(\us01/n2 ) );
  INVX4 \us01/U42  ( .A(\us01/n6 ), .Y(\us01/n18 ) );
  AOI21XL \us01/U41  ( .A0(\us01/n18 ), .A1(\us01/n162 ), .B0(\us01/n25 ), .Y(
        \us01/n161 ) );
  INVX4 \us01/U40  ( .A(sa01[2]), .Y(\us01/n69 ) );
  NOR2X4 \us01/U39  ( .A(\us01/n226 ), .B(\us01/n4 ), .Y(\us01/n40 ) );
  CLKINVX3 \us01/U38  ( .A(sa01[3]), .Y(\us01/n136 ) );
  NOR2X2 \us01/U37  ( .A(\us01/n136 ), .B(sa01[4]), .Y(\us01/n145 ) );
  CLKINVX3 \us01/U36  ( .A(sa01[4]), .Y(\us01/n58 ) );
  NOR2X2 \us01/U35  ( .A(\us01/n58 ), .B(sa01[3]), .Y(\us01/n159 ) );
  NOR2X2 \us01/U34  ( .A(\us01/n136 ), .B(\us01/n58 ), .Y(\us01/n259 ) );
  NOR2X2 \us01/U33  ( .A(sa01[4]), .B(sa01[3]), .Y(\us01/n278 ) );
  NOR2X2 \us01/U32  ( .A(\us01/n259 ), .B(\us01/n278 ), .Y(\us01/n47 ) );
  CLKINVX3 \us01/U31  ( .A(\us01/n259 ), .Y(\us01/n44 ) );
  NOR2X2 \us01/U30  ( .A(\us01/n44 ), .B(sa01[1]), .Y(\us01/n137 ) );
  AOI21XL \us01/U29  ( .A0(\us01/n44 ), .A1(\us01/n111 ), .B0(\us01/n4 ), .Y(
        \us01/n177 ) );
  AOI22XL \us01/U28  ( .A0(\us01/n23 ), .A1(\us01/n24 ), .B0(\us01/n25 ), .B1(
        sa01[2]), .Y(\us01/n22 ) );
  AOI22XL \us01/U27  ( .A0(\us01/n33 ), .A1(sa01[3]), .B0(\us01/n24 ), .B1(
        \us01/n58 ), .Y(\us01/n277 ) );
  NAND2XL \us01/U26  ( .A(\us01/n198 ), .B(\us01/n24 ), .Y(\us01/n132 ) );
  OAI2BB2XL \us01/U25  ( .B0(\us01/n20 ), .B1(\us01/n111 ), .A0N(\us01/n125 ), 
        .A1N(\us01/n24 ), .Y(\us01/n220 ) );
  NAND2XL \us01/U24  ( .A(\us01/n111 ), .B(\us01/n101 ), .Y(\us01/n21 ) );
  NAND2XL \us01/U23  ( .A(\us01/n111 ), .B(\us01/n300 ), .Y(\us01/n187 ) );
  NAND2XL \us01/U22  ( .A(\us01/n111 ), .B(\us01/n121 ), .Y(\us01/n303 ) );
  AOI221XL \us01/U21  ( .A0(\us01/n43 ), .A1(\us01/n151 ), .B0(\us01/n25 ), 
        .B1(\us01/n69 ), .C0(\us01/n275 ), .Y(\us01/n274 ) );
  NOR2BXL \us01/U20  ( .AN(\us01/n101 ), .B(\us01/n25 ), .Y(\us01/n172 ) );
  NAND2X2 \us01/U19  ( .A(\us01/n58 ), .B(\us01/n226 ), .Y(\us01/n34 ) );
  OAI222X1 \us01/U18  ( .A0(\us01/n27 ), .A1(\us01/n34 ), .B0(\us01/n69 ), 
        .B1(\us01/n205 ), .C0(\us01/n20 ), .C1(\us01/n79 ), .Y(\us01/n260 ) );
  OAI222X1 \us01/U17  ( .A0(\us01/n20 ), .A1(\us01/n99 ), .B0(\us01/n27 ), 
        .B1(\us01/n101 ), .C0(\us01/n184 ), .C1(\us01/n4 ), .Y(\us01/n250 ) );
  OAI222X1 \us01/U16  ( .A0(\us01/n4 ), .A1(\us01/n37 ), .B0(\us01/n38 ), .B1(
        \us01/n20 ), .C0(sa01[4]), .C1(\us01/n39 ), .Y(\us01/n35 ) );
  AOI221X1 \us01/U15  ( .A0(\us01/n5 ), .A1(\us01/n19 ), .B0(\us01/n33 ), .B1(
        \us01/n34 ), .C0(\us01/n35 ), .Y(\us01/n11 ) );
  OR2X2 \us01/U14  ( .A(sa01[2]), .B(sa01[7]), .Y(\us01/n1 ) );
  AOI221XL \us01/U13  ( .A0(\us01/n70 ), .A1(\us01/n43 ), .B0(\us01/n24 ), 
        .B1(\us01/n71 ), .C0(\us01/n72 ), .Y(\us01/n53 ) );
  AOI221XL \us01/U12  ( .A0(\us01/n59 ), .A1(\us01/n33 ), .B0(\us01/n43 ), 
        .B1(\us01/n126 ), .C0(\us01/n127 ), .Y(\us01/n113 ) );
  AOI222XL \us01/U11  ( .A0(\us01/n185 ), .A1(\us01/n43 ), .B0(\us01/n186 ), 
        .B1(\us01/n187 ), .C0(\us01/n6 ), .C1(\us01/n188 ), .Y(\us01/n164 ) );
  AOI221X1 \us01/U10  ( .A0(\us01/n313 ), .A1(\us01/n5 ), .B0(\us01/n23 ), 
        .B1(\us01/n2 ), .C0(\us01/n328 ), .Y(\us01/n320 ) );
  AOI221X1 \us01/U9  ( .A0(\us01/n40 ), .A1(\us01/n136 ), .B0(\us01/n33 ), 
        .B1(\us01/n178 ), .C0(\us01/n338 ), .Y(\us01/n337 ) );
  AOI222XL \us01/U8  ( .A0(\us01/n278 ), .A1(\us01/n24 ), .B0(\us01/n42 ), 
        .B1(\us01/n33 ), .C0(\us01/n43 ), .C1(\us01/n136 ), .Y(\us01/n351 ) );
  AOI31X1 \us01/U7  ( .A0(sa01[2]), .A1(\us01/n58 ), .A2(sa01[1]), .B0(
        \us01/n40 ), .Y(\us01/n350 ) );
  AOI31X1 \us01/U6  ( .A0(\us01/n44 ), .A1(\us01/n129 ), .A2(\us01/n130 ), 
        .B0(\us01/n131 ), .Y(\us01/n128 ) );
  AOI221X1 \us01/U5  ( .A0(\us01/n40 ), .A1(\us01/n136 ), .B0(\us01/n33 ), 
        .B1(\us01/n47 ), .C0(\us01/n156 ), .Y(\us01/n141 ) );
  OAI32X1 \us01/U4  ( .A0(\us01/n210 ), .A1(\us01/n145 ), .A2(\us01/n18 ), 
        .B0(\us01/n27 ), .B1(\us01/n211 ), .Y(\us01/n209 ) );
  AOI221X1 \us01/U3  ( .A0(\us01/n278 ), .A1(\us01/n40 ), .B0(\us01/n185 ), 
        .B1(\us01/n2 ), .C0(\us01/n279 ), .Y(\us01/n273 ) );
  OAI32X1 \us01/U2  ( .A0(\us01/n18 ), .A1(sa01[1]), .A2(\us01/n159 ), .B0(
        sa01[4]), .B1(\us01/n182 ), .Y(\us01/n318 ) );
  AOI31XL \us01/U1  ( .A0(\us01/n79 ), .A1(\us01/n44 ), .A2(\us01/n2 ), .B0(
        \us01/n280 ), .Y(\us01/n339 ) );
  NAND2X1 \us02/U366  ( .A(\us02/n47 ), .B(\us02/n226 ), .Y(\us02/n189 ) );
  NOR2X1 \us02/U365  ( .A(\us02/n226 ), .B(sa02[3]), .Y(\us02/n242 ) );
  INVX1 \us02/U364  ( .A(\us02/n242 ), .Y(\us02/n205 ) );
  AND2X1 \us02/U363  ( .A(\us02/n189 ), .B(\us02/n205 ), .Y(\us02/n65 ) );
  NOR2X1 \us02/U362  ( .A(\us02/n226 ), .B(\us02/n47 ), .Y(\us02/n45 ) );
  NOR2X1 \us02/U361  ( .A(\us02/n259 ), .B(\us02/n45 ), .Y(\us02/n73 ) );
  NAND2BX1 \us02/U360  ( .AN(\us02/n73 ), .B(\us02/n6 ), .Y(\us02/n158 ) );
  NOR2X1 \us02/U359  ( .A(\us02/n226 ), .B(\us02/n159 ), .Y(\us02/n95 ) );
  INVX1 \us02/U358  ( .A(\us02/n95 ), .Y(\us02/n111 ) );
  NOR2X1 \us02/U357  ( .A(\us02/n145 ), .B(sa02[1]), .Y(\us02/n42 ) );
  INVX1 \us02/U356  ( .A(\us02/n42 ), .Y(\us02/n121 ) );
  INVX1 \us02/U355  ( .A(\us02/n47 ), .Y(\us02/n96 ) );
  OAI211X1 \us02/U354  ( .A0(\us02/n65 ), .A1(\us02/n27 ), .B0(\us02/n158 ), 
        .C0(\us02/n358 ), .Y(\us02/n355 ) );
  NOR2X1 \us02/U353  ( .A(\us02/n226 ), .B(\us02/n145 ), .Y(\us02/n59 ) );
  NOR2X1 \us02/U352  ( .A(\us02/n96 ), .B(\us02/n59 ), .Y(\us02/n271 ) );
  NOR2X1 \us02/U351  ( .A(\us02/n226 ), .B(\us02/n278 ), .Y(\us02/n217 ) );
  INVX1 \us02/U350  ( .A(\us02/n217 ), .Y(\us02/n150 ) );
  NAND2X1 \us02/U349  ( .A(\us02/n44 ), .B(\us02/n150 ), .Y(\us02/n147 ) );
  NAND2X1 \us02/U348  ( .A(sa02[4]), .B(\us02/n226 ), .Y(\us02/n101 ) );
  INVX1 \us02/U347  ( .A(\us02/n159 ), .Y(\us02/n188 ) );
  NOR2X1 \us02/U346  ( .A(\us02/n188 ), .B(\us02/n226 ), .Y(\us02/n25 ) );
  INVX1 \us02/U345  ( .A(\us02/n172 ), .Y(\us02/n107 ) );
  AOI22X1 \us02/U344  ( .A0(\us02/n33 ), .A1(\us02/n147 ), .B0(\us02/n24 ), 
        .B1(\us02/n107 ), .Y(\us02/n357 ) );
  OAI221XL \us02/U343  ( .A0(\us02/n18 ), .A1(\us02/n121 ), .B0(\us02/n271 ), 
        .B1(\us02/n20 ), .C0(\us02/n357 ), .Y(\us02/n356 ) );
  MXI2X1 \us02/U342  ( .A(\us02/n355 ), .B(\us02/n356 ), .S0(\us02/n252 ), .Y(
        \us02/n331 ) );
  INVX1 \us02/U341  ( .A(\us02/n59 ), .Y(\us02/n79 ) );
  AND2X1 \us02/U340  ( .A(\us02/n101 ), .B(\us02/n79 ), .Y(\us02/n325 ) );
  XNOR2X1 \us02/U339  ( .A(sa02[5]), .B(\us02/n226 ), .Y(\us02/n352 ) );
  NOR2X1 \us02/U338  ( .A(\us02/n226 ), .B(\us02/n136 ), .Y(\us02/n281 ) );
  INVX1 \us02/U337  ( .A(\us02/n281 ), .Y(\us02/n19 ) );
  NAND2X1 \us02/U336  ( .A(\us02/n145 ), .B(\us02/n226 ), .Y(\us02/n223 ) );
  AOI21X1 \us02/U335  ( .A0(\us02/n19 ), .A1(\us02/n223 ), .B0(\us02/n27 ), 
        .Y(\us02/n354 ) );
  AOI31X1 \us02/U334  ( .A0(\us02/n6 ), .A1(\us02/n352 ), .A2(\us02/n259 ), 
        .B0(\us02/n354 ), .Y(\us02/n353 ) );
  OAI221XL \us02/U333  ( .A0(\us02/n20 ), .A1(\us02/n34 ), .B0(\us02/n325 ), 
        .B1(\us02/n4 ), .C0(\us02/n353 ), .Y(\us02/n347 ) );
  INVX1 \us02/U332  ( .A(\us02/n352 ), .Y(\us02/n349 ) );
  NAND2X1 \us02/U331  ( .A(\us02/n278 ), .B(\us02/n6 ), .Y(\us02/n74 ) );
  OAI211X1 \us02/U330  ( .A0(\us02/n349 ), .A1(\us02/n74 ), .B0(\us02/n350 ), 
        .C0(\us02/n351 ), .Y(\us02/n348 ) );
  MXI2X1 \us02/U329  ( .A(\us02/n347 ), .B(\us02/n348 ), .S0(\us02/n252 ), .Y(
        \us02/n332 ) );
  NOR2X1 \us02/U328  ( .A(\us02/n44 ), .B(\us02/n226 ), .Y(\us02/n157 ) );
  INVX1 \us02/U327  ( .A(\us02/n157 ), .Y(\us02/n240 ) );
  NAND2X1 \us02/U326  ( .A(\us02/n240 ), .B(\us02/n189 ), .Y(\us02/n68 ) );
  NOR2X1 \us02/U325  ( .A(\us02/n20 ), .B(\us02/n159 ), .Y(\us02/n225 ) );
  NOR2X1 \us02/U324  ( .A(\us02/n225 ), .B(\us02/n40 ), .Y(\us02/n345 ) );
  INVX1 \us02/U323  ( .A(\us02/n278 ), .Y(\us02/n94 ) );
  NAND2X1 \us02/U322  ( .A(\us02/n94 ), .B(\us02/n226 ), .Y(\us02/n199 ) );
  NAND2X1 \us02/U321  ( .A(\us02/n199 ), .B(\us02/n205 ), .Y(\us02/n82 ) );
  NAND2X1 \us02/U320  ( .A(\us02/n19 ), .B(\us02/n199 ), .Y(\us02/n295 ) );
  NOR2X1 \us02/U319  ( .A(\us02/n226 ), .B(\us02/n259 ), .Y(\us02/n210 ) );
  NOR2X1 \us02/U318  ( .A(\us02/n27 ), .B(\us02/n210 ), .Y(\us02/n173 ) );
  MXI2X1 \us02/U317  ( .A(\us02/n345 ), .B(\us02/n346 ), .S0(\us02/n252 ), .Y(
        \us02/n342 ) );
  NOR2X1 \us02/U316  ( .A(sa02[1]), .B(sa02[3]), .Y(\us02/n163 ) );
  INVX1 \us02/U315  ( .A(\us02/n163 ), .Y(\us02/n37 ) );
  INVX1 \us02/U314  ( .A(\us02/n173 ), .Y(\us02/n344 ) );
  AOI21X1 \us02/U313  ( .A0(\us02/n240 ), .A1(\us02/n37 ), .B0(\us02/n344 ), 
        .Y(\us02/n343 ) );
  AOI211X1 \us02/U312  ( .A0(\us02/n5 ), .A1(\us02/n68 ), .B0(\us02/n342 ), 
        .C0(\us02/n343 ), .Y(\us02/n333 ) );
  NOR2X1 \us02/U311  ( .A(\us02/n18 ), .B(\us02/n226 ), .Y(\us02/n258 ) );
  NAND2X1 \us02/U310  ( .A(\us02/n278 ), .B(sa02[1]), .Y(\us02/n204 ) );
  NOR2X1 \us02/U309  ( .A(\us02/n188 ), .B(sa02[1]), .Y(\us02/n179 ) );
  INVX1 \us02/U308  ( .A(\us02/n179 ), .Y(\us02/n330 ) );
  NAND2X1 \us02/U307  ( .A(\us02/n204 ), .B(\us02/n330 ), .Y(\us02/n239 ) );
  NOR2X1 \us02/U306  ( .A(\us02/n136 ), .B(sa02[1]), .Y(\us02/n299 ) );
  NOR2X1 \us02/U305  ( .A(\us02/n299 ), .B(\us02/n210 ), .Y(\us02/n341 ) );
  OAI32X1 \us02/U304  ( .A0(\us02/n27 ), .A1(\us02/n278 ), .A2(\us02/n95 ), 
        .B0(\us02/n341 ), .B1(\us02/n4 ), .Y(\us02/n340 ) );
  INVX1 \us02/U303  ( .A(\us02/n45 ), .Y(\us02/n126 ) );
  NAND2X1 \us02/U302  ( .A(\us02/n126 ), .B(\us02/n101 ), .Y(\us02/n178 ) );
  NOR2X1 \us02/U301  ( .A(\us02/n18 ), .B(\us02/n136 ), .Y(\us02/n280 ) );
  OAI21XL \us02/U300  ( .A0(\us02/n4 ), .A1(\us02/n121 ), .B0(\us02/n339 ), 
        .Y(\us02/n338 ) );
  MXI2X1 \us02/U299  ( .A(\us02/n336 ), .B(\us02/n337 ), .S0(\us02/n252 ), .Y(
        \us02/n335 ) );
  NOR2X1 \us02/U298  ( .A(\us02/n258 ), .B(\us02/n335 ), .Y(\us02/n334 ) );
  MX4X1 \us02/U297  ( .A(\us02/n331 ), .B(\us02/n332 ), .C(\us02/n333 ), .D(
        \us02/n334 ), .S0(sa02[6]), .S1(\us02/n234 ), .Y(sa02_sr[0]) );
  INVX1 \us02/U296  ( .A(\us02/n299 ), .Y(\us02/n80 ) );
  NOR2X1 \us02/U295  ( .A(\us02/n111 ), .B(\us02/n18 ), .Y(\us02/n269 ) );
  INVX1 \us02/U294  ( .A(\us02/n269 ), .Y(\us02/n75 ) );
  OAI221XL \us02/U293  ( .A0(\us02/n18 ), .A1(\us02/n330 ), .B0(\us02/n20 ), 
        .B1(\us02/n80 ), .C0(\us02/n75 ), .Y(\us02/n329 ) );
  AOI221X1 \us02/U292  ( .A0(\us02/n325 ), .A1(\us02/n33 ), .B0(\us02/n24 ), 
        .B1(\us02/n303 ), .C0(\us02/n329 ), .Y(\us02/n319 ) );
  NOR2X1 \us02/U291  ( .A(\us02/n234 ), .B(sa02[5]), .Y(\us02/n14 ) );
  NOR2X1 \us02/U290  ( .A(\us02/n25 ), .B(\us02/n299 ), .Y(\us02/n313 ) );
  NAND2X1 \us02/U289  ( .A(\us02/n44 ), .B(\us02/n226 ), .Y(\us02/n300 ) );
  AND2X1 \us02/U288  ( .A(\us02/n300 ), .B(\us02/n240 ), .Y(\us02/n23 ) );
  OAI32X1 \us02/U287  ( .A0(\us02/n4 ), .A1(\us02/n145 ), .A2(\us02/n210 ), 
        .B0(\us02/n137 ), .B1(\us02/n27 ), .Y(\us02/n328 ) );
  NOR2X1 \us02/U286  ( .A(sa02[0]), .B(sa02[5]), .Y(\us02/n16 ) );
  INVX1 \us02/U285  ( .A(\us02/n16 ), .Y(\us02/n114 ) );
  INVX1 \us02/U284  ( .A(\us02/n145 ), .Y(\us02/n149 ) );
  NOR2X1 \us02/U283  ( .A(\us02/n47 ), .B(sa02[1]), .Y(\us02/n98 ) );
  INVX1 \us02/U282  ( .A(\us02/n98 ), .Y(\us02/n284 ) );
  OAI21XL \us02/U281  ( .A0(\us02/n69 ), .A1(\us02/n284 ), .B0(\us02/n27 ), 
        .Y(\us02/n327 ) );
  AOI31X1 \us02/U280  ( .A0(\us02/n111 ), .A1(\us02/n149 ), .A2(\us02/n327 ), 
        .B0(\us02/n225 ), .Y(\us02/n326 ) );
  OAI21XL \us02/U279  ( .A0(\us02/n325 ), .A1(\us02/n18 ), .B0(\us02/n326 ), 
        .Y(\us02/n322 ) );
  NAND2X1 \us02/U278  ( .A(\us02/n19 ), .B(\us02/n189 ), .Y(\us02/n71 ) );
  NOR2X1 \us02/U277  ( .A(\us02/n71 ), .B(\us02/n18 ), .Y(\us02/n135 ) );
  AOI21X1 \us02/U276  ( .A0(\us02/n40 ), .A1(sa02[4]), .B0(\us02/n135 ), .Y(
        \us02/n324 ) );
  OAI221XL \us02/U275  ( .A0(\us02/n47 ), .A1(\us02/n27 ), .B0(\us02/n65 ), 
        .B1(\us02/n20 ), .C0(\us02/n324 ), .Y(\us02/n323 ) );
  AOI22X1 \us02/U274  ( .A0(\us02/n55 ), .A1(\us02/n322 ), .B0(\us02/n89 ), 
        .B1(\us02/n323 ), .Y(\us02/n321 ) );
  OAI221XL \us02/U273  ( .A0(\us02/n319 ), .A1(\us02/n52 ), .B0(\us02/n320 ), 
        .B1(\us02/n114 ), .C0(\us02/n321 ), .Y(\us02/n304 ) );
  NOR2X1 \us02/U272  ( .A(\us02/n226 ), .B(\us02/n58 ), .Y(\us02/n290 ) );
  INVX1 \us02/U271  ( .A(\us02/n290 ), .Y(\us02/n200 ) );
  NAND2X1 \us02/U270  ( .A(\us02/n34 ), .B(\us02/n200 ), .Y(\us02/n120 ) );
  INVX1 \us02/U269  ( .A(\us02/n210 ), .Y(\us02/n100 ) );
  OAI221XL \us02/U268  ( .A0(\us02/n20 ), .A1(\us02/n100 ), .B0(sa02[3]), .B1(
        \us02/n4 ), .C0(\us02/n262 ), .Y(\us02/n317 ) );
  INVX1 \us02/U267  ( .A(\us02/n258 ), .Y(\us02/n182 ) );
  AOI211X1 \us02/U266  ( .A0(\us02/n33 ), .A1(\us02/n120 ), .B0(\us02/n317 ), 
        .C0(\us02/n318 ), .Y(\us02/n306 ) );
  NAND2X1 \us02/U265  ( .A(\us02/n100 ), .B(\us02/n199 ), .Y(\us02/n151 ) );
  INVX1 \us02/U264  ( .A(\us02/n151 ), .Y(\us02/n314 ) );
  NOR2X1 \us02/U263  ( .A(\us02/n45 ), .B(\us02/n163 ), .Y(\us02/n160 ) );
  INVX1 \us02/U262  ( .A(\us02/n295 ), .Y(\us02/n92 ) );
  AOI21X1 \us02/U261  ( .A0(sa02[1]), .A1(\us02/n58 ), .B0(\us02/n98 ), .Y(
        \us02/n316 ) );
  OAI22X1 \us02/U260  ( .A0(\us02/n92 ), .A1(\us02/n18 ), .B0(\us02/n316 ), 
        .B1(\us02/n27 ), .Y(\us02/n315 ) );
  NOR2X1 \us02/U259  ( .A(\us02/n149 ), .B(\us02/n226 ), .Y(\us02/n41 ) );
  INVX1 \us02/U258  ( .A(\us02/n41 ), .Y(\us02/n105 ) );
  NAND2X1 \us02/U257  ( .A(\us02/n284 ), .B(\us02/n105 ), .Y(\us02/n227 ) );
  AOI21X1 \us02/U256  ( .A0(\us02/n313 ), .A1(\us02/n33 ), .B0(\us02/n269 ), 
        .Y(\us02/n312 ) );
  OAI221XL \us02/U255  ( .A0(\us02/n149 ), .A1(\us02/n20 ), .B0(\us02/n4 ), 
        .B1(\us02/n227 ), .C0(\us02/n312 ), .Y(\us02/n309 ) );
  AOI21X1 \us02/U254  ( .A0(\us02/n226 ), .A1(\us02/n188 ), .B0(\us02/n242 ), 
        .Y(\us02/n185 ) );
  INVX1 \us02/U253  ( .A(\us02/n185 ), .Y(\us02/n48 ) );
  AND2X1 \us02/U252  ( .A(\us02/n223 ), .B(\us02/n240 ), .Y(\us02/n28 ) );
  OAI221XL \us02/U251  ( .A0(\us02/n27 ), .A1(\us02/n44 ), .B0(\us02/n4 ), 
        .B1(\us02/n48 ), .C0(\us02/n311 ), .Y(\us02/n310 ) );
  AOI22X1 \us02/U250  ( .A0(\us02/n89 ), .A1(\us02/n309 ), .B0(\us02/n55 ), 
        .B1(\us02/n310 ), .Y(\us02/n308 ) );
  OAI221XL \us02/U249  ( .A0(\us02/n306 ), .A1(\us02/n52 ), .B0(\us02/n307 ), 
        .B1(\us02/n114 ), .C0(\us02/n308 ), .Y(\us02/n305 ) );
  MX2X1 \us02/U248  ( .A(\us02/n304 ), .B(\us02/n305 ), .S0(sa02[6]), .Y(
        sa02_sr[1]) );
  INVX1 \us02/U247  ( .A(\us02/n187 ), .Y(\us02/n61 ) );
  MXI2X1 \us02/U246  ( .A(\us02/n303 ), .B(\us02/n61 ), .S0(\us02/n69 ), .Y(
        \us02/n301 ) );
  MXI2X1 \us02/U245  ( .A(\us02/n301 ), .B(\us02/n147 ), .S0(\us02/n302 ), .Y(
        \us02/n285 ) );
  NAND2X1 \us02/U244  ( .A(\us02/n200 ), .B(\us02/n300 ), .Y(\us02/n99 ) );
  INVX1 \us02/U243  ( .A(\us02/n99 ), .Y(\us02/n296 ) );
  NOR2X1 \us02/U242  ( .A(\us02/n299 ), .B(\us02/n242 ), .Y(\us02/n298 ) );
  NAND2X1 \us02/U241  ( .A(sa02[1]), .B(\us02/n47 ), .Y(\us02/n122 ) );
  NOR2X1 \us02/U240  ( .A(\us02/n159 ), .B(\us02/n217 ), .Y(\us02/n198 ) );
  OAI221XL \us02/U239  ( .A0(\us02/n298 ), .A1(\us02/n27 ), .B0(\us02/n20 ), 
        .B1(\us02/n122 ), .C0(\us02/n132 ), .Y(\us02/n297 ) );
  AOI221X1 \us02/U238  ( .A0(\us02/n225 ), .A1(\us02/n226 ), .B0(\us02/n296 ), 
        .B1(\us02/n6 ), .C0(\us02/n297 ), .Y(\us02/n291 ) );
  OAI2BB2X1 \us02/U237  ( .B0(\us02/n27 ), .B1(\us02/n295 ), .A0N(\us02/n34 ), 
        .A1N(\us02/n24 ), .Y(\us02/n293 ) );
  AOI21X1 \us02/U236  ( .A0(\us02/n101 ), .A1(\us02/n150 ), .B0(\us02/n20 ), 
        .Y(\us02/n294 ) );
  AOI211X1 \us02/U235  ( .A0(\us02/n5 ), .A1(\us02/n79 ), .B0(\us02/n293 ), 
        .C0(\us02/n294 ), .Y(\us02/n292 ) );
  INVX1 \us02/U234  ( .A(\us02/n89 ), .Y(\us02/n10 ) );
  OAI22X1 \us02/U233  ( .A0(\us02/n291 ), .A1(\us02/n114 ), .B0(\us02/n292 ), 
        .B1(\us02/n10 ), .Y(\us02/n286 ) );
  INVX1 \us02/U232  ( .A(\us02/n225 ), .Y(\us02/n288 ) );
  NAND2X1 \us02/U231  ( .A(\us02/n200 ), .B(\us02/n284 ), .Y(\us02/n102 ) );
  NOR2X1 \us02/U230  ( .A(\us02/n290 ), .B(\us02/n163 ), .Y(\us02/n184 ) );
  AOI22X1 \us02/U229  ( .A0(\us02/n102 ), .A1(\us02/n69 ), .B0(\us02/n184 ), 
        .B1(\us02/n33 ), .Y(\us02/n289 ) );
  AOI31X1 \us02/U228  ( .A0(\us02/n132 ), .A1(\us02/n288 ), .A2(\us02/n289 ), 
        .B0(\us02/n52 ), .Y(\us02/n287 ) );
  AOI211X1 \us02/U227  ( .A0(\us02/n285 ), .A1(\us02/n55 ), .B0(\us02/n286 ), 
        .C0(\us02/n287 ), .Y(\us02/n263 ) );
  NAND2X1 \us02/U226  ( .A(\us02/n284 ), .B(\us02/n122 ), .Y(\us02/n125 ) );
  NOR2X1 \us02/U225  ( .A(\us02/n199 ), .B(\us02/n4 ), .Y(\us02/n50 ) );
  AOI21X1 \us02/U224  ( .A0(\us02/n200 ), .A1(\us02/n223 ), .B0(\us02/n20 ), 
        .Y(\us02/n283 ) );
  AOI211X1 \us02/U223  ( .A0(\us02/n5 ), .A1(\us02/n125 ), .B0(\us02/n50 ), 
        .C0(\us02/n283 ), .Y(\us02/n282 ) );
  OAI221XL \us02/U222  ( .A0(\us02/n281 ), .A1(\us02/n27 ), .B0(\us02/n4 ), 
        .B1(\us02/n111 ), .C0(\us02/n282 ), .Y(\us02/n265 ) );
  INVX1 \us02/U221  ( .A(\us02/n280 ), .Y(\us02/n247 ) );
  NAND2X1 \us02/U220  ( .A(\us02/n41 ), .B(\us02/n33 ), .Y(\us02/n272 ) );
  OAI221XL \us02/U219  ( .A0(sa02[1]), .A1(\us02/n247 ), .B0(\us02/n4 ), .B1(
        \us02/n189 ), .C0(\us02/n272 ), .Y(\us02/n279 ) );
  NAND2X1 \us02/U218  ( .A(sa02[2]), .B(\us02/n149 ), .Y(\us02/n276 ) );
  XNOR2X1 \us02/U217  ( .A(\us02/n129 ), .B(sa02[1]), .Y(\us02/n155 ) );
  MXI2X1 \us02/U216  ( .A(\us02/n276 ), .B(\us02/n277 ), .S0(\us02/n155 ), .Y(
        \us02/n275 ) );
  OAI22X1 \us02/U215  ( .A0(\us02/n273 ), .A1(\us02/n10 ), .B0(\us02/n274 ), 
        .B1(\us02/n52 ), .Y(\us02/n266 ) );
  NOR2X1 \us02/U214  ( .A(\us02/n20 ), .B(\us02/n226 ), .Y(\us02/n176 ) );
  OAI21XL \us02/U213  ( .A0(\us02/n4 ), .A1(\us02/n271 ), .B0(\us02/n272 ), 
        .Y(\us02/n270 ) );
  OAI31X1 \us02/U212  ( .A0(\us02/n176 ), .A1(\us02/n269 ), .A2(\us02/n270 ), 
        .B0(\us02/n16 ), .Y(\us02/n268 ) );
  INVX1 \us02/U211  ( .A(\us02/n268 ), .Y(\us02/n267 ) );
  AOI211X1 \us02/U210  ( .A0(\us02/n55 ), .A1(\us02/n265 ), .B0(\us02/n266 ), 
        .C0(\us02/n267 ), .Y(\us02/n264 ) );
  MXI2X1 \us02/U209  ( .A(\us02/n263 ), .B(\us02/n264 ), .S0(sa02[6]), .Y(
        sa02_sr[2]) );
  NOR2X1 \us02/U208  ( .A(\us02/n94 ), .B(sa02[1]), .Y(\us02/n211 ) );
  INVX1 \us02/U207  ( .A(\us02/n262 ), .Y(\us02/n261 ) );
  AOI211X1 \us02/U206  ( .A0(\us02/n259 ), .A1(\us02/n24 ), .B0(\us02/n260 ), 
        .C0(\us02/n261 ), .Y(\us02/n255 ) );
  OAI22X1 \us02/U205  ( .A0(\us02/n20 ), .A1(\us02/n68 ), .B0(\us02/n27 ), 
        .B1(\us02/n37 ), .Y(\us02/n257 ) );
  NOR3X1 \us02/U204  ( .A(\us02/n257 ), .B(\us02/n258 ), .C(\us02/n50 ), .Y(
        \us02/n256 ) );
  MXI2X1 \us02/U203  ( .A(\us02/n255 ), .B(\us02/n256 ), .S0(\us02/n252 ), .Y(
        \us02/n254 ) );
  AOI221X1 \us02/U202  ( .A0(\us02/n211 ), .A1(\us02/n5 ), .B0(\us02/n40 ), 
        .B1(sa02[4]), .C0(\us02/n254 ), .Y(\us02/n248 ) );
  INVX1 \us02/U201  ( .A(\us02/n211 ), .Y(\us02/n106 ) );
  NAND2X1 \us02/U200  ( .A(\us02/n200 ), .B(\us02/n106 ), .Y(\us02/n83 ) );
  NAND2X1 \us02/U199  ( .A(\us02/n199 ), .B(\us02/n204 ), .Y(\us02/n169 ) );
  AOI2BB2X1 \us02/U198  ( .B0(\us02/n65 ), .B1(\us02/n24 ), .A0N(\us02/n169 ), 
        .A1N(\us02/n20 ), .Y(\us02/n253 ) );
  OAI221XL \us02/U197  ( .A0(\us02/n172 ), .A1(\us02/n18 ), .B0(\us02/n27 ), 
        .B1(\us02/n83 ), .C0(\us02/n253 ), .Y(\us02/n251 ) );
  MXI2X1 \us02/U196  ( .A(\us02/n250 ), .B(\us02/n251 ), .S0(\us02/n252 ), .Y(
        \us02/n249 ) );
  MXI2X1 \us02/U195  ( .A(\us02/n248 ), .B(\us02/n249 ), .S0(\us02/n234 ), .Y(
        \us02/n228 ) );
  OAI21XL \us02/U194  ( .A0(\us02/n58 ), .A1(\us02/n27 ), .B0(\us02/n247 ), 
        .Y(\us02/n245 ) );
  NOR2X1 \us02/U193  ( .A(sa02[7]), .B(\us02/n145 ), .Y(\us02/n246 ) );
  XNOR2X1 \us02/U192  ( .A(\us02/n69 ), .B(sa02[1]), .Y(\us02/n130 ) );
  MXI2X1 \us02/U191  ( .A(\us02/n245 ), .B(\us02/n246 ), .S0(\us02/n130 ), .Y(
        \us02/n243 ) );
  OAI211X1 \us02/U190  ( .A0(\us02/n4 ), .A1(\us02/n149 ), .B0(\us02/n243 ), 
        .C0(\us02/n244 ), .Y(\us02/n230 ) );
  NOR2X1 \us02/U189  ( .A(\us02/n242 ), .B(\us02/n137 ), .Y(\us02/n70 ) );
  OAI221XL \us02/U188  ( .A0(\us02/n159 ), .A1(\us02/n27 ), .B0(\us02/n20 ), 
        .B1(\us02/n34 ), .C0(\us02/n241 ), .Y(\us02/n231 ) );
  NAND2X1 \us02/U187  ( .A(\us02/n101 ), .B(\us02/n240 ), .Y(\us02/n76 ) );
  AOI21X1 \us02/U186  ( .A0(\us02/n122 ), .A1(\us02/n106 ), .B0(\us02/n129 ), 
        .Y(\us02/n237 ) );
  INVX1 \us02/U185  ( .A(\us02/n239 ), .Y(\us02/n238 ) );
  OAI21XL \us02/U184  ( .A0(\us02/n237 ), .A1(\us02/n43 ), .B0(\us02/n238 ), 
        .Y(\us02/n236 ) );
  OAI221XL \us02/U183  ( .A0(\us02/n18 ), .A1(\us02/n76 ), .B0(\us02/n59 ), 
        .B1(\us02/n27 ), .C0(\us02/n236 ), .Y(\us02/n232 ) );
  AOI2BB2X1 \us02/U182  ( .B0(\us02/n24 ), .B1(\us02/n187 ), .A0N(\us02/n227 ), 
        .A1N(\us02/n20 ), .Y(\us02/n235 ) );
  OAI211X1 \us02/U181  ( .A0(\us02/n27 ), .A1(\us02/n122 ), .B0(\us02/n158 ), 
        .C0(\us02/n235 ), .Y(\us02/n233 ) );
  MX4X1 \us02/U180  ( .A(\us02/n230 ), .B(\us02/n231 ), .C(\us02/n232 ), .D(
        \us02/n233 ), .S0(\us02/n234 ), .S1(sa02[5]), .Y(\us02/n229 ) );
  MX2X1 \us02/U179  ( .A(\us02/n228 ), .B(\us02/n229 ), .S0(sa02[6]), .Y(
        sa02_sr[3]) );
  NOR2BX1 \us02/U178  ( .AN(\us02/n204 ), .B(\us02/n137 ), .Y(\us02/n110 ) );
  INVX1 \us02/U177  ( .A(\us02/n110 ), .Y(\us02/n64 ) );
  AOI22X1 \us02/U176  ( .A0(\us02/n225 ), .A1(\us02/n226 ), .B0(\us02/n6 ), 
        .B1(\us02/n227 ), .Y(\us02/n224 ) );
  OAI221XL \us02/U175  ( .A0(\us02/n27 ), .A1(\us02/n64 ), .B0(\us02/n4 ), 
        .B1(\us02/n83 ), .C0(\us02/n224 ), .Y(\us02/n212 ) );
  NAND2X1 \us02/U174  ( .A(\us02/n34 ), .B(\us02/n204 ), .Y(\us02/n221 ) );
  OAI21XL \us02/U173  ( .A0(\us02/n69 ), .A1(\us02/n223 ), .B0(\us02/n27 ), 
        .Y(\us02/n222 ) );
  NOR2X1 \us02/U172  ( .A(\us02/n217 ), .B(\us02/n42 ), .Y(\us02/n208 ) );
  AOI211X1 \us02/U171  ( .A0(\us02/n208 ), .A1(\us02/n5 ), .B0(\us02/n220 ), 
        .C0(\us02/n173 ), .Y(\us02/n219 ) );
  OAI22X1 \us02/U170  ( .A0(\us02/n218 ), .A1(\us02/n10 ), .B0(\us02/n219 ), 
        .B1(\us02/n114 ), .Y(\us02/n213 ) );
  INVX1 \us02/U169  ( .A(\us02/n135 ), .Y(\us02/n215 ) );
  NOR2X1 \us02/U168  ( .A(\us02/n4 ), .B(\us02/n159 ), .Y(\us02/n31 ) );
  INVX1 \us02/U167  ( .A(\us02/n31 ), .Y(\us02/n196 ) );
  AOI31X1 \us02/U166  ( .A0(\us02/n215 ), .A1(\us02/n196 ), .A2(\us02/n216 ), 
        .B0(\us02/n52 ), .Y(\us02/n214 ) );
  AOI211X1 \us02/U165  ( .A0(\us02/n55 ), .A1(\us02/n212 ), .B0(\us02/n213 ), 
        .C0(\us02/n214 ), .Y(\us02/n190 ) );
  INVX1 \us02/U164  ( .A(\us02/n207 ), .Y(\us02/n192 ) );
  NOR2X1 \us02/U163  ( .A(\us02/n25 ), .B(\us02/n98 ), .Y(\us02/n32 ) );
  OAI22X1 \us02/U162  ( .A0(\us02/n28 ), .A1(\us02/n4 ), .B0(\us02/n188 ), 
        .B1(\us02/n27 ), .Y(\us02/n206 ) );
  NAND2X1 \us02/U161  ( .A(\us02/n204 ), .B(\us02/n80 ), .Y(\us02/n118 ) );
  INVX1 \us02/U160  ( .A(\us02/n118 ), .Y(\us02/n123 ) );
  NAND2X1 \us02/U159  ( .A(\us02/n94 ), .B(\us02/n79 ), .Y(\us02/n203 ) );
  OAI2BB1X1 \us02/U158  ( .A0N(\us02/n199 ), .A1N(\us02/n200 ), .B0(\us02/n33 ), .Y(\us02/n195 ) );
  INVX1 \us02/U157  ( .A(\us02/n55 ), .Y(\us02/n12 ) );
  AOI31X1 \us02/U156  ( .A0(\us02/n195 ), .A1(\us02/n196 ), .A2(\us02/n197 ), 
        .B0(\us02/n12 ), .Y(\us02/n194 ) );
  AOI211X1 \us02/U155  ( .A0(\us02/n89 ), .A1(\us02/n192 ), .B0(\us02/n193 ), 
        .C0(\us02/n194 ), .Y(\us02/n191 ) );
  MXI2X1 \us02/U154  ( .A(\us02/n190 ), .B(\us02/n191 ), .S0(sa02[6]), .Y(
        sa02_sr[4]) );
  OAI21XL \us02/U153  ( .A0(\us02/n69 ), .A1(\us02/n189 ), .B0(\us02/n27 ), 
        .Y(\us02/n186 ) );
  INVX1 \us02/U152  ( .A(\us02/n183 ), .Y(\us02/n180 ) );
  NAND2X1 \us02/U151  ( .A(\us02/n74 ), .B(\us02/n182 ), .Y(\us02/n181 ) );
  AOI211X1 \us02/U150  ( .A0(\us02/n179 ), .A1(\us02/n24 ), .B0(\us02/n180 ), 
        .C0(\us02/n181 ), .Y(\us02/n165 ) );
  INVX1 \us02/U149  ( .A(\us02/n178 ), .Y(\us02/n175 ) );
  AOI211X1 \us02/U148  ( .A0(\us02/n175 ), .A1(\us02/n5 ), .B0(\us02/n176 ), 
        .C0(\us02/n177 ), .Y(\us02/n174 ) );
  OAI221XL \us02/U147  ( .A0(\us02/n159 ), .A1(\us02/n27 ), .B0(\us02/n145 ), 
        .B1(\us02/n20 ), .C0(\us02/n174 ), .Y(\us02/n167 ) );
  MXI2X1 \us02/U146  ( .A(\us02/n40 ), .B(\us02/n173 ), .S0(\us02/n96 ), .Y(
        \us02/n170 ) );
  AOI22X1 \us02/U145  ( .A0(\us02/n137 ), .A1(\us02/n24 ), .B0(\us02/n172 ), 
        .B1(\us02/n6 ), .Y(\us02/n171 ) );
  OAI211X1 \us02/U144  ( .A0(\us02/n20 ), .A1(\us02/n169 ), .B0(\us02/n170 ), 
        .C0(\us02/n171 ), .Y(\us02/n168 ) );
  AOI22X1 \us02/U143  ( .A0(\us02/n89 ), .A1(\us02/n167 ), .B0(\us02/n55 ), 
        .B1(\us02/n168 ), .Y(\us02/n166 ) );
  OAI221XL \us02/U142  ( .A0(\us02/n164 ), .A1(\us02/n114 ), .B0(\us02/n165 ), 
        .B1(\us02/n52 ), .C0(\us02/n166 ), .Y(\us02/n138 ) );
  OAI21XL \us02/U141  ( .A0(\us02/n41 ), .A1(\us02/n163 ), .B0(\us02/n69 ), 
        .Y(\us02/n162 ) );
  AOI221X1 \us02/U140  ( .A0(\us02/n159 ), .A1(\us02/n24 ), .B0(\us02/n160 ), 
        .B1(\us02/n33 ), .C0(\us02/n161 ), .Y(\us02/n140 ) );
  OAI21XL \us02/U139  ( .A0(\us02/n157 ), .A1(\us02/n20 ), .B0(\us02/n158 ), 
        .Y(\us02/n156 ) );
  NOR2X1 \us02/U138  ( .A(\us02/n4 ), .B(\us02/n136 ), .Y(\us02/n153 ) );
  NOR2X1 \us02/U137  ( .A(\us02/n145 ), .B(\us02/n69 ), .Y(\us02/n154 ) );
  MXI2X1 \us02/U136  ( .A(\us02/n153 ), .B(\us02/n154 ), .S0(\us02/n155 ), .Y(
        \us02/n152 ) );
  OAI221XL \us02/U135  ( .A0(\us02/n110 ), .A1(\us02/n18 ), .B0(\us02/n20 ), 
        .B1(\us02/n151 ), .C0(\us02/n152 ), .Y(\us02/n143 ) );
  AOI21X1 \us02/U134  ( .A0(\us02/n149 ), .A1(\us02/n150 ), .B0(\us02/n18 ), 
        .Y(\us02/n148 ) );
  AOI2BB1X1 \us02/U133  ( .A0N(\us02/n147 ), .A1N(\us02/n27 ), .B0(\us02/n148 ), .Y(\us02/n146 ) );
  OAI221XL \us02/U132  ( .A0(\us02/n145 ), .A1(\us02/n20 ), .B0(\us02/n4 ), 
        .B1(\us02/n34 ), .C0(\us02/n146 ), .Y(\us02/n144 ) );
  AOI22X1 \us02/U131  ( .A0(\us02/n89 ), .A1(\us02/n143 ), .B0(\us02/n14 ), 
        .B1(\us02/n144 ), .Y(\us02/n142 ) );
  OAI221XL \us02/U130  ( .A0(\us02/n140 ), .A1(\us02/n12 ), .B0(\us02/n141 ), 
        .B1(\us02/n114 ), .C0(\us02/n142 ), .Y(\us02/n139 ) );
  MX2X1 \us02/U129  ( .A(\us02/n138 ), .B(\us02/n139 ), .S0(sa02[6]), .Y(
        sa02_sr[5]) );
  INVX1 \us02/U128  ( .A(\us02/n70 ), .Y(\us02/n133 ) );
  OAI22X1 \us02/U127  ( .A0(\us02/n4 ), .A1(\us02/n136 ), .B0(\us02/n137 ), 
        .B1(\us02/n27 ), .Y(\us02/n134 ) );
  AOI211X1 \us02/U126  ( .A0(\us02/n133 ), .A1(\us02/n69 ), .B0(\us02/n134 ), 
        .C0(\us02/n135 ), .Y(\us02/n112 ) );
  INVX1 \us02/U125  ( .A(\us02/n132 ), .Y(\us02/n131 ) );
  OAI21XL \us02/U124  ( .A0(\us02/n18 ), .A1(\us02/n37 ), .B0(\us02/n128 ), 
        .Y(\us02/n127 ) );
  OAI221XL \us02/U123  ( .A0(\us02/n18 ), .A1(\us02/n105 ), .B0(\us02/n123 ), 
        .B1(\us02/n27 ), .C0(\us02/n124 ), .Y(\us02/n116 ) );
  NAND2X1 \us02/U122  ( .A(\us02/n121 ), .B(\us02/n122 ), .Y(\us02/n30 ) );
  OAI221XL \us02/U121  ( .A0(\us02/n18 ), .A1(\us02/n118 ), .B0(\us02/n27 ), 
        .B1(\us02/n30 ), .C0(\us02/n119 ), .Y(\us02/n117 ) );
  AOI22X1 \us02/U120  ( .A0(\us02/n89 ), .A1(\us02/n116 ), .B0(\us02/n55 ), 
        .B1(\us02/n117 ), .Y(\us02/n115 ) );
  OAI221XL \us02/U119  ( .A0(\us02/n112 ), .A1(\us02/n52 ), .B0(\us02/n113 ), 
        .B1(\us02/n114 ), .C0(\us02/n115 ), .Y(\us02/n84 ) );
  OAI22X1 \us02/U118  ( .A0(\us02/n110 ), .A1(\us02/n4 ), .B0(\us02/n20 ), 
        .B1(\us02/n21 ), .Y(\us02/n108 ) );
  AOI21X1 \us02/U117  ( .A0(sa02[1]), .A1(\us02/n58 ), .B0(\us02/n27 ), .Y(
        \us02/n109 ) );
  AOI211X1 \us02/U116  ( .A0(\us02/n5 ), .A1(\us02/n107 ), .B0(\us02/n108 ), 
        .C0(\us02/n109 ), .Y(\us02/n86 ) );
  OAI22X1 \us02/U115  ( .A0(\us02/n45 ), .A1(\us02/n4 ), .B0(sa02[4]), .B1(
        \us02/n18 ), .Y(\us02/n103 ) );
  AOI21X1 \us02/U114  ( .A0(\us02/n105 ), .A1(\us02/n106 ), .B0(\us02/n20 ), 
        .Y(\us02/n104 ) );
  AOI211X1 \us02/U113  ( .A0(\us02/n33 ), .A1(\us02/n102 ), .B0(\us02/n103 ), 
        .C0(\us02/n104 ), .Y(\us02/n87 ) );
  NAND2X1 \us02/U112  ( .A(\us02/n100 ), .B(\us02/n101 ), .Y(\us02/n62 ) );
  OAI221XL \us02/U111  ( .A0(\us02/n27 ), .A1(\us02/n62 ), .B0(\us02/n4 ), 
        .B1(\us02/n21 ), .C0(\us02/n97 ), .Y(\us02/n90 ) );
  NOR3X1 \us02/U110  ( .A(\us02/n4 ), .B(\us02/n95 ), .C(\us02/n96 ), .Y(
        \us02/n67 ) );
  AOI31X1 \us02/U109  ( .A0(\us02/n79 ), .A1(\us02/n94 ), .A2(\us02/n6 ), .B0(
        \us02/n67 ), .Y(\us02/n93 ) );
  OAI221XL \us02/U108  ( .A0(\us02/n73 ), .A1(\us02/n27 ), .B0(\us02/n92 ), 
        .B1(\us02/n20 ), .C0(\us02/n93 ), .Y(\us02/n91 ) );
  AOI22X1 \us02/U107  ( .A0(\us02/n89 ), .A1(\us02/n90 ), .B0(\us02/n16 ), 
        .B1(\us02/n91 ), .Y(\us02/n88 ) );
  OAI221XL \us02/U106  ( .A0(\us02/n86 ), .A1(\us02/n52 ), .B0(\us02/n87 ), 
        .B1(\us02/n12 ), .C0(\us02/n88 ), .Y(\us02/n85 ) );
  MX2X1 \us02/U105  ( .A(\us02/n84 ), .B(\us02/n85 ), .S0(sa02[6]), .Y(
        sa02_sr[6]) );
  INVX1 \us02/U104  ( .A(\us02/n81 ), .Y(\us02/n77 ) );
  AOI21X1 \us02/U103  ( .A0(\us02/n79 ), .A1(\us02/n80 ), .B0(\us02/n27 ), .Y(
        \us02/n78 ) );
  AOI211X1 \us02/U102  ( .A0(\us02/n5 ), .A1(\us02/n76 ), .B0(\us02/n77 ), 
        .C0(\us02/n78 ), .Y(\us02/n51 ) );
  OAI211X1 \us02/U101  ( .A0(\us02/n73 ), .A1(\us02/n27 ), .B0(\us02/n74 ), 
        .C0(\us02/n75 ), .Y(\us02/n72 ) );
  AOI21X1 \us02/U100  ( .A0(\us02/n68 ), .A1(\us02/n69 ), .B0(\us02/n6 ), .Y(
        \us02/n63 ) );
  INVX1 \us02/U99  ( .A(\us02/n67 ), .Y(\us02/n66 ) );
  OAI221XL \us02/U98  ( .A0(\us02/n63 ), .A1(\us02/n64 ), .B0(\us02/n65 ), 
        .B1(\us02/n27 ), .C0(\us02/n66 ), .Y(\us02/n56 ) );
  AOI2BB2X1 \us02/U97  ( .B0(\us02/n61 ), .B1(\us02/n24 ), .A0N(\us02/n62 ), 
        .A1N(\us02/n20 ), .Y(\us02/n60 ) );
  OAI221XL \us02/U96  ( .A0(\us02/n58 ), .A1(\us02/n18 ), .B0(\us02/n59 ), 
        .B1(\us02/n27 ), .C0(\us02/n60 ), .Y(\us02/n57 ) );
  AOI22X1 \us02/U95  ( .A0(\us02/n55 ), .A1(\us02/n56 ), .B0(\us02/n16 ), .B1(
        \us02/n57 ), .Y(\us02/n54 ) );
  OAI221XL \us02/U94  ( .A0(\us02/n51 ), .A1(\us02/n52 ), .B0(\us02/n53 ), 
        .B1(\us02/n10 ), .C0(\us02/n54 ), .Y(\us02/n7 ) );
  INVX1 \us02/U93  ( .A(\us02/n50 ), .Y(\us02/n49 ) );
  OAI221XL \us02/U92  ( .A0(\us02/n47 ), .A1(\us02/n18 ), .B0(\us02/n27 ), 
        .B1(\us02/n48 ), .C0(\us02/n49 ), .Y(\us02/n46 ) );
  NOR2X1 \us02/U91  ( .A(\us02/n41 ), .B(\us02/n42 ), .Y(\us02/n38 ) );
  INVX1 \us02/U90  ( .A(\us02/n40 ), .Y(\us02/n39 ) );
  INVX1 \us02/U89  ( .A(\us02/n32 ), .Y(\us02/n26 ) );
  AOI21X1 \us02/U88  ( .A0(\us02/n5 ), .A1(\us02/n30 ), .B0(\us02/n31 ), .Y(
        \us02/n29 ) );
  OAI221XL \us02/U87  ( .A0(\us02/n26 ), .A1(\us02/n27 ), .B0(\us02/n28 ), 
        .B1(\us02/n20 ), .C0(\us02/n29 ), .Y(\us02/n15 ) );
  OAI221XL \us02/U86  ( .A0(\us02/n18 ), .A1(\us02/n19 ), .B0(\us02/n20 ), 
        .B1(\us02/n21 ), .C0(\us02/n22 ), .Y(\us02/n17 ) );
  AOI22X1 \us02/U85  ( .A0(\us02/n14 ), .A1(\us02/n15 ), .B0(\us02/n16 ), .B1(
        \us02/n17 ), .Y(\us02/n13 ) );
  OAI221XL \us02/U84  ( .A0(\us02/n9 ), .A1(\us02/n10 ), .B0(\us02/n11 ), .B1(
        \us02/n12 ), .C0(\us02/n13 ), .Y(\us02/n8 ) );
  MX2X1 \us02/U83  ( .A(\us02/n7 ), .B(\us02/n8 ), .S0(sa02[6]), .Y(sa02_sr[7]) );
  NOR2X4 \us02/U82  ( .A(\us02/n129 ), .B(sa02[2]), .Y(\us02/n43 ) );
  CLKINVX3 \us02/U81  ( .A(\us02/n14 ), .Y(\us02/n52 ) );
  OAI22XL \us02/U80  ( .A0(\us02/n201 ), .A1(\us02/n52 ), .B0(\us02/n202 ), 
        .B1(\us02/n114 ), .Y(\us02/n193 ) );
  CLKINVX3 \us02/U79  ( .A(sa02[5]), .Y(\us02/n252 ) );
  NOR2X2 \us02/U78  ( .A(\us02/n252 ), .B(\us02/n234 ), .Y(\us02/n55 ) );
  CLKINVX3 \us02/U77  ( .A(sa02[7]), .Y(\us02/n129 ) );
  NOR2X4 \us02/U76  ( .A(\us02/n129 ), .B(\us02/n69 ), .Y(\us02/n24 ) );
  AOI22XL \us02/U75  ( .A0(\us02/n70 ), .A1(\us02/n24 ), .B0(\us02/n96 ), .B1(
        \us02/n129 ), .Y(\us02/n241 ) );
  NOR2X2 \us02/U74  ( .A(\us02/n252 ), .B(sa02[0]), .Y(\us02/n89 ) );
  CLKINVX3 \us02/U73  ( .A(sa02[0]), .Y(\us02/n234 ) );
  NOR2X4 \us02/U72  ( .A(\us02/n69 ), .B(sa02[7]), .Y(\us02/n33 ) );
  INVX12 \us02/U71  ( .A(\us02/n33 ), .Y(\us02/n27 ) );
  CLKINVX3 \us02/U70  ( .A(\us02/n1 ), .Y(\us02/n6 ) );
  CLKINVX3 \us02/U69  ( .A(\us02/n1 ), .Y(\us02/n5 ) );
  INVXL \us02/U68  ( .A(\us02/n24 ), .Y(\us02/n36 ) );
  INVX4 \us02/U67  ( .A(\us02/n3 ), .Y(\us02/n4 ) );
  INVXL \us02/U66  ( .A(\us02/n36 ), .Y(\us02/n3 ) );
  INVX4 \us02/U65  ( .A(sa02[1]), .Y(\us02/n226 ) );
  INVX4 \us02/U64  ( .A(\us02/n43 ), .Y(\us02/n20 ) );
  AOI221X4 \us02/U63  ( .A0(\us02/n24 ), .A1(\us02/n82 ), .B0(\us02/n43 ), 
        .B1(\us02/n295 ), .C0(\us02/n173 ), .Y(\us02/n346 ) );
  AOI221X4 \us02/U62  ( .A0(\us02/n5 ), .A1(\us02/n96 ), .B0(\us02/n43 ), .B1(
        \us02/n239 ), .C0(\us02/n340 ), .Y(\us02/n336 ) );
  AOI222X4 \us02/U61  ( .A0(\us02/n59 ), .A1(\us02/n43 ), .B0(\us02/n6 ), .B1(
        \us02/n221 ), .C0(\us02/n222 ), .C1(\us02/n187 ), .Y(\us02/n218 ) );
  AOI222X4 \us02/U60  ( .A0(\us02/n123 ), .A1(\us02/n43 ), .B0(sa02[2]), .B1(
        \us02/n203 ), .C0(\us02/n6 ), .C1(\us02/n71 ), .Y(\us02/n202 ) );
  AOI221X4 \us02/U59  ( .A0(\us02/n314 ), .A1(\us02/n43 ), .B0(\us02/n160 ), 
        .B1(\us02/n24 ), .C0(\us02/n315 ), .Y(\us02/n307 ) );
  AOI221X4 \us02/U58  ( .A0(\us02/n43 ), .A1(\us02/n208 ), .B0(\us02/n76 ), 
        .B1(\us02/n24 ), .C0(\us02/n209 ), .Y(\us02/n207 ) );
  AOI221X4 \us02/U57  ( .A0(\us02/n43 ), .A1(\us02/n205 ), .B0(\us02/n32 ), 
        .B1(\us02/n6 ), .C0(\us02/n206 ), .Y(\us02/n201 ) );
  AOI221X4 \us02/U56  ( .A0(\us02/n43 ), .A1(\us02/n44 ), .B0(\us02/n45 ), 
        .B1(\us02/n24 ), .C0(\us02/n46 ), .Y(\us02/n9 ) );
  AOI22XL \us02/U55  ( .A0(\us02/n217 ), .A1(\us02/n43 ), .B0(\us02/n33 ), 
        .B1(\us02/n47 ), .Y(\us02/n216 ) );
  AOI22XL \us02/U54  ( .A0(\us02/n98 ), .A1(\us02/n43 ), .B0(\us02/n6 ), .B1(
        \us02/n99 ), .Y(\us02/n97 ) );
  AOI22XL \us02/U53  ( .A0(\us02/n82 ), .A1(\us02/n43 ), .B0(\us02/n83 ), .B1(
        \us02/n24 ), .Y(\us02/n81 ) );
  AOI2BB2XL \us02/U52  ( .B0(\us02/n43 ), .B1(\us02/n94 ), .A0N(\us02/n120 ), 
        .A1N(\us02/n4 ), .Y(\us02/n119 ) );
  AOI222X4 \us02/U51  ( .A0(\us02/n125 ), .A1(\us02/n33 ), .B0(\us02/n145 ), 
        .B1(\us02/n40 ), .C0(\us02/n43 ), .C1(\us02/n184 ), .Y(\us02/n183 ) );
  AOI22XL \us02/U50  ( .A0(\us02/n43 ), .A1(\us02/n303 ), .B0(\us02/n24 ), 
        .B1(\us02/n96 ), .Y(\us02/n358 ) );
  AOI22XL \us02/U49  ( .A0(\us02/n43 ), .A1(\us02/n100 ), .B0(\us02/n24 ), 
        .B1(\us02/n125 ), .Y(\us02/n124 ) );
  AOI21XL \us02/U48  ( .A0(\us02/n159 ), .A1(\us02/n43 ), .B0(\us02/n40 ), .Y(
        \us02/n262 ) );
  AOI22XL \us02/U47  ( .A0(\us02/n40 ), .A1(\us02/n94 ), .B0(\us02/n43 ), .B1(
        \us02/n187 ), .Y(\us02/n244 ) );
  AOI22XL \us02/U46  ( .A0(\us02/n184 ), .A1(\us02/n5 ), .B0(\us02/n198 ), 
        .B1(\us02/n43 ), .Y(\us02/n197 ) );
  NOR2XL \us02/U45  ( .A(\us02/n33 ), .B(\us02/n2 ), .Y(\us02/n302 ) );
  MXI2XL \us02/U44  ( .A(\us02/n2 ), .B(\us02/n6 ), .S0(\us02/n28 ), .Y(
        \us02/n311 ) );
  INVXL \us02/U43  ( .A(\us02/n20 ), .Y(\us02/n2 ) );
  INVX4 \us02/U42  ( .A(\us02/n6 ), .Y(\us02/n18 ) );
  AOI21XL \us02/U41  ( .A0(\us02/n18 ), .A1(\us02/n162 ), .B0(\us02/n25 ), .Y(
        \us02/n161 ) );
  INVX4 \us02/U40  ( .A(sa02[2]), .Y(\us02/n69 ) );
  NOR2X4 \us02/U39  ( .A(\us02/n226 ), .B(\us02/n4 ), .Y(\us02/n40 ) );
  CLKINVX3 \us02/U38  ( .A(sa02[3]), .Y(\us02/n136 ) );
  NOR2X2 \us02/U37  ( .A(\us02/n136 ), .B(sa02[4]), .Y(\us02/n145 ) );
  CLKINVX3 \us02/U36  ( .A(sa02[4]), .Y(\us02/n58 ) );
  NOR2X2 \us02/U35  ( .A(\us02/n58 ), .B(sa02[3]), .Y(\us02/n159 ) );
  NOR2X2 \us02/U34  ( .A(\us02/n136 ), .B(\us02/n58 ), .Y(\us02/n259 ) );
  NOR2X2 \us02/U33  ( .A(sa02[4]), .B(sa02[3]), .Y(\us02/n278 ) );
  NOR2X2 \us02/U32  ( .A(\us02/n259 ), .B(\us02/n278 ), .Y(\us02/n47 ) );
  CLKINVX3 \us02/U31  ( .A(\us02/n259 ), .Y(\us02/n44 ) );
  NOR2X2 \us02/U30  ( .A(\us02/n44 ), .B(sa02[1]), .Y(\us02/n137 ) );
  AOI21XL \us02/U29  ( .A0(\us02/n44 ), .A1(\us02/n111 ), .B0(\us02/n4 ), .Y(
        \us02/n177 ) );
  AOI22XL \us02/U28  ( .A0(\us02/n23 ), .A1(\us02/n24 ), .B0(\us02/n25 ), .B1(
        sa02[2]), .Y(\us02/n22 ) );
  AOI22XL \us02/U27  ( .A0(\us02/n33 ), .A1(sa02[3]), .B0(\us02/n24 ), .B1(
        \us02/n58 ), .Y(\us02/n277 ) );
  NAND2XL \us02/U26  ( .A(\us02/n198 ), .B(\us02/n24 ), .Y(\us02/n132 ) );
  OAI2BB2XL \us02/U25  ( .B0(\us02/n20 ), .B1(\us02/n111 ), .A0N(\us02/n125 ), 
        .A1N(\us02/n24 ), .Y(\us02/n220 ) );
  NAND2XL \us02/U24  ( .A(\us02/n111 ), .B(\us02/n101 ), .Y(\us02/n21 ) );
  NAND2XL \us02/U23  ( .A(\us02/n111 ), .B(\us02/n300 ), .Y(\us02/n187 ) );
  NAND2XL \us02/U22  ( .A(\us02/n111 ), .B(\us02/n121 ), .Y(\us02/n303 ) );
  AOI221XL \us02/U21  ( .A0(\us02/n43 ), .A1(\us02/n151 ), .B0(\us02/n25 ), 
        .B1(\us02/n69 ), .C0(\us02/n275 ), .Y(\us02/n274 ) );
  NOR2BXL \us02/U20  ( .AN(\us02/n101 ), .B(\us02/n25 ), .Y(\us02/n172 ) );
  NAND2X2 \us02/U19  ( .A(\us02/n58 ), .B(\us02/n226 ), .Y(\us02/n34 ) );
  OAI222X1 \us02/U18  ( .A0(\us02/n27 ), .A1(\us02/n34 ), .B0(\us02/n69 ), 
        .B1(\us02/n205 ), .C0(\us02/n20 ), .C1(\us02/n79 ), .Y(\us02/n260 ) );
  OAI222X1 \us02/U17  ( .A0(\us02/n20 ), .A1(\us02/n99 ), .B0(\us02/n27 ), 
        .B1(\us02/n101 ), .C0(\us02/n184 ), .C1(\us02/n4 ), .Y(\us02/n250 ) );
  OAI222X1 \us02/U16  ( .A0(\us02/n4 ), .A1(\us02/n37 ), .B0(\us02/n38 ), .B1(
        \us02/n20 ), .C0(sa02[4]), .C1(\us02/n39 ), .Y(\us02/n35 ) );
  AOI221X1 \us02/U15  ( .A0(\us02/n5 ), .A1(\us02/n19 ), .B0(\us02/n33 ), .B1(
        \us02/n34 ), .C0(\us02/n35 ), .Y(\us02/n11 ) );
  OR2X2 \us02/U14  ( .A(sa02[2]), .B(sa02[7]), .Y(\us02/n1 ) );
  AOI221XL \us02/U13  ( .A0(\us02/n70 ), .A1(\us02/n43 ), .B0(\us02/n24 ), 
        .B1(\us02/n71 ), .C0(\us02/n72 ), .Y(\us02/n53 ) );
  AOI221XL \us02/U12  ( .A0(\us02/n59 ), .A1(\us02/n33 ), .B0(\us02/n43 ), 
        .B1(\us02/n126 ), .C0(\us02/n127 ), .Y(\us02/n113 ) );
  AOI222XL \us02/U11  ( .A0(\us02/n185 ), .A1(\us02/n43 ), .B0(\us02/n186 ), 
        .B1(\us02/n187 ), .C0(\us02/n6 ), .C1(\us02/n188 ), .Y(\us02/n164 ) );
  AOI221X1 \us02/U10  ( .A0(\us02/n313 ), .A1(\us02/n5 ), .B0(\us02/n23 ), 
        .B1(\us02/n2 ), .C0(\us02/n328 ), .Y(\us02/n320 ) );
  AOI221X1 \us02/U9  ( .A0(\us02/n40 ), .A1(\us02/n136 ), .B0(\us02/n33 ), 
        .B1(\us02/n178 ), .C0(\us02/n338 ), .Y(\us02/n337 ) );
  AOI222XL \us02/U8  ( .A0(\us02/n278 ), .A1(\us02/n24 ), .B0(\us02/n42 ), 
        .B1(\us02/n33 ), .C0(\us02/n43 ), .C1(\us02/n136 ), .Y(\us02/n351 ) );
  AOI31X1 \us02/U7  ( .A0(sa02[2]), .A1(\us02/n58 ), .A2(sa02[1]), .B0(
        \us02/n40 ), .Y(\us02/n350 ) );
  AOI31X1 \us02/U6  ( .A0(\us02/n44 ), .A1(\us02/n129 ), .A2(\us02/n130 ), 
        .B0(\us02/n131 ), .Y(\us02/n128 ) );
  AOI221X1 \us02/U5  ( .A0(\us02/n40 ), .A1(\us02/n136 ), .B0(\us02/n33 ), 
        .B1(\us02/n47 ), .C0(\us02/n156 ), .Y(\us02/n141 ) );
  OAI32X1 \us02/U4  ( .A0(\us02/n210 ), .A1(\us02/n145 ), .A2(\us02/n18 ), 
        .B0(\us02/n27 ), .B1(\us02/n211 ), .Y(\us02/n209 ) );
  AOI221X1 \us02/U3  ( .A0(\us02/n278 ), .A1(\us02/n40 ), .B0(\us02/n185 ), 
        .B1(\us02/n2 ), .C0(\us02/n279 ), .Y(\us02/n273 ) );
  OAI32X1 \us02/U2  ( .A0(\us02/n18 ), .A1(sa02[1]), .A2(\us02/n159 ), .B0(
        sa02[4]), .B1(\us02/n182 ), .Y(\us02/n318 ) );
  AOI31XL \us02/U1  ( .A0(\us02/n79 ), .A1(\us02/n44 ), .A2(\us02/n2 ), .B0(
        \us02/n280 ), .Y(\us02/n339 ) );
  NAND2X1 \us03/U366  ( .A(\us03/n47 ), .B(\us03/n226 ), .Y(\us03/n189 ) );
  NOR2X1 \us03/U365  ( .A(\us03/n226 ), .B(sa03[3]), .Y(\us03/n242 ) );
  INVX1 \us03/U364  ( .A(\us03/n242 ), .Y(\us03/n205 ) );
  AND2X1 \us03/U363  ( .A(\us03/n189 ), .B(\us03/n205 ), .Y(\us03/n65 ) );
  NOR2X1 \us03/U362  ( .A(\us03/n226 ), .B(\us03/n47 ), .Y(\us03/n45 ) );
  NOR2X1 \us03/U361  ( .A(\us03/n259 ), .B(\us03/n45 ), .Y(\us03/n73 ) );
  NAND2BX1 \us03/U360  ( .AN(\us03/n73 ), .B(\us03/n6 ), .Y(\us03/n158 ) );
  NOR2X1 \us03/U359  ( .A(\us03/n226 ), .B(\us03/n159 ), .Y(\us03/n95 ) );
  INVX1 \us03/U358  ( .A(\us03/n95 ), .Y(\us03/n111 ) );
  NOR2X1 \us03/U357  ( .A(\us03/n145 ), .B(sa03[1]), .Y(\us03/n42 ) );
  INVX1 \us03/U356  ( .A(\us03/n42 ), .Y(\us03/n121 ) );
  INVX1 \us03/U355  ( .A(\us03/n47 ), .Y(\us03/n96 ) );
  OAI211X1 \us03/U354  ( .A0(\us03/n65 ), .A1(\us03/n27 ), .B0(\us03/n158 ), 
        .C0(\us03/n358 ), .Y(\us03/n355 ) );
  NOR2X1 \us03/U353  ( .A(\us03/n226 ), .B(\us03/n145 ), .Y(\us03/n59 ) );
  NOR2X1 \us03/U352  ( .A(\us03/n96 ), .B(\us03/n59 ), .Y(\us03/n271 ) );
  NOR2X1 \us03/U351  ( .A(\us03/n226 ), .B(\us03/n278 ), .Y(\us03/n217 ) );
  INVX1 \us03/U350  ( .A(\us03/n217 ), .Y(\us03/n150 ) );
  NAND2X1 \us03/U349  ( .A(\us03/n44 ), .B(\us03/n150 ), .Y(\us03/n147 ) );
  NAND2X1 \us03/U348  ( .A(sa03[4]), .B(\us03/n226 ), .Y(\us03/n101 ) );
  INVX1 \us03/U347  ( .A(\us03/n159 ), .Y(\us03/n188 ) );
  NOR2X1 \us03/U346  ( .A(\us03/n188 ), .B(\us03/n226 ), .Y(\us03/n25 ) );
  INVX1 \us03/U345  ( .A(\us03/n172 ), .Y(\us03/n107 ) );
  AOI22X1 \us03/U344  ( .A0(\us03/n33 ), .A1(\us03/n147 ), .B0(\us03/n24 ), 
        .B1(\us03/n107 ), .Y(\us03/n357 ) );
  OAI221XL \us03/U343  ( .A0(\us03/n18 ), .A1(\us03/n121 ), .B0(\us03/n271 ), 
        .B1(\us03/n20 ), .C0(\us03/n357 ), .Y(\us03/n356 ) );
  MXI2X1 \us03/U342  ( .A(\us03/n355 ), .B(\us03/n356 ), .S0(\us03/n252 ), .Y(
        \us03/n331 ) );
  INVX1 \us03/U341  ( .A(\us03/n59 ), .Y(\us03/n79 ) );
  AND2X1 \us03/U340  ( .A(\us03/n101 ), .B(\us03/n79 ), .Y(\us03/n325 ) );
  XNOR2X1 \us03/U339  ( .A(sa03[5]), .B(\us03/n226 ), .Y(\us03/n352 ) );
  NOR2X1 \us03/U338  ( .A(\us03/n226 ), .B(\us03/n136 ), .Y(\us03/n281 ) );
  INVX1 \us03/U337  ( .A(\us03/n281 ), .Y(\us03/n19 ) );
  NAND2X1 \us03/U336  ( .A(\us03/n145 ), .B(\us03/n226 ), .Y(\us03/n223 ) );
  AOI21X1 \us03/U335  ( .A0(\us03/n19 ), .A1(\us03/n223 ), .B0(\us03/n27 ), 
        .Y(\us03/n354 ) );
  AOI31X1 \us03/U334  ( .A0(\us03/n6 ), .A1(\us03/n352 ), .A2(\us03/n259 ), 
        .B0(\us03/n354 ), .Y(\us03/n353 ) );
  OAI221XL \us03/U333  ( .A0(\us03/n20 ), .A1(\us03/n34 ), .B0(\us03/n325 ), 
        .B1(\us03/n4 ), .C0(\us03/n353 ), .Y(\us03/n347 ) );
  INVX1 \us03/U332  ( .A(\us03/n352 ), .Y(\us03/n349 ) );
  NAND2X1 \us03/U331  ( .A(\us03/n278 ), .B(\us03/n6 ), .Y(\us03/n74 ) );
  OAI211X1 \us03/U330  ( .A0(\us03/n349 ), .A1(\us03/n74 ), .B0(\us03/n350 ), 
        .C0(\us03/n351 ), .Y(\us03/n348 ) );
  MXI2X1 \us03/U329  ( .A(\us03/n347 ), .B(\us03/n348 ), .S0(\us03/n252 ), .Y(
        \us03/n332 ) );
  NOR2X1 \us03/U328  ( .A(\us03/n44 ), .B(\us03/n226 ), .Y(\us03/n157 ) );
  INVX1 \us03/U327  ( .A(\us03/n157 ), .Y(\us03/n240 ) );
  NAND2X1 \us03/U326  ( .A(\us03/n240 ), .B(\us03/n189 ), .Y(\us03/n68 ) );
  NOR2X1 \us03/U325  ( .A(\us03/n20 ), .B(\us03/n159 ), .Y(\us03/n225 ) );
  NOR2X1 \us03/U324  ( .A(\us03/n225 ), .B(\us03/n40 ), .Y(\us03/n345 ) );
  INVX1 \us03/U323  ( .A(\us03/n278 ), .Y(\us03/n94 ) );
  NAND2X1 \us03/U322  ( .A(\us03/n94 ), .B(\us03/n226 ), .Y(\us03/n199 ) );
  NAND2X1 \us03/U321  ( .A(\us03/n199 ), .B(\us03/n205 ), .Y(\us03/n82 ) );
  NAND2X1 \us03/U320  ( .A(\us03/n19 ), .B(\us03/n199 ), .Y(\us03/n295 ) );
  NOR2X1 \us03/U319  ( .A(\us03/n226 ), .B(\us03/n259 ), .Y(\us03/n210 ) );
  NOR2X1 \us03/U318  ( .A(\us03/n27 ), .B(\us03/n210 ), .Y(\us03/n173 ) );
  MXI2X1 \us03/U317  ( .A(\us03/n345 ), .B(\us03/n346 ), .S0(\us03/n252 ), .Y(
        \us03/n342 ) );
  NOR2X1 \us03/U316  ( .A(sa03[1]), .B(sa03[3]), .Y(\us03/n163 ) );
  INVX1 \us03/U315  ( .A(\us03/n163 ), .Y(\us03/n37 ) );
  INVX1 \us03/U314  ( .A(\us03/n173 ), .Y(\us03/n344 ) );
  AOI21X1 \us03/U313  ( .A0(\us03/n240 ), .A1(\us03/n37 ), .B0(\us03/n344 ), 
        .Y(\us03/n343 ) );
  AOI211X1 \us03/U312  ( .A0(\us03/n5 ), .A1(\us03/n68 ), .B0(\us03/n342 ), 
        .C0(\us03/n343 ), .Y(\us03/n333 ) );
  NOR2X1 \us03/U311  ( .A(\us03/n18 ), .B(\us03/n226 ), .Y(\us03/n258 ) );
  NAND2X1 \us03/U310  ( .A(\us03/n278 ), .B(sa03[1]), .Y(\us03/n204 ) );
  NOR2X1 \us03/U309  ( .A(\us03/n188 ), .B(sa03[1]), .Y(\us03/n179 ) );
  INVX1 \us03/U308  ( .A(\us03/n179 ), .Y(\us03/n330 ) );
  NAND2X1 \us03/U307  ( .A(\us03/n204 ), .B(\us03/n330 ), .Y(\us03/n239 ) );
  NOR2X1 \us03/U306  ( .A(\us03/n136 ), .B(sa03[1]), .Y(\us03/n299 ) );
  NOR2X1 \us03/U305  ( .A(\us03/n299 ), .B(\us03/n210 ), .Y(\us03/n341 ) );
  OAI32X1 \us03/U304  ( .A0(\us03/n27 ), .A1(\us03/n278 ), .A2(\us03/n95 ), 
        .B0(\us03/n341 ), .B1(\us03/n4 ), .Y(\us03/n340 ) );
  INVX1 \us03/U303  ( .A(\us03/n45 ), .Y(\us03/n126 ) );
  NAND2X1 \us03/U302  ( .A(\us03/n126 ), .B(\us03/n101 ), .Y(\us03/n178 ) );
  NOR2X1 \us03/U301  ( .A(\us03/n18 ), .B(\us03/n136 ), .Y(\us03/n280 ) );
  OAI21XL \us03/U300  ( .A0(\us03/n4 ), .A1(\us03/n121 ), .B0(\us03/n339 ), 
        .Y(\us03/n338 ) );
  MXI2X1 \us03/U299  ( .A(\us03/n336 ), .B(\us03/n337 ), .S0(\us03/n252 ), .Y(
        \us03/n335 ) );
  NOR2X1 \us03/U298  ( .A(\us03/n258 ), .B(\us03/n335 ), .Y(\us03/n334 ) );
  MX4X1 \us03/U297  ( .A(\us03/n331 ), .B(\us03/n332 ), .C(\us03/n333 ), .D(
        \us03/n334 ), .S0(sa03[6]), .S1(\us03/n234 ), .Y(sa03_sr[0]) );
  INVX1 \us03/U296  ( .A(\us03/n299 ), .Y(\us03/n80 ) );
  NOR2X1 \us03/U295  ( .A(\us03/n111 ), .B(\us03/n18 ), .Y(\us03/n269 ) );
  INVX1 \us03/U294  ( .A(\us03/n269 ), .Y(\us03/n75 ) );
  OAI221XL \us03/U293  ( .A0(\us03/n18 ), .A1(\us03/n330 ), .B0(\us03/n20 ), 
        .B1(\us03/n80 ), .C0(\us03/n75 ), .Y(\us03/n329 ) );
  AOI221X1 \us03/U292  ( .A0(\us03/n325 ), .A1(\us03/n33 ), .B0(\us03/n24 ), 
        .B1(\us03/n303 ), .C0(\us03/n329 ), .Y(\us03/n319 ) );
  NOR2X1 \us03/U291  ( .A(\us03/n234 ), .B(sa03[5]), .Y(\us03/n14 ) );
  NOR2X1 \us03/U290  ( .A(\us03/n25 ), .B(\us03/n299 ), .Y(\us03/n313 ) );
  NAND2X1 \us03/U289  ( .A(\us03/n44 ), .B(\us03/n226 ), .Y(\us03/n300 ) );
  AND2X1 \us03/U288  ( .A(\us03/n300 ), .B(\us03/n240 ), .Y(\us03/n23 ) );
  OAI32X1 \us03/U287  ( .A0(\us03/n4 ), .A1(\us03/n145 ), .A2(\us03/n210 ), 
        .B0(\us03/n137 ), .B1(\us03/n27 ), .Y(\us03/n328 ) );
  NOR2X1 \us03/U286  ( .A(sa03[0]), .B(sa03[5]), .Y(\us03/n16 ) );
  INVX1 \us03/U285  ( .A(\us03/n16 ), .Y(\us03/n114 ) );
  INVX1 \us03/U284  ( .A(\us03/n145 ), .Y(\us03/n149 ) );
  NOR2X1 \us03/U283  ( .A(\us03/n47 ), .B(sa03[1]), .Y(\us03/n98 ) );
  INVX1 \us03/U282  ( .A(\us03/n98 ), .Y(\us03/n284 ) );
  OAI21XL \us03/U281  ( .A0(\us03/n69 ), .A1(\us03/n284 ), .B0(\us03/n27 ), 
        .Y(\us03/n327 ) );
  AOI31X1 \us03/U280  ( .A0(\us03/n111 ), .A1(\us03/n149 ), .A2(\us03/n327 ), 
        .B0(\us03/n225 ), .Y(\us03/n326 ) );
  OAI21XL \us03/U279  ( .A0(\us03/n325 ), .A1(\us03/n18 ), .B0(\us03/n326 ), 
        .Y(\us03/n322 ) );
  NAND2X1 \us03/U278  ( .A(\us03/n19 ), .B(\us03/n189 ), .Y(\us03/n71 ) );
  NOR2X1 \us03/U277  ( .A(\us03/n71 ), .B(\us03/n18 ), .Y(\us03/n135 ) );
  AOI21X1 \us03/U276  ( .A0(\us03/n40 ), .A1(sa03[4]), .B0(\us03/n135 ), .Y(
        \us03/n324 ) );
  OAI221XL \us03/U275  ( .A0(\us03/n47 ), .A1(\us03/n27 ), .B0(\us03/n65 ), 
        .B1(\us03/n20 ), .C0(\us03/n324 ), .Y(\us03/n323 ) );
  AOI22X1 \us03/U274  ( .A0(\us03/n55 ), .A1(\us03/n322 ), .B0(\us03/n89 ), 
        .B1(\us03/n323 ), .Y(\us03/n321 ) );
  OAI221XL \us03/U273  ( .A0(\us03/n319 ), .A1(\us03/n52 ), .B0(\us03/n320 ), 
        .B1(\us03/n114 ), .C0(\us03/n321 ), .Y(\us03/n304 ) );
  NOR2X1 \us03/U272  ( .A(\us03/n226 ), .B(\us03/n58 ), .Y(\us03/n290 ) );
  INVX1 \us03/U271  ( .A(\us03/n290 ), .Y(\us03/n200 ) );
  NAND2X1 \us03/U270  ( .A(\us03/n34 ), .B(\us03/n200 ), .Y(\us03/n120 ) );
  INVX1 \us03/U269  ( .A(\us03/n210 ), .Y(\us03/n100 ) );
  OAI221XL \us03/U268  ( .A0(\us03/n20 ), .A1(\us03/n100 ), .B0(sa03[3]), .B1(
        \us03/n4 ), .C0(\us03/n262 ), .Y(\us03/n317 ) );
  INVX1 \us03/U267  ( .A(\us03/n258 ), .Y(\us03/n182 ) );
  AOI211X1 \us03/U266  ( .A0(\us03/n33 ), .A1(\us03/n120 ), .B0(\us03/n317 ), 
        .C0(\us03/n318 ), .Y(\us03/n306 ) );
  NAND2X1 \us03/U265  ( .A(\us03/n100 ), .B(\us03/n199 ), .Y(\us03/n151 ) );
  INVX1 \us03/U264  ( .A(\us03/n151 ), .Y(\us03/n314 ) );
  NOR2X1 \us03/U263  ( .A(\us03/n45 ), .B(\us03/n163 ), .Y(\us03/n160 ) );
  INVX1 \us03/U262  ( .A(\us03/n295 ), .Y(\us03/n92 ) );
  AOI21X1 \us03/U261  ( .A0(sa03[1]), .A1(\us03/n58 ), .B0(\us03/n98 ), .Y(
        \us03/n316 ) );
  OAI22X1 \us03/U260  ( .A0(\us03/n92 ), .A1(\us03/n18 ), .B0(\us03/n316 ), 
        .B1(\us03/n27 ), .Y(\us03/n315 ) );
  NOR2X1 \us03/U259  ( .A(\us03/n149 ), .B(\us03/n226 ), .Y(\us03/n41 ) );
  INVX1 \us03/U258  ( .A(\us03/n41 ), .Y(\us03/n105 ) );
  NAND2X1 \us03/U257  ( .A(\us03/n284 ), .B(\us03/n105 ), .Y(\us03/n227 ) );
  AOI21X1 \us03/U256  ( .A0(\us03/n313 ), .A1(\us03/n33 ), .B0(\us03/n269 ), 
        .Y(\us03/n312 ) );
  OAI221XL \us03/U255  ( .A0(\us03/n149 ), .A1(\us03/n20 ), .B0(\us03/n4 ), 
        .B1(\us03/n227 ), .C0(\us03/n312 ), .Y(\us03/n309 ) );
  AOI21X1 \us03/U254  ( .A0(\us03/n226 ), .A1(\us03/n188 ), .B0(\us03/n242 ), 
        .Y(\us03/n185 ) );
  INVX1 \us03/U253  ( .A(\us03/n185 ), .Y(\us03/n48 ) );
  AND2X1 \us03/U252  ( .A(\us03/n223 ), .B(\us03/n240 ), .Y(\us03/n28 ) );
  OAI221XL \us03/U251  ( .A0(\us03/n27 ), .A1(\us03/n44 ), .B0(\us03/n4 ), 
        .B1(\us03/n48 ), .C0(\us03/n311 ), .Y(\us03/n310 ) );
  AOI22X1 \us03/U250  ( .A0(\us03/n89 ), .A1(\us03/n309 ), .B0(\us03/n55 ), 
        .B1(\us03/n310 ), .Y(\us03/n308 ) );
  OAI221XL \us03/U249  ( .A0(\us03/n306 ), .A1(\us03/n52 ), .B0(\us03/n307 ), 
        .B1(\us03/n114 ), .C0(\us03/n308 ), .Y(\us03/n305 ) );
  MX2X1 \us03/U248  ( .A(\us03/n304 ), .B(\us03/n305 ), .S0(sa03[6]), .Y(
        sa03_sr[1]) );
  INVX1 \us03/U247  ( .A(\us03/n187 ), .Y(\us03/n61 ) );
  MXI2X1 \us03/U246  ( .A(\us03/n303 ), .B(\us03/n61 ), .S0(\us03/n69 ), .Y(
        \us03/n301 ) );
  MXI2X1 \us03/U245  ( .A(\us03/n301 ), .B(\us03/n147 ), .S0(\us03/n302 ), .Y(
        \us03/n285 ) );
  NAND2X1 \us03/U244  ( .A(\us03/n200 ), .B(\us03/n300 ), .Y(\us03/n99 ) );
  INVX1 \us03/U243  ( .A(\us03/n99 ), .Y(\us03/n296 ) );
  NOR2X1 \us03/U242  ( .A(\us03/n299 ), .B(\us03/n242 ), .Y(\us03/n298 ) );
  NAND2X1 \us03/U241  ( .A(sa03[1]), .B(\us03/n47 ), .Y(\us03/n122 ) );
  NOR2X1 \us03/U240  ( .A(\us03/n159 ), .B(\us03/n217 ), .Y(\us03/n198 ) );
  OAI221XL \us03/U239  ( .A0(\us03/n298 ), .A1(\us03/n27 ), .B0(\us03/n20 ), 
        .B1(\us03/n122 ), .C0(\us03/n132 ), .Y(\us03/n297 ) );
  AOI221X1 \us03/U238  ( .A0(\us03/n225 ), .A1(\us03/n226 ), .B0(\us03/n296 ), 
        .B1(\us03/n6 ), .C0(\us03/n297 ), .Y(\us03/n291 ) );
  OAI2BB2X1 \us03/U237  ( .B0(\us03/n27 ), .B1(\us03/n295 ), .A0N(\us03/n34 ), 
        .A1N(\us03/n24 ), .Y(\us03/n293 ) );
  AOI21X1 \us03/U236  ( .A0(\us03/n101 ), .A1(\us03/n150 ), .B0(\us03/n20 ), 
        .Y(\us03/n294 ) );
  AOI211X1 \us03/U235  ( .A0(\us03/n5 ), .A1(\us03/n79 ), .B0(\us03/n293 ), 
        .C0(\us03/n294 ), .Y(\us03/n292 ) );
  INVX1 \us03/U234  ( .A(\us03/n89 ), .Y(\us03/n10 ) );
  OAI22X1 \us03/U233  ( .A0(\us03/n291 ), .A1(\us03/n114 ), .B0(\us03/n292 ), 
        .B1(\us03/n10 ), .Y(\us03/n286 ) );
  INVX1 \us03/U232  ( .A(\us03/n225 ), .Y(\us03/n288 ) );
  NAND2X1 \us03/U231  ( .A(\us03/n200 ), .B(\us03/n284 ), .Y(\us03/n102 ) );
  NOR2X1 \us03/U230  ( .A(\us03/n290 ), .B(\us03/n163 ), .Y(\us03/n184 ) );
  AOI22X1 \us03/U229  ( .A0(\us03/n102 ), .A1(\us03/n69 ), .B0(\us03/n184 ), 
        .B1(\us03/n33 ), .Y(\us03/n289 ) );
  AOI31X1 \us03/U228  ( .A0(\us03/n132 ), .A1(\us03/n288 ), .A2(\us03/n289 ), 
        .B0(\us03/n52 ), .Y(\us03/n287 ) );
  AOI211X1 \us03/U227  ( .A0(\us03/n285 ), .A1(\us03/n55 ), .B0(\us03/n286 ), 
        .C0(\us03/n287 ), .Y(\us03/n263 ) );
  NAND2X1 \us03/U226  ( .A(\us03/n284 ), .B(\us03/n122 ), .Y(\us03/n125 ) );
  NOR2X1 \us03/U225  ( .A(\us03/n199 ), .B(\us03/n4 ), .Y(\us03/n50 ) );
  AOI21X1 \us03/U224  ( .A0(\us03/n200 ), .A1(\us03/n223 ), .B0(\us03/n20 ), 
        .Y(\us03/n283 ) );
  AOI211X1 \us03/U223  ( .A0(\us03/n5 ), .A1(\us03/n125 ), .B0(\us03/n50 ), 
        .C0(\us03/n283 ), .Y(\us03/n282 ) );
  OAI221XL \us03/U222  ( .A0(\us03/n281 ), .A1(\us03/n27 ), .B0(\us03/n4 ), 
        .B1(\us03/n111 ), .C0(\us03/n282 ), .Y(\us03/n265 ) );
  INVX1 \us03/U221  ( .A(\us03/n280 ), .Y(\us03/n247 ) );
  NAND2X1 \us03/U220  ( .A(\us03/n41 ), .B(\us03/n33 ), .Y(\us03/n272 ) );
  OAI221XL \us03/U219  ( .A0(sa03[1]), .A1(\us03/n247 ), .B0(\us03/n4 ), .B1(
        \us03/n189 ), .C0(\us03/n272 ), .Y(\us03/n279 ) );
  NAND2X1 \us03/U218  ( .A(sa03[2]), .B(\us03/n149 ), .Y(\us03/n276 ) );
  XNOR2X1 \us03/U217  ( .A(\us03/n129 ), .B(sa03[1]), .Y(\us03/n155 ) );
  MXI2X1 \us03/U216  ( .A(\us03/n276 ), .B(\us03/n277 ), .S0(\us03/n155 ), .Y(
        \us03/n275 ) );
  OAI22X1 \us03/U215  ( .A0(\us03/n273 ), .A1(\us03/n10 ), .B0(\us03/n274 ), 
        .B1(\us03/n52 ), .Y(\us03/n266 ) );
  NOR2X1 \us03/U214  ( .A(\us03/n20 ), .B(\us03/n226 ), .Y(\us03/n176 ) );
  OAI21XL \us03/U213  ( .A0(\us03/n4 ), .A1(\us03/n271 ), .B0(\us03/n272 ), 
        .Y(\us03/n270 ) );
  OAI31X1 \us03/U212  ( .A0(\us03/n176 ), .A1(\us03/n269 ), .A2(\us03/n270 ), 
        .B0(\us03/n16 ), .Y(\us03/n268 ) );
  INVX1 \us03/U211  ( .A(\us03/n268 ), .Y(\us03/n267 ) );
  AOI211X1 \us03/U210  ( .A0(\us03/n55 ), .A1(\us03/n265 ), .B0(\us03/n266 ), 
        .C0(\us03/n267 ), .Y(\us03/n264 ) );
  MXI2X1 \us03/U209  ( .A(\us03/n263 ), .B(\us03/n264 ), .S0(sa03[6]), .Y(
        sa03_sr[2]) );
  NOR2X1 \us03/U208  ( .A(\us03/n94 ), .B(sa03[1]), .Y(\us03/n211 ) );
  INVX1 \us03/U207  ( .A(\us03/n262 ), .Y(\us03/n261 ) );
  AOI211X1 \us03/U206  ( .A0(\us03/n259 ), .A1(\us03/n24 ), .B0(\us03/n260 ), 
        .C0(\us03/n261 ), .Y(\us03/n255 ) );
  OAI22X1 \us03/U205  ( .A0(\us03/n20 ), .A1(\us03/n68 ), .B0(\us03/n27 ), 
        .B1(\us03/n37 ), .Y(\us03/n257 ) );
  NOR3X1 \us03/U204  ( .A(\us03/n257 ), .B(\us03/n258 ), .C(\us03/n50 ), .Y(
        \us03/n256 ) );
  MXI2X1 \us03/U203  ( .A(\us03/n255 ), .B(\us03/n256 ), .S0(\us03/n252 ), .Y(
        \us03/n254 ) );
  AOI221X1 \us03/U202  ( .A0(\us03/n211 ), .A1(\us03/n5 ), .B0(\us03/n40 ), 
        .B1(sa03[4]), .C0(\us03/n254 ), .Y(\us03/n248 ) );
  INVX1 \us03/U201  ( .A(\us03/n211 ), .Y(\us03/n106 ) );
  NAND2X1 \us03/U200  ( .A(\us03/n200 ), .B(\us03/n106 ), .Y(\us03/n83 ) );
  NAND2X1 \us03/U199  ( .A(\us03/n199 ), .B(\us03/n204 ), .Y(\us03/n169 ) );
  AOI2BB2X1 \us03/U198  ( .B0(\us03/n65 ), .B1(\us03/n24 ), .A0N(\us03/n169 ), 
        .A1N(\us03/n20 ), .Y(\us03/n253 ) );
  OAI221XL \us03/U197  ( .A0(\us03/n172 ), .A1(\us03/n18 ), .B0(\us03/n27 ), 
        .B1(\us03/n83 ), .C0(\us03/n253 ), .Y(\us03/n251 ) );
  MXI2X1 \us03/U196  ( .A(\us03/n250 ), .B(\us03/n251 ), .S0(\us03/n252 ), .Y(
        \us03/n249 ) );
  MXI2X1 \us03/U195  ( .A(\us03/n248 ), .B(\us03/n249 ), .S0(\us03/n234 ), .Y(
        \us03/n228 ) );
  OAI21XL \us03/U194  ( .A0(\us03/n58 ), .A1(\us03/n27 ), .B0(\us03/n247 ), 
        .Y(\us03/n245 ) );
  NOR2X1 \us03/U193  ( .A(sa03[7]), .B(\us03/n145 ), .Y(\us03/n246 ) );
  XNOR2X1 \us03/U192  ( .A(\us03/n69 ), .B(sa03[1]), .Y(\us03/n130 ) );
  MXI2X1 \us03/U191  ( .A(\us03/n245 ), .B(\us03/n246 ), .S0(\us03/n130 ), .Y(
        \us03/n243 ) );
  OAI211X1 \us03/U190  ( .A0(\us03/n4 ), .A1(\us03/n149 ), .B0(\us03/n243 ), 
        .C0(\us03/n244 ), .Y(\us03/n230 ) );
  NOR2X1 \us03/U189  ( .A(\us03/n242 ), .B(\us03/n137 ), .Y(\us03/n70 ) );
  OAI221XL \us03/U188  ( .A0(\us03/n159 ), .A1(\us03/n27 ), .B0(\us03/n20 ), 
        .B1(\us03/n34 ), .C0(\us03/n241 ), .Y(\us03/n231 ) );
  NAND2X1 \us03/U187  ( .A(\us03/n101 ), .B(\us03/n240 ), .Y(\us03/n76 ) );
  AOI21X1 \us03/U186  ( .A0(\us03/n122 ), .A1(\us03/n106 ), .B0(\us03/n129 ), 
        .Y(\us03/n237 ) );
  INVX1 \us03/U185  ( .A(\us03/n239 ), .Y(\us03/n238 ) );
  OAI21XL \us03/U184  ( .A0(\us03/n237 ), .A1(\us03/n43 ), .B0(\us03/n238 ), 
        .Y(\us03/n236 ) );
  OAI221XL \us03/U183  ( .A0(\us03/n18 ), .A1(\us03/n76 ), .B0(\us03/n59 ), 
        .B1(\us03/n27 ), .C0(\us03/n236 ), .Y(\us03/n232 ) );
  AOI2BB2X1 \us03/U182  ( .B0(\us03/n24 ), .B1(\us03/n187 ), .A0N(\us03/n227 ), 
        .A1N(\us03/n20 ), .Y(\us03/n235 ) );
  OAI211X1 \us03/U181  ( .A0(\us03/n27 ), .A1(\us03/n122 ), .B0(\us03/n158 ), 
        .C0(\us03/n235 ), .Y(\us03/n233 ) );
  MX4X1 \us03/U180  ( .A(\us03/n230 ), .B(\us03/n231 ), .C(\us03/n232 ), .D(
        \us03/n233 ), .S0(\us03/n234 ), .S1(sa03[5]), .Y(\us03/n229 ) );
  MX2X1 \us03/U179  ( .A(\us03/n228 ), .B(\us03/n229 ), .S0(sa03[6]), .Y(
        sa03_sr[3]) );
  NOR2BX1 \us03/U178  ( .AN(\us03/n204 ), .B(\us03/n137 ), .Y(\us03/n110 ) );
  INVX1 \us03/U177  ( .A(\us03/n110 ), .Y(\us03/n64 ) );
  AOI22X1 \us03/U176  ( .A0(\us03/n225 ), .A1(\us03/n226 ), .B0(\us03/n6 ), 
        .B1(\us03/n227 ), .Y(\us03/n224 ) );
  OAI221XL \us03/U175  ( .A0(\us03/n27 ), .A1(\us03/n64 ), .B0(\us03/n4 ), 
        .B1(\us03/n83 ), .C0(\us03/n224 ), .Y(\us03/n212 ) );
  NAND2X1 \us03/U174  ( .A(\us03/n34 ), .B(\us03/n204 ), .Y(\us03/n221 ) );
  OAI21XL \us03/U173  ( .A0(\us03/n69 ), .A1(\us03/n223 ), .B0(\us03/n27 ), 
        .Y(\us03/n222 ) );
  NOR2X1 \us03/U172  ( .A(\us03/n217 ), .B(\us03/n42 ), .Y(\us03/n208 ) );
  AOI211X1 \us03/U171  ( .A0(\us03/n208 ), .A1(\us03/n5 ), .B0(\us03/n220 ), 
        .C0(\us03/n173 ), .Y(\us03/n219 ) );
  OAI22X1 \us03/U170  ( .A0(\us03/n218 ), .A1(\us03/n10 ), .B0(\us03/n219 ), 
        .B1(\us03/n114 ), .Y(\us03/n213 ) );
  INVX1 \us03/U169  ( .A(\us03/n135 ), .Y(\us03/n215 ) );
  NOR2X1 \us03/U168  ( .A(\us03/n4 ), .B(\us03/n159 ), .Y(\us03/n31 ) );
  INVX1 \us03/U167  ( .A(\us03/n31 ), .Y(\us03/n196 ) );
  AOI31X1 \us03/U166  ( .A0(\us03/n215 ), .A1(\us03/n196 ), .A2(\us03/n216 ), 
        .B0(\us03/n52 ), .Y(\us03/n214 ) );
  AOI211X1 \us03/U165  ( .A0(\us03/n55 ), .A1(\us03/n212 ), .B0(\us03/n213 ), 
        .C0(\us03/n214 ), .Y(\us03/n190 ) );
  INVX1 \us03/U164  ( .A(\us03/n207 ), .Y(\us03/n192 ) );
  NOR2X1 \us03/U163  ( .A(\us03/n25 ), .B(\us03/n98 ), .Y(\us03/n32 ) );
  OAI22X1 \us03/U162  ( .A0(\us03/n28 ), .A1(\us03/n4 ), .B0(\us03/n188 ), 
        .B1(\us03/n27 ), .Y(\us03/n206 ) );
  NAND2X1 \us03/U161  ( .A(\us03/n204 ), .B(\us03/n80 ), .Y(\us03/n118 ) );
  INVX1 \us03/U160  ( .A(\us03/n118 ), .Y(\us03/n123 ) );
  NAND2X1 \us03/U159  ( .A(\us03/n94 ), .B(\us03/n79 ), .Y(\us03/n203 ) );
  OAI2BB1X1 \us03/U158  ( .A0N(\us03/n199 ), .A1N(\us03/n200 ), .B0(\us03/n33 ), .Y(\us03/n195 ) );
  INVX1 \us03/U157  ( .A(\us03/n55 ), .Y(\us03/n12 ) );
  AOI31X1 \us03/U156  ( .A0(\us03/n195 ), .A1(\us03/n196 ), .A2(\us03/n197 ), 
        .B0(\us03/n12 ), .Y(\us03/n194 ) );
  AOI211X1 \us03/U155  ( .A0(\us03/n89 ), .A1(\us03/n192 ), .B0(\us03/n193 ), 
        .C0(\us03/n194 ), .Y(\us03/n191 ) );
  MXI2X1 \us03/U154  ( .A(\us03/n190 ), .B(\us03/n191 ), .S0(sa03[6]), .Y(
        sa03_sr[4]) );
  OAI21XL \us03/U153  ( .A0(\us03/n69 ), .A1(\us03/n189 ), .B0(\us03/n27 ), 
        .Y(\us03/n186 ) );
  INVX1 \us03/U152  ( .A(\us03/n183 ), .Y(\us03/n180 ) );
  NAND2X1 \us03/U151  ( .A(\us03/n74 ), .B(\us03/n182 ), .Y(\us03/n181 ) );
  AOI211X1 \us03/U150  ( .A0(\us03/n179 ), .A1(\us03/n24 ), .B0(\us03/n180 ), 
        .C0(\us03/n181 ), .Y(\us03/n165 ) );
  INVX1 \us03/U149  ( .A(\us03/n178 ), .Y(\us03/n175 ) );
  AOI211X1 \us03/U148  ( .A0(\us03/n175 ), .A1(\us03/n5 ), .B0(\us03/n176 ), 
        .C0(\us03/n177 ), .Y(\us03/n174 ) );
  OAI221XL \us03/U147  ( .A0(\us03/n159 ), .A1(\us03/n27 ), .B0(\us03/n145 ), 
        .B1(\us03/n20 ), .C0(\us03/n174 ), .Y(\us03/n167 ) );
  MXI2X1 \us03/U146  ( .A(\us03/n40 ), .B(\us03/n173 ), .S0(\us03/n96 ), .Y(
        \us03/n170 ) );
  AOI22X1 \us03/U145  ( .A0(\us03/n137 ), .A1(\us03/n24 ), .B0(\us03/n172 ), 
        .B1(\us03/n6 ), .Y(\us03/n171 ) );
  OAI211X1 \us03/U144  ( .A0(\us03/n20 ), .A1(\us03/n169 ), .B0(\us03/n170 ), 
        .C0(\us03/n171 ), .Y(\us03/n168 ) );
  AOI22X1 \us03/U143  ( .A0(\us03/n89 ), .A1(\us03/n167 ), .B0(\us03/n55 ), 
        .B1(\us03/n168 ), .Y(\us03/n166 ) );
  OAI221XL \us03/U142  ( .A0(\us03/n164 ), .A1(\us03/n114 ), .B0(\us03/n165 ), 
        .B1(\us03/n52 ), .C0(\us03/n166 ), .Y(\us03/n138 ) );
  OAI21XL \us03/U141  ( .A0(\us03/n41 ), .A1(\us03/n163 ), .B0(\us03/n69 ), 
        .Y(\us03/n162 ) );
  AOI221X1 \us03/U140  ( .A0(\us03/n159 ), .A1(\us03/n24 ), .B0(\us03/n160 ), 
        .B1(\us03/n33 ), .C0(\us03/n161 ), .Y(\us03/n140 ) );
  OAI21XL \us03/U139  ( .A0(\us03/n157 ), .A1(\us03/n20 ), .B0(\us03/n158 ), 
        .Y(\us03/n156 ) );
  NOR2X1 \us03/U138  ( .A(\us03/n4 ), .B(\us03/n136 ), .Y(\us03/n153 ) );
  NOR2X1 \us03/U137  ( .A(\us03/n145 ), .B(\us03/n69 ), .Y(\us03/n154 ) );
  MXI2X1 \us03/U136  ( .A(\us03/n153 ), .B(\us03/n154 ), .S0(\us03/n155 ), .Y(
        \us03/n152 ) );
  OAI221XL \us03/U135  ( .A0(\us03/n110 ), .A1(\us03/n18 ), .B0(\us03/n20 ), 
        .B1(\us03/n151 ), .C0(\us03/n152 ), .Y(\us03/n143 ) );
  AOI21X1 \us03/U134  ( .A0(\us03/n149 ), .A1(\us03/n150 ), .B0(\us03/n18 ), 
        .Y(\us03/n148 ) );
  AOI2BB1X1 \us03/U133  ( .A0N(\us03/n147 ), .A1N(\us03/n27 ), .B0(\us03/n148 ), .Y(\us03/n146 ) );
  OAI221XL \us03/U132  ( .A0(\us03/n145 ), .A1(\us03/n20 ), .B0(\us03/n4 ), 
        .B1(\us03/n34 ), .C0(\us03/n146 ), .Y(\us03/n144 ) );
  AOI22X1 \us03/U131  ( .A0(\us03/n89 ), .A1(\us03/n143 ), .B0(\us03/n14 ), 
        .B1(\us03/n144 ), .Y(\us03/n142 ) );
  OAI221XL \us03/U130  ( .A0(\us03/n140 ), .A1(\us03/n12 ), .B0(\us03/n141 ), 
        .B1(\us03/n114 ), .C0(\us03/n142 ), .Y(\us03/n139 ) );
  MX2X1 \us03/U129  ( .A(\us03/n138 ), .B(\us03/n139 ), .S0(sa03[6]), .Y(
        sa03_sr[5]) );
  INVX1 \us03/U128  ( .A(\us03/n70 ), .Y(\us03/n133 ) );
  OAI22X1 \us03/U127  ( .A0(\us03/n4 ), .A1(\us03/n136 ), .B0(\us03/n137 ), 
        .B1(\us03/n27 ), .Y(\us03/n134 ) );
  AOI211X1 \us03/U126  ( .A0(\us03/n133 ), .A1(\us03/n69 ), .B0(\us03/n134 ), 
        .C0(\us03/n135 ), .Y(\us03/n112 ) );
  INVX1 \us03/U125  ( .A(\us03/n132 ), .Y(\us03/n131 ) );
  OAI21XL \us03/U124  ( .A0(\us03/n18 ), .A1(\us03/n37 ), .B0(\us03/n128 ), 
        .Y(\us03/n127 ) );
  OAI221XL \us03/U123  ( .A0(\us03/n18 ), .A1(\us03/n105 ), .B0(\us03/n123 ), 
        .B1(\us03/n27 ), .C0(\us03/n124 ), .Y(\us03/n116 ) );
  NAND2X1 \us03/U122  ( .A(\us03/n121 ), .B(\us03/n122 ), .Y(\us03/n30 ) );
  OAI221XL \us03/U121  ( .A0(\us03/n18 ), .A1(\us03/n118 ), .B0(\us03/n27 ), 
        .B1(\us03/n30 ), .C0(\us03/n119 ), .Y(\us03/n117 ) );
  AOI22X1 \us03/U120  ( .A0(\us03/n89 ), .A1(\us03/n116 ), .B0(\us03/n55 ), 
        .B1(\us03/n117 ), .Y(\us03/n115 ) );
  OAI221XL \us03/U119  ( .A0(\us03/n112 ), .A1(\us03/n52 ), .B0(\us03/n113 ), 
        .B1(\us03/n114 ), .C0(\us03/n115 ), .Y(\us03/n84 ) );
  OAI22X1 \us03/U118  ( .A0(\us03/n110 ), .A1(\us03/n4 ), .B0(\us03/n20 ), 
        .B1(\us03/n21 ), .Y(\us03/n108 ) );
  AOI21X1 \us03/U117  ( .A0(sa03[1]), .A1(\us03/n58 ), .B0(\us03/n27 ), .Y(
        \us03/n109 ) );
  AOI211X1 \us03/U116  ( .A0(\us03/n5 ), .A1(\us03/n107 ), .B0(\us03/n108 ), 
        .C0(\us03/n109 ), .Y(\us03/n86 ) );
  OAI22X1 \us03/U115  ( .A0(\us03/n45 ), .A1(\us03/n4 ), .B0(sa03[4]), .B1(
        \us03/n18 ), .Y(\us03/n103 ) );
  AOI21X1 \us03/U114  ( .A0(\us03/n105 ), .A1(\us03/n106 ), .B0(\us03/n20 ), 
        .Y(\us03/n104 ) );
  AOI211X1 \us03/U113  ( .A0(\us03/n33 ), .A1(\us03/n102 ), .B0(\us03/n103 ), 
        .C0(\us03/n104 ), .Y(\us03/n87 ) );
  NAND2X1 \us03/U112  ( .A(\us03/n100 ), .B(\us03/n101 ), .Y(\us03/n62 ) );
  OAI221XL \us03/U111  ( .A0(\us03/n27 ), .A1(\us03/n62 ), .B0(\us03/n4 ), 
        .B1(\us03/n21 ), .C0(\us03/n97 ), .Y(\us03/n90 ) );
  NOR3X1 \us03/U110  ( .A(\us03/n4 ), .B(\us03/n95 ), .C(\us03/n96 ), .Y(
        \us03/n67 ) );
  AOI31X1 \us03/U109  ( .A0(\us03/n79 ), .A1(\us03/n94 ), .A2(\us03/n6 ), .B0(
        \us03/n67 ), .Y(\us03/n93 ) );
  OAI221XL \us03/U108  ( .A0(\us03/n73 ), .A1(\us03/n27 ), .B0(\us03/n92 ), 
        .B1(\us03/n20 ), .C0(\us03/n93 ), .Y(\us03/n91 ) );
  AOI22X1 \us03/U107  ( .A0(\us03/n89 ), .A1(\us03/n90 ), .B0(\us03/n16 ), 
        .B1(\us03/n91 ), .Y(\us03/n88 ) );
  OAI221XL \us03/U106  ( .A0(\us03/n86 ), .A1(\us03/n52 ), .B0(\us03/n87 ), 
        .B1(\us03/n12 ), .C0(\us03/n88 ), .Y(\us03/n85 ) );
  MX2X1 \us03/U105  ( .A(\us03/n84 ), .B(\us03/n85 ), .S0(sa03[6]), .Y(
        sa03_sr[6]) );
  INVX1 \us03/U104  ( .A(\us03/n81 ), .Y(\us03/n77 ) );
  AOI21X1 \us03/U103  ( .A0(\us03/n79 ), .A1(\us03/n80 ), .B0(\us03/n27 ), .Y(
        \us03/n78 ) );
  AOI211X1 \us03/U102  ( .A0(\us03/n5 ), .A1(\us03/n76 ), .B0(\us03/n77 ), 
        .C0(\us03/n78 ), .Y(\us03/n51 ) );
  OAI211X1 \us03/U101  ( .A0(\us03/n73 ), .A1(\us03/n27 ), .B0(\us03/n74 ), 
        .C0(\us03/n75 ), .Y(\us03/n72 ) );
  AOI21X1 \us03/U100  ( .A0(\us03/n68 ), .A1(\us03/n69 ), .B0(\us03/n6 ), .Y(
        \us03/n63 ) );
  INVX1 \us03/U99  ( .A(\us03/n67 ), .Y(\us03/n66 ) );
  OAI221XL \us03/U98  ( .A0(\us03/n63 ), .A1(\us03/n64 ), .B0(\us03/n65 ), 
        .B1(\us03/n27 ), .C0(\us03/n66 ), .Y(\us03/n56 ) );
  AOI2BB2X1 \us03/U97  ( .B0(\us03/n61 ), .B1(\us03/n24 ), .A0N(\us03/n62 ), 
        .A1N(\us03/n20 ), .Y(\us03/n60 ) );
  OAI221XL \us03/U96  ( .A0(\us03/n58 ), .A1(\us03/n18 ), .B0(\us03/n59 ), 
        .B1(\us03/n27 ), .C0(\us03/n60 ), .Y(\us03/n57 ) );
  AOI22X1 \us03/U95  ( .A0(\us03/n55 ), .A1(\us03/n56 ), .B0(\us03/n16 ), .B1(
        \us03/n57 ), .Y(\us03/n54 ) );
  OAI221XL \us03/U94  ( .A0(\us03/n51 ), .A1(\us03/n52 ), .B0(\us03/n53 ), 
        .B1(\us03/n10 ), .C0(\us03/n54 ), .Y(\us03/n7 ) );
  INVX1 \us03/U93  ( .A(\us03/n50 ), .Y(\us03/n49 ) );
  OAI221XL \us03/U92  ( .A0(\us03/n47 ), .A1(\us03/n18 ), .B0(\us03/n27 ), 
        .B1(\us03/n48 ), .C0(\us03/n49 ), .Y(\us03/n46 ) );
  NOR2X1 \us03/U91  ( .A(\us03/n41 ), .B(\us03/n42 ), .Y(\us03/n38 ) );
  INVX1 \us03/U90  ( .A(\us03/n40 ), .Y(\us03/n39 ) );
  INVX1 \us03/U89  ( .A(\us03/n32 ), .Y(\us03/n26 ) );
  AOI21X1 \us03/U88  ( .A0(\us03/n5 ), .A1(\us03/n30 ), .B0(\us03/n31 ), .Y(
        \us03/n29 ) );
  OAI221XL \us03/U87  ( .A0(\us03/n26 ), .A1(\us03/n27 ), .B0(\us03/n28 ), 
        .B1(\us03/n20 ), .C0(\us03/n29 ), .Y(\us03/n15 ) );
  OAI221XL \us03/U86  ( .A0(\us03/n18 ), .A1(\us03/n19 ), .B0(\us03/n20 ), 
        .B1(\us03/n21 ), .C0(\us03/n22 ), .Y(\us03/n17 ) );
  AOI22X1 \us03/U85  ( .A0(\us03/n14 ), .A1(\us03/n15 ), .B0(\us03/n16 ), .B1(
        \us03/n17 ), .Y(\us03/n13 ) );
  OAI221XL \us03/U84  ( .A0(\us03/n9 ), .A1(\us03/n10 ), .B0(\us03/n11 ), .B1(
        \us03/n12 ), .C0(\us03/n13 ), .Y(\us03/n8 ) );
  MX2X1 \us03/U83  ( .A(\us03/n7 ), .B(\us03/n8 ), .S0(sa03[6]), .Y(sa03_sr[7]) );
  NOR2X4 \us03/U82  ( .A(\us03/n129 ), .B(sa03[2]), .Y(\us03/n43 ) );
  CLKINVX3 \us03/U81  ( .A(\us03/n14 ), .Y(\us03/n52 ) );
  OAI22XL \us03/U80  ( .A0(\us03/n201 ), .A1(\us03/n52 ), .B0(\us03/n202 ), 
        .B1(\us03/n114 ), .Y(\us03/n193 ) );
  CLKINVX3 \us03/U79  ( .A(sa03[5]), .Y(\us03/n252 ) );
  NOR2X2 \us03/U78  ( .A(\us03/n252 ), .B(\us03/n234 ), .Y(\us03/n55 ) );
  CLKINVX3 \us03/U77  ( .A(sa03[7]), .Y(\us03/n129 ) );
  NOR2X4 \us03/U76  ( .A(\us03/n129 ), .B(\us03/n69 ), .Y(\us03/n24 ) );
  AOI22XL \us03/U75  ( .A0(\us03/n70 ), .A1(\us03/n24 ), .B0(\us03/n96 ), .B1(
        \us03/n129 ), .Y(\us03/n241 ) );
  NOR2X2 \us03/U74  ( .A(\us03/n252 ), .B(sa03[0]), .Y(\us03/n89 ) );
  CLKINVX3 \us03/U73  ( .A(sa03[0]), .Y(\us03/n234 ) );
  NOR2X4 \us03/U72  ( .A(\us03/n69 ), .B(sa03[7]), .Y(\us03/n33 ) );
  INVX12 \us03/U71  ( .A(\us03/n33 ), .Y(\us03/n27 ) );
  CLKINVX3 \us03/U70  ( .A(\us03/n1 ), .Y(\us03/n6 ) );
  CLKINVX3 \us03/U69  ( .A(\us03/n1 ), .Y(\us03/n5 ) );
  INVXL \us03/U68  ( .A(\us03/n24 ), .Y(\us03/n36 ) );
  INVX4 \us03/U67  ( .A(\us03/n3 ), .Y(\us03/n4 ) );
  INVXL \us03/U66  ( .A(\us03/n36 ), .Y(\us03/n3 ) );
  INVX4 \us03/U65  ( .A(sa03[1]), .Y(\us03/n226 ) );
  INVX4 \us03/U64  ( .A(\us03/n43 ), .Y(\us03/n20 ) );
  AOI221X4 \us03/U63  ( .A0(\us03/n24 ), .A1(\us03/n82 ), .B0(\us03/n43 ), 
        .B1(\us03/n295 ), .C0(\us03/n173 ), .Y(\us03/n346 ) );
  AOI221X4 \us03/U62  ( .A0(\us03/n5 ), .A1(\us03/n96 ), .B0(\us03/n43 ), .B1(
        \us03/n239 ), .C0(\us03/n340 ), .Y(\us03/n336 ) );
  AOI222X4 \us03/U61  ( .A0(\us03/n59 ), .A1(\us03/n43 ), .B0(\us03/n6 ), .B1(
        \us03/n221 ), .C0(\us03/n222 ), .C1(\us03/n187 ), .Y(\us03/n218 ) );
  AOI222X4 \us03/U60  ( .A0(\us03/n123 ), .A1(\us03/n43 ), .B0(sa03[2]), .B1(
        \us03/n203 ), .C0(\us03/n6 ), .C1(\us03/n71 ), .Y(\us03/n202 ) );
  AOI221X4 \us03/U59  ( .A0(\us03/n314 ), .A1(\us03/n43 ), .B0(\us03/n160 ), 
        .B1(\us03/n24 ), .C0(\us03/n315 ), .Y(\us03/n307 ) );
  AOI221X4 \us03/U58  ( .A0(\us03/n43 ), .A1(\us03/n208 ), .B0(\us03/n76 ), 
        .B1(\us03/n24 ), .C0(\us03/n209 ), .Y(\us03/n207 ) );
  AOI221X4 \us03/U57  ( .A0(\us03/n43 ), .A1(\us03/n205 ), .B0(\us03/n32 ), 
        .B1(\us03/n6 ), .C0(\us03/n206 ), .Y(\us03/n201 ) );
  AOI221X4 \us03/U56  ( .A0(\us03/n43 ), .A1(\us03/n44 ), .B0(\us03/n45 ), 
        .B1(\us03/n24 ), .C0(\us03/n46 ), .Y(\us03/n9 ) );
  AOI22XL \us03/U55  ( .A0(\us03/n217 ), .A1(\us03/n43 ), .B0(\us03/n33 ), 
        .B1(\us03/n47 ), .Y(\us03/n216 ) );
  AOI22XL \us03/U54  ( .A0(\us03/n98 ), .A1(\us03/n43 ), .B0(\us03/n6 ), .B1(
        \us03/n99 ), .Y(\us03/n97 ) );
  AOI22XL \us03/U53  ( .A0(\us03/n82 ), .A1(\us03/n43 ), .B0(\us03/n83 ), .B1(
        \us03/n24 ), .Y(\us03/n81 ) );
  AOI2BB2XL \us03/U52  ( .B0(\us03/n43 ), .B1(\us03/n94 ), .A0N(\us03/n120 ), 
        .A1N(\us03/n4 ), .Y(\us03/n119 ) );
  AOI222X4 \us03/U51  ( .A0(\us03/n125 ), .A1(\us03/n33 ), .B0(\us03/n145 ), 
        .B1(\us03/n40 ), .C0(\us03/n43 ), .C1(\us03/n184 ), .Y(\us03/n183 ) );
  AOI22XL \us03/U50  ( .A0(\us03/n43 ), .A1(\us03/n303 ), .B0(\us03/n24 ), 
        .B1(\us03/n96 ), .Y(\us03/n358 ) );
  AOI22XL \us03/U49  ( .A0(\us03/n43 ), .A1(\us03/n100 ), .B0(\us03/n24 ), 
        .B1(\us03/n125 ), .Y(\us03/n124 ) );
  AOI21XL \us03/U48  ( .A0(\us03/n159 ), .A1(\us03/n43 ), .B0(\us03/n40 ), .Y(
        \us03/n262 ) );
  AOI22XL \us03/U47  ( .A0(\us03/n40 ), .A1(\us03/n94 ), .B0(\us03/n43 ), .B1(
        \us03/n187 ), .Y(\us03/n244 ) );
  AOI22XL \us03/U46  ( .A0(\us03/n184 ), .A1(\us03/n5 ), .B0(\us03/n198 ), 
        .B1(\us03/n43 ), .Y(\us03/n197 ) );
  NOR2XL \us03/U45  ( .A(\us03/n33 ), .B(\us03/n2 ), .Y(\us03/n302 ) );
  MXI2XL \us03/U44  ( .A(\us03/n2 ), .B(\us03/n6 ), .S0(\us03/n28 ), .Y(
        \us03/n311 ) );
  INVXL \us03/U43  ( .A(\us03/n20 ), .Y(\us03/n2 ) );
  INVX4 \us03/U42  ( .A(\us03/n6 ), .Y(\us03/n18 ) );
  AOI21XL \us03/U41  ( .A0(\us03/n18 ), .A1(\us03/n162 ), .B0(\us03/n25 ), .Y(
        \us03/n161 ) );
  INVX4 \us03/U40  ( .A(sa03[2]), .Y(\us03/n69 ) );
  NOR2X4 \us03/U39  ( .A(\us03/n226 ), .B(\us03/n4 ), .Y(\us03/n40 ) );
  CLKINVX3 \us03/U38  ( .A(sa03[3]), .Y(\us03/n136 ) );
  NOR2X2 \us03/U37  ( .A(\us03/n136 ), .B(sa03[4]), .Y(\us03/n145 ) );
  CLKINVX3 \us03/U36  ( .A(sa03[4]), .Y(\us03/n58 ) );
  NOR2X2 \us03/U35  ( .A(\us03/n58 ), .B(sa03[3]), .Y(\us03/n159 ) );
  NOR2X2 \us03/U34  ( .A(\us03/n136 ), .B(\us03/n58 ), .Y(\us03/n259 ) );
  NOR2X2 \us03/U33  ( .A(sa03[4]), .B(sa03[3]), .Y(\us03/n278 ) );
  NOR2X2 \us03/U32  ( .A(\us03/n259 ), .B(\us03/n278 ), .Y(\us03/n47 ) );
  CLKINVX3 \us03/U31  ( .A(\us03/n259 ), .Y(\us03/n44 ) );
  NOR2X2 \us03/U30  ( .A(\us03/n44 ), .B(sa03[1]), .Y(\us03/n137 ) );
  AOI21XL \us03/U29  ( .A0(\us03/n44 ), .A1(\us03/n111 ), .B0(\us03/n4 ), .Y(
        \us03/n177 ) );
  AOI22XL \us03/U28  ( .A0(\us03/n23 ), .A1(\us03/n24 ), .B0(\us03/n25 ), .B1(
        sa03[2]), .Y(\us03/n22 ) );
  AOI22XL \us03/U27  ( .A0(\us03/n33 ), .A1(sa03[3]), .B0(\us03/n24 ), .B1(
        \us03/n58 ), .Y(\us03/n277 ) );
  NAND2XL \us03/U26  ( .A(\us03/n198 ), .B(\us03/n24 ), .Y(\us03/n132 ) );
  OAI2BB2XL \us03/U25  ( .B0(\us03/n20 ), .B1(\us03/n111 ), .A0N(\us03/n125 ), 
        .A1N(\us03/n24 ), .Y(\us03/n220 ) );
  NAND2XL \us03/U24  ( .A(\us03/n111 ), .B(\us03/n101 ), .Y(\us03/n21 ) );
  NAND2XL \us03/U23  ( .A(\us03/n111 ), .B(\us03/n300 ), .Y(\us03/n187 ) );
  NAND2XL \us03/U22  ( .A(\us03/n111 ), .B(\us03/n121 ), .Y(\us03/n303 ) );
  AOI221XL \us03/U21  ( .A0(\us03/n43 ), .A1(\us03/n151 ), .B0(\us03/n25 ), 
        .B1(\us03/n69 ), .C0(\us03/n275 ), .Y(\us03/n274 ) );
  NOR2BXL \us03/U20  ( .AN(\us03/n101 ), .B(\us03/n25 ), .Y(\us03/n172 ) );
  NAND2X2 \us03/U19  ( .A(\us03/n58 ), .B(\us03/n226 ), .Y(\us03/n34 ) );
  OAI222X1 \us03/U18  ( .A0(\us03/n27 ), .A1(\us03/n34 ), .B0(\us03/n69 ), 
        .B1(\us03/n205 ), .C0(\us03/n20 ), .C1(\us03/n79 ), .Y(\us03/n260 ) );
  OAI222X1 \us03/U17  ( .A0(\us03/n20 ), .A1(\us03/n99 ), .B0(\us03/n27 ), 
        .B1(\us03/n101 ), .C0(\us03/n184 ), .C1(\us03/n4 ), .Y(\us03/n250 ) );
  OAI222X1 \us03/U16  ( .A0(\us03/n4 ), .A1(\us03/n37 ), .B0(\us03/n38 ), .B1(
        \us03/n20 ), .C0(sa03[4]), .C1(\us03/n39 ), .Y(\us03/n35 ) );
  AOI221X1 \us03/U15  ( .A0(\us03/n5 ), .A1(\us03/n19 ), .B0(\us03/n33 ), .B1(
        \us03/n34 ), .C0(\us03/n35 ), .Y(\us03/n11 ) );
  OR2X2 \us03/U14  ( .A(sa03[2]), .B(sa03[7]), .Y(\us03/n1 ) );
  AOI221XL \us03/U13  ( .A0(\us03/n70 ), .A1(\us03/n43 ), .B0(\us03/n24 ), 
        .B1(\us03/n71 ), .C0(\us03/n72 ), .Y(\us03/n53 ) );
  AOI221XL \us03/U12  ( .A0(\us03/n59 ), .A1(\us03/n33 ), .B0(\us03/n43 ), 
        .B1(\us03/n126 ), .C0(\us03/n127 ), .Y(\us03/n113 ) );
  AOI222XL \us03/U11  ( .A0(\us03/n185 ), .A1(\us03/n43 ), .B0(\us03/n186 ), 
        .B1(\us03/n187 ), .C0(\us03/n6 ), .C1(\us03/n188 ), .Y(\us03/n164 ) );
  AOI221X1 \us03/U10  ( .A0(\us03/n313 ), .A1(\us03/n5 ), .B0(\us03/n23 ), 
        .B1(\us03/n2 ), .C0(\us03/n328 ), .Y(\us03/n320 ) );
  AOI221X1 \us03/U9  ( .A0(\us03/n40 ), .A1(\us03/n136 ), .B0(\us03/n33 ), 
        .B1(\us03/n178 ), .C0(\us03/n338 ), .Y(\us03/n337 ) );
  AOI222XL \us03/U8  ( .A0(\us03/n278 ), .A1(\us03/n24 ), .B0(\us03/n42 ), 
        .B1(\us03/n33 ), .C0(\us03/n43 ), .C1(\us03/n136 ), .Y(\us03/n351 ) );
  AOI31X1 \us03/U7  ( .A0(sa03[2]), .A1(\us03/n58 ), .A2(sa03[1]), .B0(
        \us03/n40 ), .Y(\us03/n350 ) );
  AOI31X1 \us03/U6  ( .A0(\us03/n44 ), .A1(\us03/n129 ), .A2(\us03/n130 ), 
        .B0(\us03/n131 ), .Y(\us03/n128 ) );
  AOI221X1 \us03/U5  ( .A0(\us03/n40 ), .A1(\us03/n136 ), .B0(\us03/n33 ), 
        .B1(\us03/n47 ), .C0(\us03/n156 ), .Y(\us03/n141 ) );
  OAI32X1 \us03/U4  ( .A0(\us03/n210 ), .A1(\us03/n145 ), .A2(\us03/n18 ), 
        .B0(\us03/n27 ), .B1(\us03/n211 ), .Y(\us03/n209 ) );
  AOI221X1 \us03/U3  ( .A0(\us03/n278 ), .A1(\us03/n40 ), .B0(\us03/n185 ), 
        .B1(\us03/n2 ), .C0(\us03/n279 ), .Y(\us03/n273 ) );
  OAI32X1 \us03/U2  ( .A0(\us03/n18 ), .A1(sa03[1]), .A2(\us03/n159 ), .B0(
        sa03[4]), .B1(\us03/n182 ), .Y(\us03/n318 ) );
  AOI31XL \us03/U1  ( .A0(\us03/n79 ), .A1(\us03/n44 ), .A2(\us03/n2 ), .B0(
        \us03/n280 ), .Y(\us03/n339 ) );
  NAND2X1 \us10/U366  ( .A(\us10/n47 ), .B(\us10/n226 ), .Y(\us10/n189 ) );
  NOR2X1 \us10/U365  ( .A(\us10/n226 ), .B(sa10[3]), .Y(\us10/n242 ) );
  INVX1 \us10/U364  ( .A(\us10/n242 ), .Y(\us10/n205 ) );
  AND2X1 \us10/U363  ( .A(\us10/n189 ), .B(\us10/n205 ), .Y(\us10/n65 ) );
  NOR2X1 \us10/U362  ( .A(\us10/n226 ), .B(\us10/n47 ), .Y(\us10/n45 ) );
  NOR2X1 \us10/U361  ( .A(\us10/n259 ), .B(\us10/n45 ), .Y(\us10/n73 ) );
  NAND2BX1 \us10/U360  ( .AN(\us10/n73 ), .B(\us10/n6 ), .Y(\us10/n158 ) );
  NOR2X1 \us10/U359  ( .A(\us10/n226 ), .B(\us10/n159 ), .Y(\us10/n95 ) );
  INVX1 \us10/U358  ( .A(\us10/n95 ), .Y(\us10/n111 ) );
  NOR2X1 \us10/U357  ( .A(\us10/n145 ), .B(sa10[1]), .Y(\us10/n42 ) );
  INVX1 \us10/U356  ( .A(\us10/n42 ), .Y(\us10/n121 ) );
  INVX1 \us10/U355  ( .A(\us10/n47 ), .Y(\us10/n96 ) );
  OAI211X1 \us10/U354  ( .A0(\us10/n65 ), .A1(\us10/n27 ), .B0(\us10/n158 ), 
        .C0(\us10/n358 ), .Y(\us10/n355 ) );
  NOR2X1 \us10/U353  ( .A(\us10/n226 ), .B(\us10/n145 ), .Y(\us10/n59 ) );
  NOR2X1 \us10/U352  ( .A(\us10/n96 ), .B(\us10/n59 ), .Y(\us10/n271 ) );
  NOR2X1 \us10/U351  ( .A(\us10/n226 ), .B(\us10/n278 ), .Y(\us10/n217 ) );
  INVX1 \us10/U350  ( .A(\us10/n217 ), .Y(\us10/n150 ) );
  NAND2X1 \us10/U349  ( .A(\us10/n44 ), .B(\us10/n150 ), .Y(\us10/n147 ) );
  NAND2X1 \us10/U348  ( .A(sa10[4]), .B(\us10/n226 ), .Y(\us10/n101 ) );
  INVX1 \us10/U347  ( .A(\us10/n159 ), .Y(\us10/n188 ) );
  NOR2X1 \us10/U346  ( .A(\us10/n188 ), .B(\us10/n226 ), .Y(\us10/n25 ) );
  INVX1 \us10/U345  ( .A(\us10/n172 ), .Y(\us10/n107 ) );
  AOI22X1 \us10/U344  ( .A0(\us10/n33 ), .A1(\us10/n147 ), .B0(\us10/n24 ), 
        .B1(\us10/n107 ), .Y(\us10/n357 ) );
  OAI221XL \us10/U343  ( .A0(\us10/n18 ), .A1(\us10/n121 ), .B0(\us10/n271 ), 
        .B1(\us10/n20 ), .C0(\us10/n357 ), .Y(\us10/n356 ) );
  MXI2X1 \us10/U342  ( .A(\us10/n355 ), .B(\us10/n356 ), .S0(\us10/n252 ), .Y(
        \us10/n331 ) );
  INVX1 \us10/U341  ( .A(\us10/n59 ), .Y(\us10/n79 ) );
  AND2X1 \us10/U340  ( .A(\us10/n101 ), .B(\us10/n79 ), .Y(\us10/n325 ) );
  XNOR2X1 \us10/U339  ( .A(sa10[5]), .B(\us10/n226 ), .Y(\us10/n352 ) );
  NOR2X1 \us10/U338  ( .A(\us10/n226 ), .B(\us10/n136 ), .Y(\us10/n281 ) );
  INVX1 \us10/U337  ( .A(\us10/n281 ), .Y(\us10/n19 ) );
  NAND2X1 \us10/U336  ( .A(\us10/n145 ), .B(\us10/n226 ), .Y(\us10/n223 ) );
  AOI21X1 \us10/U335  ( .A0(\us10/n19 ), .A1(\us10/n223 ), .B0(\us10/n27 ), 
        .Y(\us10/n354 ) );
  AOI31X1 \us10/U334  ( .A0(\us10/n6 ), .A1(\us10/n352 ), .A2(\us10/n259 ), 
        .B0(\us10/n354 ), .Y(\us10/n353 ) );
  OAI221XL \us10/U333  ( .A0(\us10/n20 ), .A1(\us10/n34 ), .B0(\us10/n325 ), 
        .B1(\us10/n4 ), .C0(\us10/n353 ), .Y(\us10/n347 ) );
  INVX1 \us10/U332  ( .A(\us10/n352 ), .Y(\us10/n349 ) );
  NAND2X1 \us10/U331  ( .A(\us10/n278 ), .B(\us10/n6 ), .Y(\us10/n74 ) );
  OAI211X1 \us10/U330  ( .A0(\us10/n349 ), .A1(\us10/n74 ), .B0(\us10/n350 ), 
        .C0(\us10/n351 ), .Y(\us10/n348 ) );
  MXI2X1 \us10/U329  ( .A(\us10/n347 ), .B(\us10/n348 ), .S0(\us10/n252 ), .Y(
        \us10/n332 ) );
  NOR2X1 \us10/U328  ( .A(\us10/n44 ), .B(\us10/n226 ), .Y(\us10/n157 ) );
  INVX1 \us10/U327  ( .A(\us10/n157 ), .Y(\us10/n240 ) );
  NAND2X1 \us10/U326  ( .A(\us10/n240 ), .B(\us10/n189 ), .Y(\us10/n68 ) );
  NOR2X1 \us10/U325  ( .A(\us10/n20 ), .B(\us10/n159 ), .Y(\us10/n225 ) );
  NOR2X1 \us10/U324  ( .A(\us10/n225 ), .B(\us10/n40 ), .Y(\us10/n345 ) );
  INVX1 \us10/U323  ( .A(\us10/n278 ), .Y(\us10/n94 ) );
  NAND2X1 \us10/U322  ( .A(\us10/n94 ), .B(\us10/n226 ), .Y(\us10/n199 ) );
  NAND2X1 \us10/U321  ( .A(\us10/n199 ), .B(\us10/n205 ), .Y(\us10/n82 ) );
  NAND2X1 \us10/U320  ( .A(\us10/n19 ), .B(\us10/n199 ), .Y(\us10/n295 ) );
  NOR2X1 \us10/U319  ( .A(\us10/n226 ), .B(\us10/n259 ), .Y(\us10/n210 ) );
  NOR2X1 \us10/U318  ( .A(\us10/n27 ), .B(\us10/n210 ), .Y(\us10/n173 ) );
  MXI2X1 \us10/U317  ( .A(\us10/n345 ), .B(\us10/n346 ), .S0(\us10/n252 ), .Y(
        \us10/n342 ) );
  NOR2X1 \us10/U316  ( .A(sa10[1]), .B(sa10[3]), .Y(\us10/n163 ) );
  INVX1 \us10/U315  ( .A(\us10/n163 ), .Y(\us10/n37 ) );
  INVX1 \us10/U314  ( .A(\us10/n173 ), .Y(\us10/n344 ) );
  AOI21X1 \us10/U313  ( .A0(\us10/n240 ), .A1(\us10/n37 ), .B0(\us10/n344 ), 
        .Y(\us10/n343 ) );
  AOI211X1 \us10/U312  ( .A0(\us10/n5 ), .A1(\us10/n68 ), .B0(\us10/n342 ), 
        .C0(\us10/n343 ), .Y(\us10/n333 ) );
  NOR2X1 \us10/U311  ( .A(\us10/n18 ), .B(\us10/n226 ), .Y(\us10/n258 ) );
  NAND2X1 \us10/U310  ( .A(\us10/n278 ), .B(sa10[1]), .Y(\us10/n204 ) );
  NOR2X1 \us10/U309  ( .A(\us10/n188 ), .B(sa10[1]), .Y(\us10/n179 ) );
  INVX1 \us10/U308  ( .A(\us10/n179 ), .Y(\us10/n330 ) );
  NAND2X1 \us10/U307  ( .A(\us10/n204 ), .B(\us10/n330 ), .Y(\us10/n239 ) );
  NOR2X1 \us10/U306  ( .A(\us10/n136 ), .B(sa10[1]), .Y(\us10/n299 ) );
  NOR2X1 \us10/U305  ( .A(\us10/n299 ), .B(\us10/n210 ), .Y(\us10/n341 ) );
  OAI32X1 \us10/U304  ( .A0(\us10/n27 ), .A1(\us10/n278 ), .A2(\us10/n95 ), 
        .B0(\us10/n341 ), .B1(\us10/n4 ), .Y(\us10/n340 ) );
  INVX1 \us10/U303  ( .A(\us10/n45 ), .Y(\us10/n126 ) );
  NAND2X1 \us10/U302  ( .A(\us10/n126 ), .B(\us10/n101 ), .Y(\us10/n178 ) );
  NOR2X1 \us10/U301  ( .A(\us10/n18 ), .B(\us10/n136 ), .Y(\us10/n280 ) );
  OAI21XL \us10/U300  ( .A0(\us10/n4 ), .A1(\us10/n121 ), .B0(\us10/n339 ), 
        .Y(\us10/n338 ) );
  MXI2X1 \us10/U299  ( .A(\us10/n336 ), .B(\us10/n337 ), .S0(\us10/n252 ), .Y(
        \us10/n335 ) );
  NOR2X1 \us10/U298  ( .A(\us10/n258 ), .B(\us10/n335 ), .Y(\us10/n334 ) );
  MX4X1 \us10/U297  ( .A(\us10/n331 ), .B(\us10/n332 ), .C(\us10/n333 ), .D(
        \us10/n334 ), .S0(sa10[6]), .S1(\us10/n234 ), .Y(sa13_sr[0]) );
  INVX1 \us10/U296  ( .A(\us10/n299 ), .Y(\us10/n80 ) );
  NOR2X1 \us10/U295  ( .A(\us10/n111 ), .B(\us10/n18 ), .Y(\us10/n269 ) );
  INVX1 \us10/U294  ( .A(\us10/n269 ), .Y(\us10/n75 ) );
  OAI221XL \us10/U293  ( .A0(\us10/n18 ), .A1(\us10/n330 ), .B0(\us10/n20 ), 
        .B1(\us10/n80 ), .C0(\us10/n75 ), .Y(\us10/n329 ) );
  AOI221X1 \us10/U292  ( .A0(\us10/n325 ), .A1(\us10/n33 ), .B0(\us10/n24 ), 
        .B1(\us10/n303 ), .C0(\us10/n329 ), .Y(\us10/n319 ) );
  NOR2X1 \us10/U291  ( .A(\us10/n234 ), .B(sa10[5]), .Y(\us10/n14 ) );
  NOR2X1 \us10/U290  ( .A(\us10/n25 ), .B(\us10/n299 ), .Y(\us10/n313 ) );
  NAND2X1 \us10/U289  ( .A(\us10/n44 ), .B(\us10/n226 ), .Y(\us10/n300 ) );
  AND2X1 \us10/U288  ( .A(\us10/n300 ), .B(\us10/n240 ), .Y(\us10/n23 ) );
  OAI32X1 \us10/U287  ( .A0(\us10/n4 ), .A1(\us10/n145 ), .A2(\us10/n210 ), 
        .B0(\us10/n137 ), .B1(\us10/n27 ), .Y(\us10/n328 ) );
  NOR2X1 \us10/U286  ( .A(sa10[0]), .B(sa10[5]), .Y(\us10/n16 ) );
  INVX1 \us10/U285  ( .A(\us10/n16 ), .Y(\us10/n114 ) );
  INVX1 \us10/U284  ( .A(\us10/n145 ), .Y(\us10/n149 ) );
  NOR2X1 \us10/U283  ( .A(\us10/n47 ), .B(sa10[1]), .Y(\us10/n98 ) );
  INVX1 \us10/U282  ( .A(\us10/n98 ), .Y(\us10/n284 ) );
  OAI21XL \us10/U281  ( .A0(\us10/n69 ), .A1(\us10/n284 ), .B0(\us10/n27 ), 
        .Y(\us10/n327 ) );
  AOI31X1 \us10/U280  ( .A0(\us10/n111 ), .A1(\us10/n149 ), .A2(\us10/n327 ), 
        .B0(\us10/n225 ), .Y(\us10/n326 ) );
  OAI21XL \us10/U279  ( .A0(\us10/n325 ), .A1(\us10/n18 ), .B0(\us10/n326 ), 
        .Y(\us10/n322 ) );
  NAND2X1 \us10/U278  ( .A(\us10/n19 ), .B(\us10/n189 ), .Y(\us10/n71 ) );
  NOR2X1 \us10/U277  ( .A(\us10/n71 ), .B(\us10/n18 ), .Y(\us10/n135 ) );
  AOI21X1 \us10/U276  ( .A0(\us10/n40 ), .A1(sa10[4]), .B0(\us10/n135 ), .Y(
        \us10/n324 ) );
  OAI221XL \us10/U275  ( .A0(\us10/n47 ), .A1(\us10/n27 ), .B0(\us10/n65 ), 
        .B1(\us10/n20 ), .C0(\us10/n324 ), .Y(\us10/n323 ) );
  AOI22X1 \us10/U274  ( .A0(\us10/n55 ), .A1(\us10/n322 ), .B0(\us10/n89 ), 
        .B1(\us10/n323 ), .Y(\us10/n321 ) );
  OAI221XL \us10/U273  ( .A0(\us10/n319 ), .A1(\us10/n52 ), .B0(\us10/n320 ), 
        .B1(\us10/n114 ), .C0(\us10/n321 ), .Y(\us10/n304 ) );
  NOR2X1 \us10/U272  ( .A(\us10/n226 ), .B(\us10/n58 ), .Y(\us10/n290 ) );
  INVX1 \us10/U271  ( .A(\us10/n290 ), .Y(\us10/n200 ) );
  NAND2X1 \us10/U270  ( .A(\us10/n34 ), .B(\us10/n200 ), .Y(\us10/n120 ) );
  INVX1 \us10/U269  ( .A(\us10/n210 ), .Y(\us10/n100 ) );
  OAI221XL \us10/U268  ( .A0(\us10/n20 ), .A1(\us10/n100 ), .B0(sa10[3]), .B1(
        \us10/n4 ), .C0(\us10/n262 ), .Y(\us10/n317 ) );
  INVX1 \us10/U267  ( .A(\us10/n258 ), .Y(\us10/n182 ) );
  AOI211X1 \us10/U266  ( .A0(\us10/n33 ), .A1(\us10/n120 ), .B0(\us10/n317 ), 
        .C0(\us10/n318 ), .Y(\us10/n306 ) );
  NAND2X1 \us10/U265  ( .A(\us10/n100 ), .B(\us10/n199 ), .Y(\us10/n151 ) );
  INVX1 \us10/U264  ( .A(\us10/n151 ), .Y(\us10/n314 ) );
  NOR2X1 \us10/U263  ( .A(\us10/n45 ), .B(\us10/n163 ), .Y(\us10/n160 ) );
  INVX1 \us10/U262  ( .A(\us10/n295 ), .Y(\us10/n92 ) );
  AOI21X1 \us10/U261  ( .A0(sa10[1]), .A1(\us10/n58 ), .B0(\us10/n98 ), .Y(
        \us10/n316 ) );
  OAI22X1 \us10/U260  ( .A0(\us10/n92 ), .A1(\us10/n18 ), .B0(\us10/n316 ), 
        .B1(\us10/n27 ), .Y(\us10/n315 ) );
  NOR2X1 \us10/U259  ( .A(\us10/n149 ), .B(\us10/n226 ), .Y(\us10/n41 ) );
  INVX1 \us10/U258  ( .A(\us10/n41 ), .Y(\us10/n105 ) );
  NAND2X1 \us10/U257  ( .A(\us10/n284 ), .B(\us10/n105 ), .Y(\us10/n227 ) );
  AOI21X1 \us10/U256  ( .A0(\us10/n313 ), .A1(\us10/n33 ), .B0(\us10/n269 ), 
        .Y(\us10/n312 ) );
  OAI221XL \us10/U255  ( .A0(\us10/n149 ), .A1(\us10/n20 ), .B0(\us10/n4 ), 
        .B1(\us10/n227 ), .C0(\us10/n312 ), .Y(\us10/n309 ) );
  AOI21X1 \us10/U254  ( .A0(\us10/n226 ), .A1(\us10/n188 ), .B0(\us10/n242 ), 
        .Y(\us10/n185 ) );
  INVX1 \us10/U253  ( .A(\us10/n185 ), .Y(\us10/n48 ) );
  AND2X1 \us10/U252  ( .A(\us10/n223 ), .B(\us10/n240 ), .Y(\us10/n28 ) );
  OAI221XL \us10/U251  ( .A0(\us10/n27 ), .A1(\us10/n44 ), .B0(\us10/n4 ), 
        .B1(\us10/n48 ), .C0(\us10/n311 ), .Y(\us10/n310 ) );
  AOI22X1 \us10/U250  ( .A0(\us10/n89 ), .A1(\us10/n309 ), .B0(\us10/n55 ), 
        .B1(\us10/n310 ), .Y(\us10/n308 ) );
  OAI221XL \us10/U249  ( .A0(\us10/n306 ), .A1(\us10/n52 ), .B0(\us10/n307 ), 
        .B1(\us10/n114 ), .C0(\us10/n308 ), .Y(\us10/n305 ) );
  MX2X1 \us10/U248  ( .A(\us10/n304 ), .B(\us10/n305 ), .S0(sa10[6]), .Y(
        sa13_sr[1]) );
  INVX1 \us10/U247  ( .A(\us10/n187 ), .Y(\us10/n61 ) );
  MXI2X1 \us10/U246  ( .A(\us10/n303 ), .B(\us10/n61 ), .S0(\us10/n69 ), .Y(
        \us10/n301 ) );
  MXI2X1 \us10/U245  ( .A(\us10/n301 ), .B(\us10/n147 ), .S0(\us10/n302 ), .Y(
        \us10/n285 ) );
  NAND2X1 \us10/U244  ( .A(\us10/n200 ), .B(\us10/n300 ), .Y(\us10/n99 ) );
  INVX1 \us10/U243  ( .A(\us10/n99 ), .Y(\us10/n296 ) );
  NOR2X1 \us10/U242  ( .A(\us10/n299 ), .B(\us10/n242 ), .Y(\us10/n298 ) );
  NAND2X1 \us10/U241  ( .A(sa10[1]), .B(\us10/n47 ), .Y(\us10/n122 ) );
  NOR2X1 \us10/U240  ( .A(\us10/n159 ), .B(\us10/n217 ), .Y(\us10/n198 ) );
  OAI221XL \us10/U239  ( .A0(\us10/n298 ), .A1(\us10/n27 ), .B0(\us10/n20 ), 
        .B1(\us10/n122 ), .C0(\us10/n132 ), .Y(\us10/n297 ) );
  AOI221X1 \us10/U238  ( .A0(\us10/n225 ), .A1(\us10/n226 ), .B0(\us10/n296 ), 
        .B1(\us10/n6 ), .C0(\us10/n297 ), .Y(\us10/n291 ) );
  OAI2BB2X1 \us10/U237  ( .B0(\us10/n27 ), .B1(\us10/n295 ), .A0N(\us10/n34 ), 
        .A1N(\us10/n24 ), .Y(\us10/n293 ) );
  AOI21X1 \us10/U236  ( .A0(\us10/n101 ), .A1(\us10/n150 ), .B0(\us10/n20 ), 
        .Y(\us10/n294 ) );
  AOI211X1 \us10/U235  ( .A0(\us10/n5 ), .A1(\us10/n79 ), .B0(\us10/n293 ), 
        .C0(\us10/n294 ), .Y(\us10/n292 ) );
  INVX1 \us10/U234  ( .A(\us10/n89 ), .Y(\us10/n10 ) );
  OAI22X1 \us10/U233  ( .A0(\us10/n291 ), .A1(\us10/n114 ), .B0(\us10/n292 ), 
        .B1(\us10/n10 ), .Y(\us10/n286 ) );
  INVX1 \us10/U232  ( .A(\us10/n225 ), .Y(\us10/n288 ) );
  NAND2X1 \us10/U231  ( .A(\us10/n200 ), .B(\us10/n284 ), .Y(\us10/n102 ) );
  NOR2X1 \us10/U230  ( .A(\us10/n290 ), .B(\us10/n163 ), .Y(\us10/n184 ) );
  AOI22X1 \us10/U229  ( .A0(\us10/n102 ), .A1(\us10/n69 ), .B0(\us10/n184 ), 
        .B1(\us10/n33 ), .Y(\us10/n289 ) );
  AOI31X1 \us10/U228  ( .A0(\us10/n132 ), .A1(\us10/n288 ), .A2(\us10/n289 ), 
        .B0(\us10/n52 ), .Y(\us10/n287 ) );
  AOI211X1 \us10/U227  ( .A0(\us10/n285 ), .A1(\us10/n55 ), .B0(\us10/n286 ), 
        .C0(\us10/n287 ), .Y(\us10/n263 ) );
  NAND2X1 \us10/U226  ( .A(\us10/n284 ), .B(\us10/n122 ), .Y(\us10/n125 ) );
  NOR2X1 \us10/U225  ( .A(\us10/n199 ), .B(\us10/n4 ), .Y(\us10/n50 ) );
  AOI21X1 \us10/U224  ( .A0(\us10/n200 ), .A1(\us10/n223 ), .B0(\us10/n20 ), 
        .Y(\us10/n283 ) );
  AOI211X1 \us10/U223  ( .A0(\us10/n5 ), .A1(\us10/n125 ), .B0(\us10/n50 ), 
        .C0(\us10/n283 ), .Y(\us10/n282 ) );
  OAI221XL \us10/U222  ( .A0(\us10/n281 ), .A1(\us10/n27 ), .B0(\us10/n4 ), 
        .B1(\us10/n111 ), .C0(\us10/n282 ), .Y(\us10/n265 ) );
  INVX1 \us10/U221  ( .A(\us10/n280 ), .Y(\us10/n247 ) );
  NAND2X1 \us10/U220  ( .A(\us10/n41 ), .B(\us10/n33 ), .Y(\us10/n272 ) );
  OAI221XL \us10/U219  ( .A0(sa10[1]), .A1(\us10/n247 ), .B0(\us10/n4 ), .B1(
        \us10/n189 ), .C0(\us10/n272 ), .Y(\us10/n279 ) );
  NAND2X1 \us10/U218  ( .A(sa10[2]), .B(\us10/n149 ), .Y(\us10/n276 ) );
  XNOR2X1 \us10/U217  ( .A(\us10/n129 ), .B(sa10[1]), .Y(\us10/n155 ) );
  MXI2X1 \us10/U216  ( .A(\us10/n276 ), .B(\us10/n277 ), .S0(\us10/n155 ), .Y(
        \us10/n275 ) );
  OAI22X1 \us10/U215  ( .A0(\us10/n273 ), .A1(\us10/n10 ), .B0(\us10/n274 ), 
        .B1(\us10/n52 ), .Y(\us10/n266 ) );
  NOR2X1 \us10/U214  ( .A(\us10/n20 ), .B(\us10/n226 ), .Y(\us10/n176 ) );
  OAI21XL \us10/U213  ( .A0(\us10/n4 ), .A1(\us10/n271 ), .B0(\us10/n272 ), 
        .Y(\us10/n270 ) );
  OAI31X1 \us10/U212  ( .A0(\us10/n176 ), .A1(\us10/n269 ), .A2(\us10/n270 ), 
        .B0(\us10/n16 ), .Y(\us10/n268 ) );
  INVX1 \us10/U211  ( .A(\us10/n268 ), .Y(\us10/n267 ) );
  AOI211X1 \us10/U210  ( .A0(\us10/n55 ), .A1(\us10/n265 ), .B0(\us10/n266 ), 
        .C0(\us10/n267 ), .Y(\us10/n264 ) );
  MXI2X1 \us10/U209  ( .A(\us10/n263 ), .B(\us10/n264 ), .S0(sa10[6]), .Y(
        sa13_sr[2]) );
  NOR2X1 \us10/U208  ( .A(\us10/n94 ), .B(sa10[1]), .Y(\us10/n211 ) );
  INVX1 \us10/U207  ( .A(\us10/n262 ), .Y(\us10/n261 ) );
  AOI211X1 \us10/U206  ( .A0(\us10/n259 ), .A1(\us10/n24 ), .B0(\us10/n260 ), 
        .C0(\us10/n261 ), .Y(\us10/n255 ) );
  OAI22X1 \us10/U205  ( .A0(\us10/n20 ), .A1(\us10/n68 ), .B0(\us10/n27 ), 
        .B1(\us10/n37 ), .Y(\us10/n257 ) );
  NOR3X1 \us10/U204  ( .A(\us10/n257 ), .B(\us10/n258 ), .C(\us10/n50 ), .Y(
        \us10/n256 ) );
  MXI2X1 \us10/U203  ( .A(\us10/n255 ), .B(\us10/n256 ), .S0(\us10/n252 ), .Y(
        \us10/n254 ) );
  AOI221X1 \us10/U202  ( .A0(\us10/n211 ), .A1(\us10/n5 ), .B0(\us10/n40 ), 
        .B1(sa10[4]), .C0(\us10/n254 ), .Y(\us10/n248 ) );
  INVX1 \us10/U201  ( .A(\us10/n211 ), .Y(\us10/n106 ) );
  NAND2X1 \us10/U200  ( .A(\us10/n200 ), .B(\us10/n106 ), .Y(\us10/n83 ) );
  NAND2X1 \us10/U199  ( .A(\us10/n199 ), .B(\us10/n204 ), .Y(\us10/n169 ) );
  AOI2BB2X1 \us10/U198  ( .B0(\us10/n65 ), .B1(\us10/n24 ), .A0N(\us10/n169 ), 
        .A1N(\us10/n20 ), .Y(\us10/n253 ) );
  OAI221XL \us10/U197  ( .A0(\us10/n172 ), .A1(\us10/n18 ), .B0(\us10/n27 ), 
        .B1(\us10/n83 ), .C0(\us10/n253 ), .Y(\us10/n251 ) );
  MXI2X1 \us10/U196  ( .A(\us10/n250 ), .B(\us10/n251 ), .S0(\us10/n252 ), .Y(
        \us10/n249 ) );
  MXI2X1 \us10/U195  ( .A(\us10/n248 ), .B(\us10/n249 ), .S0(\us10/n234 ), .Y(
        \us10/n228 ) );
  OAI21XL \us10/U194  ( .A0(\us10/n58 ), .A1(\us10/n27 ), .B0(\us10/n247 ), 
        .Y(\us10/n245 ) );
  NOR2X1 \us10/U193  ( .A(sa10[7]), .B(\us10/n145 ), .Y(\us10/n246 ) );
  XNOR2X1 \us10/U192  ( .A(\us10/n69 ), .B(sa10[1]), .Y(\us10/n130 ) );
  MXI2X1 \us10/U191  ( .A(\us10/n245 ), .B(\us10/n246 ), .S0(\us10/n130 ), .Y(
        \us10/n243 ) );
  OAI211X1 \us10/U190  ( .A0(\us10/n4 ), .A1(\us10/n149 ), .B0(\us10/n243 ), 
        .C0(\us10/n244 ), .Y(\us10/n230 ) );
  NOR2X1 \us10/U189  ( .A(\us10/n242 ), .B(\us10/n137 ), .Y(\us10/n70 ) );
  OAI221XL \us10/U188  ( .A0(\us10/n159 ), .A1(\us10/n27 ), .B0(\us10/n20 ), 
        .B1(\us10/n34 ), .C0(\us10/n241 ), .Y(\us10/n231 ) );
  NAND2X1 \us10/U187  ( .A(\us10/n101 ), .B(\us10/n240 ), .Y(\us10/n76 ) );
  AOI21X1 \us10/U186  ( .A0(\us10/n122 ), .A1(\us10/n106 ), .B0(\us10/n129 ), 
        .Y(\us10/n237 ) );
  INVX1 \us10/U185  ( .A(\us10/n239 ), .Y(\us10/n238 ) );
  OAI21XL \us10/U184  ( .A0(\us10/n237 ), .A1(\us10/n43 ), .B0(\us10/n238 ), 
        .Y(\us10/n236 ) );
  OAI221XL \us10/U183  ( .A0(\us10/n18 ), .A1(\us10/n76 ), .B0(\us10/n59 ), 
        .B1(\us10/n27 ), .C0(\us10/n236 ), .Y(\us10/n232 ) );
  AOI2BB2X1 \us10/U182  ( .B0(\us10/n24 ), .B1(\us10/n187 ), .A0N(\us10/n227 ), 
        .A1N(\us10/n20 ), .Y(\us10/n235 ) );
  OAI211X1 \us10/U181  ( .A0(\us10/n27 ), .A1(\us10/n122 ), .B0(\us10/n158 ), 
        .C0(\us10/n235 ), .Y(\us10/n233 ) );
  MX4X1 \us10/U180  ( .A(\us10/n230 ), .B(\us10/n231 ), .C(\us10/n232 ), .D(
        \us10/n233 ), .S0(\us10/n234 ), .S1(sa10[5]), .Y(\us10/n229 ) );
  MX2X1 \us10/U179  ( .A(\us10/n228 ), .B(\us10/n229 ), .S0(sa10[6]), .Y(
        sa13_sr[3]) );
  NOR2BX1 \us10/U178  ( .AN(\us10/n204 ), .B(\us10/n137 ), .Y(\us10/n110 ) );
  INVX1 \us10/U177  ( .A(\us10/n110 ), .Y(\us10/n64 ) );
  AOI22X1 \us10/U176  ( .A0(\us10/n225 ), .A1(\us10/n226 ), .B0(\us10/n6 ), 
        .B1(\us10/n227 ), .Y(\us10/n224 ) );
  OAI221XL \us10/U175  ( .A0(\us10/n27 ), .A1(\us10/n64 ), .B0(\us10/n4 ), 
        .B1(\us10/n83 ), .C0(\us10/n224 ), .Y(\us10/n212 ) );
  NAND2X1 \us10/U174  ( .A(\us10/n34 ), .B(\us10/n204 ), .Y(\us10/n221 ) );
  OAI21XL \us10/U173  ( .A0(\us10/n69 ), .A1(\us10/n223 ), .B0(\us10/n27 ), 
        .Y(\us10/n222 ) );
  NOR2X1 \us10/U172  ( .A(\us10/n217 ), .B(\us10/n42 ), .Y(\us10/n208 ) );
  AOI211X1 \us10/U171  ( .A0(\us10/n208 ), .A1(\us10/n5 ), .B0(\us10/n220 ), 
        .C0(\us10/n173 ), .Y(\us10/n219 ) );
  OAI22X1 \us10/U170  ( .A0(\us10/n218 ), .A1(\us10/n10 ), .B0(\us10/n219 ), 
        .B1(\us10/n114 ), .Y(\us10/n213 ) );
  INVX1 \us10/U169  ( .A(\us10/n135 ), .Y(\us10/n215 ) );
  NOR2X1 \us10/U168  ( .A(\us10/n4 ), .B(\us10/n159 ), .Y(\us10/n31 ) );
  INVX1 \us10/U167  ( .A(\us10/n31 ), .Y(\us10/n196 ) );
  AOI31X1 \us10/U166  ( .A0(\us10/n215 ), .A1(\us10/n196 ), .A2(\us10/n216 ), 
        .B0(\us10/n52 ), .Y(\us10/n214 ) );
  AOI211X1 \us10/U165  ( .A0(\us10/n55 ), .A1(\us10/n212 ), .B0(\us10/n213 ), 
        .C0(\us10/n214 ), .Y(\us10/n190 ) );
  INVX1 \us10/U164  ( .A(\us10/n207 ), .Y(\us10/n192 ) );
  NOR2X1 \us10/U163  ( .A(\us10/n25 ), .B(\us10/n98 ), .Y(\us10/n32 ) );
  OAI22X1 \us10/U162  ( .A0(\us10/n28 ), .A1(\us10/n4 ), .B0(\us10/n188 ), 
        .B1(\us10/n27 ), .Y(\us10/n206 ) );
  NAND2X1 \us10/U161  ( .A(\us10/n204 ), .B(\us10/n80 ), .Y(\us10/n118 ) );
  INVX1 \us10/U160  ( .A(\us10/n118 ), .Y(\us10/n123 ) );
  NAND2X1 \us10/U159  ( .A(\us10/n94 ), .B(\us10/n79 ), .Y(\us10/n203 ) );
  OAI2BB1X1 \us10/U158  ( .A0N(\us10/n199 ), .A1N(\us10/n200 ), .B0(\us10/n33 ), .Y(\us10/n195 ) );
  INVX1 \us10/U157  ( .A(\us10/n55 ), .Y(\us10/n12 ) );
  AOI31X1 \us10/U156  ( .A0(\us10/n195 ), .A1(\us10/n196 ), .A2(\us10/n197 ), 
        .B0(\us10/n12 ), .Y(\us10/n194 ) );
  AOI211X1 \us10/U155  ( .A0(\us10/n89 ), .A1(\us10/n192 ), .B0(\us10/n193 ), 
        .C0(\us10/n194 ), .Y(\us10/n191 ) );
  MXI2X1 \us10/U154  ( .A(\us10/n190 ), .B(\us10/n191 ), .S0(sa10[6]), .Y(
        sa13_sr[4]) );
  OAI21XL \us10/U153  ( .A0(\us10/n69 ), .A1(\us10/n189 ), .B0(\us10/n27 ), 
        .Y(\us10/n186 ) );
  INVX1 \us10/U152  ( .A(\us10/n183 ), .Y(\us10/n180 ) );
  NAND2X1 \us10/U151  ( .A(\us10/n74 ), .B(\us10/n182 ), .Y(\us10/n181 ) );
  AOI211X1 \us10/U150  ( .A0(\us10/n179 ), .A1(\us10/n24 ), .B0(\us10/n180 ), 
        .C0(\us10/n181 ), .Y(\us10/n165 ) );
  INVX1 \us10/U149  ( .A(\us10/n178 ), .Y(\us10/n175 ) );
  AOI211X1 \us10/U148  ( .A0(\us10/n175 ), .A1(\us10/n5 ), .B0(\us10/n176 ), 
        .C0(\us10/n177 ), .Y(\us10/n174 ) );
  OAI221XL \us10/U147  ( .A0(\us10/n159 ), .A1(\us10/n27 ), .B0(\us10/n145 ), 
        .B1(\us10/n20 ), .C0(\us10/n174 ), .Y(\us10/n167 ) );
  MXI2X1 \us10/U146  ( .A(\us10/n40 ), .B(\us10/n173 ), .S0(\us10/n96 ), .Y(
        \us10/n170 ) );
  AOI22X1 \us10/U145  ( .A0(\us10/n137 ), .A1(\us10/n24 ), .B0(\us10/n172 ), 
        .B1(\us10/n6 ), .Y(\us10/n171 ) );
  OAI211X1 \us10/U144  ( .A0(\us10/n20 ), .A1(\us10/n169 ), .B0(\us10/n170 ), 
        .C0(\us10/n171 ), .Y(\us10/n168 ) );
  AOI22X1 \us10/U143  ( .A0(\us10/n89 ), .A1(\us10/n167 ), .B0(\us10/n55 ), 
        .B1(\us10/n168 ), .Y(\us10/n166 ) );
  OAI221XL \us10/U142  ( .A0(\us10/n164 ), .A1(\us10/n114 ), .B0(\us10/n165 ), 
        .B1(\us10/n52 ), .C0(\us10/n166 ), .Y(\us10/n138 ) );
  OAI21XL \us10/U141  ( .A0(\us10/n41 ), .A1(\us10/n163 ), .B0(\us10/n69 ), 
        .Y(\us10/n162 ) );
  AOI221X1 \us10/U140  ( .A0(\us10/n159 ), .A1(\us10/n24 ), .B0(\us10/n160 ), 
        .B1(\us10/n33 ), .C0(\us10/n161 ), .Y(\us10/n140 ) );
  OAI21XL \us10/U139  ( .A0(\us10/n157 ), .A1(\us10/n20 ), .B0(\us10/n158 ), 
        .Y(\us10/n156 ) );
  NOR2X1 \us10/U138  ( .A(\us10/n4 ), .B(\us10/n136 ), .Y(\us10/n153 ) );
  NOR2X1 \us10/U137  ( .A(\us10/n145 ), .B(\us10/n69 ), .Y(\us10/n154 ) );
  MXI2X1 \us10/U136  ( .A(\us10/n153 ), .B(\us10/n154 ), .S0(\us10/n155 ), .Y(
        \us10/n152 ) );
  OAI221XL \us10/U135  ( .A0(\us10/n110 ), .A1(\us10/n18 ), .B0(\us10/n20 ), 
        .B1(\us10/n151 ), .C0(\us10/n152 ), .Y(\us10/n143 ) );
  AOI21X1 \us10/U134  ( .A0(\us10/n149 ), .A1(\us10/n150 ), .B0(\us10/n18 ), 
        .Y(\us10/n148 ) );
  AOI2BB1X1 \us10/U133  ( .A0N(\us10/n147 ), .A1N(\us10/n27 ), .B0(\us10/n148 ), .Y(\us10/n146 ) );
  OAI221XL \us10/U132  ( .A0(\us10/n145 ), .A1(\us10/n20 ), .B0(\us10/n4 ), 
        .B1(\us10/n34 ), .C0(\us10/n146 ), .Y(\us10/n144 ) );
  AOI22X1 \us10/U131  ( .A0(\us10/n89 ), .A1(\us10/n143 ), .B0(\us10/n14 ), 
        .B1(\us10/n144 ), .Y(\us10/n142 ) );
  OAI221XL \us10/U130  ( .A0(\us10/n140 ), .A1(\us10/n12 ), .B0(\us10/n141 ), 
        .B1(\us10/n114 ), .C0(\us10/n142 ), .Y(\us10/n139 ) );
  MX2X1 \us10/U129  ( .A(\us10/n138 ), .B(\us10/n139 ), .S0(sa10[6]), .Y(
        sa13_sr[5]) );
  INVX1 \us10/U128  ( .A(\us10/n70 ), .Y(\us10/n133 ) );
  OAI22X1 \us10/U127  ( .A0(\us10/n4 ), .A1(\us10/n136 ), .B0(\us10/n137 ), 
        .B1(\us10/n27 ), .Y(\us10/n134 ) );
  AOI211X1 \us10/U126  ( .A0(\us10/n133 ), .A1(\us10/n69 ), .B0(\us10/n134 ), 
        .C0(\us10/n135 ), .Y(\us10/n112 ) );
  INVX1 \us10/U125  ( .A(\us10/n132 ), .Y(\us10/n131 ) );
  OAI21XL \us10/U124  ( .A0(\us10/n18 ), .A1(\us10/n37 ), .B0(\us10/n128 ), 
        .Y(\us10/n127 ) );
  OAI221XL \us10/U123  ( .A0(\us10/n18 ), .A1(\us10/n105 ), .B0(\us10/n123 ), 
        .B1(\us10/n27 ), .C0(\us10/n124 ), .Y(\us10/n116 ) );
  NAND2X1 \us10/U122  ( .A(\us10/n121 ), .B(\us10/n122 ), .Y(\us10/n30 ) );
  OAI221XL \us10/U121  ( .A0(\us10/n18 ), .A1(\us10/n118 ), .B0(\us10/n27 ), 
        .B1(\us10/n30 ), .C0(\us10/n119 ), .Y(\us10/n117 ) );
  AOI22X1 \us10/U120  ( .A0(\us10/n89 ), .A1(\us10/n116 ), .B0(\us10/n55 ), 
        .B1(\us10/n117 ), .Y(\us10/n115 ) );
  OAI221XL \us10/U119  ( .A0(\us10/n112 ), .A1(\us10/n52 ), .B0(\us10/n113 ), 
        .B1(\us10/n114 ), .C0(\us10/n115 ), .Y(\us10/n84 ) );
  OAI22X1 \us10/U118  ( .A0(\us10/n110 ), .A1(\us10/n4 ), .B0(\us10/n20 ), 
        .B1(\us10/n21 ), .Y(\us10/n108 ) );
  AOI21X1 \us10/U117  ( .A0(sa10[1]), .A1(\us10/n58 ), .B0(\us10/n27 ), .Y(
        \us10/n109 ) );
  AOI211X1 \us10/U116  ( .A0(\us10/n5 ), .A1(\us10/n107 ), .B0(\us10/n108 ), 
        .C0(\us10/n109 ), .Y(\us10/n86 ) );
  OAI22X1 \us10/U115  ( .A0(\us10/n45 ), .A1(\us10/n4 ), .B0(sa10[4]), .B1(
        \us10/n18 ), .Y(\us10/n103 ) );
  AOI21X1 \us10/U114  ( .A0(\us10/n105 ), .A1(\us10/n106 ), .B0(\us10/n20 ), 
        .Y(\us10/n104 ) );
  AOI211X1 \us10/U113  ( .A0(\us10/n33 ), .A1(\us10/n102 ), .B0(\us10/n103 ), 
        .C0(\us10/n104 ), .Y(\us10/n87 ) );
  NAND2X1 \us10/U112  ( .A(\us10/n100 ), .B(\us10/n101 ), .Y(\us10/n62 ) );
  OAI221XL \us10/U111  ( .A0(\us10/n27 ), .A1(\us10/n62 ), .B0(\us10/n4 ), 
        .B1(\us10/n21 ), .C0(\us10/n97 ), .Y(\us10/n90 ) );
  NOR3X1 \us10/U110  ( .A(\us10/n4 ), .B(\us10/n95 ), .C(\us10/n96 ), .Y(
        \us10/n67 ) );
  AOI31X1 \us10/U109  ( .A0(\us10/n79 ), .A1(\us10/n94 ), .A2(\us10/n6 ), .B0(
        \us10/n67 ), .Y(\us10/n93 ) );
  OAI221XL \us10/U108  ( .A0(\us10/n73 ), .A1(\us10/n27 ), .B0(\us10/n92 ), 
        .B1(\us10/n20 ), .C0(\us10/n93 ), .Y(\us10/n91 ) );
  AOI22X1 \us10/U107  ( .A0(\us10/n89 ), .A1(\us10/n90 ), .B0(\us10/n16 ), 
        .B1(\us10/n91 ), .Y(\us10/n88 ) );
  OAI221XL \us10/U106  ( .A0(\us10/n86 ), .A1(\us10/n52 ), .B0(\us10/n87 ), 
        .B1(\us10/n12 ), .C0(\us10/n88 ), .Y(\us10/n85 ) );
  MX2X1 \us10/U105  ( .A(\us10/n84 ), .B(\us10/n85 ), .S0(sa10[6]), .Y(
        sa13_sr[6]) );
  INVX1 \us10/U104  ( .A(\us10/n81 ), .Y(\us10/n77 ) );
  AOI21X1 \us10/U103  ( .A0(\us10/n79 ), .A1(\us10/n80 ), .B0(\us10/n27 ), .Y(
        \us10/n78 ) );
  AOI211X1 \us10/U102  ( .A0(\us10/n5 ), .A1(\us10/n76 ), .B0(\us10/n77 ), 
        .C0(\us10/n78 ), .Y(\us10/n51 ) );
  OAI211X1 \us10/U101  ( .A0(\us10/n73 ), .A1(\us10/n27 ), .B0(\us10/n74 ), 
        .C0(\us10/n75 ), .Y(\us10/n72 ) );
  AOI21X1 \us10/U100  ( .A0(\us10/n68 ), .A1(\us10/n69 ), .B0(\us10/n6 ), .Y(
        \us10/n63 ) );
  INVX1 \us10/U99  ( .A(\us10/n67 ), .Y(\us10/n66 ) );
  OAI221XL \us10/U98  ( .A0(\us10/n63 ), .A1(\us10/n64 ), .B0(\us10/n65 ), 
        .B1(\us10/n27 ), .C0(\us10/n66 ), .Y(\us10/n56 ) );
  AOI2BB2X1 \us10/U97  ( .B0(\us10/n61 ), .B1(\us10/n24 ), .A0N(\us10/n62 ), 
        .A1N(\us10/n20 ), .Y(\us10/n60 ) );
  OAI221XL \us10/U96  ( .A0(\us10/n58 ), .A1(\us10/n18 ), .B0(\us10/n59 ), 
        .B1(\us10/n27 ), .C0(\us10/n60 ), .Y(\us10/n57 ) );
  AOI22X1 \us10/U95  ( .A0(\us10/n55 ), .A1(\us10/n56 ), .B0(\us10/n16 ), .B1(
        \us10/n57 ), .Y(\us10/n54 ) );
  OAI221XL \us10/U94  ( .A0(\us10/n51 ), .A1(\us10/n52 ), .B0(\us10/n53 ), 
        .B1(\us10/n10 ), .C0(\us10/n54 ), .Y(\us10/n7 ) );
  INVX1 \us10/U93  ( .A(\us10/n50 ), .Y(\us10/n49 ) );
  OAI221XL \us10/U92  ( .A0(\us10/n47 ), .A1(\us10/n18 ), .B0(\us10/n27 ), 
        .B1(\us10/n48 ), .C0(\us10/n49 ), .Y(\us10/n46 ) );
  NOR2X1 \us10/U91  ( .A(\us10/n41 ), .B(\us10/n42 ), .Y(\us10/n38 ) );
  INVX1 \us10/U90  ( .A(\us10/n40 ), .Y(\us10/n39 ) );
  INVX1 \us10/U89  ( .A(\us10/n32 ), .Y(\us10/n26 ) );
  AOI21X1 \us10/U88  ( .A0(\us10/n5 ), .A1(\us10/n30 ), .B0(\us10/n31 ), .Y(
        \us10/n29 ) );
  OAI221XL \us10/U87  ( .A0(\us10/n26 ), .A1(\us10/n27 ), .B0(\us10/n28 ), 
        .B1(\us10/n20 ), .C0(\us10/n29 ), .Y(\us10/n15 ) );
  OAI221XL \us10/U86  ( .A0(\us10/n18 ), .A1(\us10/n19 ), .B0(\us10/n20 ), 
        .B1(\us10/n21 ), .C0(\us10/n22 ), .Y(\us10/n17 ) );
  AOI22X1 \us10/U85  ( .A0(\us10/n14 ), .A1(\us10/n15 ), .B0(\us10/n16 ), .B1(
        \us10/n17 ), .Y(\us10/n13 ) );
  OAI221XL \us10/U84  ( .A0(\us10/n9 ), .A1(\us10/n10 ), .B0(\us10/n11 ), .B1(
        \us10/n12 ), .C0(\us10/n13 ), .Y(\us10/n8 ) );
  MX2X1 \us10/U83  ( .A(\us10/n7 ), .B(\us10/n8 ), .S0(sa10[6]), .Y(sa13_sr[7]) );
  NOR2X4 \us10/U82  ( .A(\us10/n129 ), .B(sa10[2]), .Y(\us10/n43 ) );
  CLKINVX3 \us10/U81  ( .A(\us10/n14 ), .Y(\us10/n52 ) );
  OAI22XL \us10/U80  ( .A0(\us10/n201 ), .A1(\us10/n52 ), .B0(\us10/n202 ), 
        .B1(\us10/n114 ), .Y(\us10/n193 ) );
  CLKINVX3 \us10/U79  ( .A(sa10[5]), .Y(\us10/n252 ) );
  NOR2X2 \us10/U78  ( .A(\us10/n252 ), .B(\us10/n234 ), .Y(\us10/n55 ) );
  CLKINVX3 \us10/U77  ( .A(sa10[7]), .Y(\us10/n129 ) );
  NOR2X4 \us10/U76  ( .A(\us10/n129 ), .B(\us10/n69 ), .Y(\us10/n24 ) );
  AOI22XL \us10/U75  ( .A0(\us10/n70 ), .A1(\us10/n24 ), .B0(\us10/n96 ), .B1(
        \us10/n129 ), .Y(\us10/n241 ) );
  NOR2X2 \us10/U74  ( .A(\us10/n252 ), .B(sa10[0]), .Y(\us10/n89 ) );
  CLKINVX3 \us10/U73  ( .A(sa10[0]), .Y(\us10/n234 ) );
  NOR2X4 \us10/U72  ( .A(\us10/n69 ), .B(sa10[7]), .Y(\us10/n33 ) );
  INVX12 \us10/U71  ( .A(\us10/n33 ), .Y(\us10/n27 ) );
  CLKINVX3 \us10/U70  ( .A(\us10/n1 ), .Y(\us10/n6 ) );
  CLKINVX3 \us10/U69  ( .A(\us10/n1 ), .Y(\us10/n5 ) );
  INVXL \us10/U68  ( .A(\us10/n24 ), .Y(\us10/n36 ) );
  INVX4 \us10/U67  ( .A(\us10/n3 ), .Y(\us10/n4 ) );
  INVXL \us10/U66  ( .A(\us10/n36 ), .Y(\us10/n3 ) );
  INVX4 \us10/U65  ( .A(sa10[1]), .Y(\us10/n226 ) );
  INVX4 \us10/U64  ( .A(\us10/n43 ), .Y(\us10/n20 ) );
  AOI221X4 \us10/U63  ( .A0(\us10/n24 ), .A1(\us10/n82 ), .B0(\us10/n43 ), 
        .B1(\us10/n295 ), .C0(\us10/n173 ), .Y(\us10/n346 ) );
  AOI221X4 \us10/U62  ( .A0(\us10/n5 ), .A1(\us10/n96 ), .B0(\us10/n43 ), .B1(
        \us10/n239 ), .C0(\us10/n340 ), .Y(\us10/n336 ) );
  AOI222X4 \us10/U61  ( .A0(\us10/n59 ), .A1(\us10/n43 ), .B0(\us10/n6 ), .B1(
        \us10/n221 ), .C0(\us10/n222 ), .C1(\us10/n187 ), .Y(\us10/n218 ) );
  AOI222X4 \us10/U60  ( .A0(\us10/n123 ), .A1(\us10/n43 ), .B0(sa10[2]), .B1(
        \us10/n203 ), .C0(\us10/n6 ), .C1(\us10/n71 ), .Y(\us10/n202 ) );
  AOI221X4 \us10/U59  ( .A0(\us10/n314 ), .A1(\us10/n43 ), .B0(\us10/n160 ), 
        .B1(\us10/n24 ), .C0(\us10/n315 ), .Y(\us10/n307 ) );
  AOI221X4 \us10/U58  ( .A0(\us10/n43 ), .A1(\us10/n208 ), .B0(\us10/n76 ), 
        .B1(\us10/n24 ), .C0(\us10/n209 ), .Y(\us10/n207 ) );
  AOI221X4 \us10/U57  ( .A0(\us10/n43 ), .A1(\us10/n205 ), .B0(\us10/n32 ), 
        .B1(\us10/n6 ), .C0(\us10/n206 ), .Y(\us10/n201 ) );
  AOI221X4 \us10/U56  ( .A0(\us10/n43 ), .A1(\us10/n44 ), .B0(\us10/n45 ), 
        .B1(\us10/n24 ), .C0(\us10/n46 ), .Y(\us10/n9 ) );
  AOI22XL \us10/U55  ( .A0(\us10/n217 ), .A1(\us10/n43 ), .B0(\us10/n33 ), 
        .B1(\us10/n47 ), .Y(\us10/n216 ) );
  AOI22XL \us10/U54  ( .A0(\us10/n98 ), .A1(\us10/n43 ), .B0(\us10/n6 ), .B1(
        \us10/n99 ), .Y(\us10/n97 ) );
  AOI22XL \us10/U53  ( .A0(\us10/n82 ), .A1(\us10/n43 ), .B0(\us10/n83 ), .B1(
        \us10/n24 ), .Y(\us10/n81 ) );
  AOI2BB2XL \us10/U52  ( .B0(\us10/n43 ), .B1(\us10/n94 ), .A0N(\us10/n120 ), 
        .A1N(\us10/n4 ), .Y(\us10/n119 ) );
  AOI222X4 \us10/U51  ( .A0(\us10/n125 ), .A1(\us10/n33 ), .B0(\us10/n145 ), 
        .B1(\us10/n40 ), .C0(\us10/n43 ), .C1(\us10/n184 ), .Y(\us10/n183 ) );
  AOI22XL \us10/U50  ( .A0(\us10/n43 ), .A1(\us10/n303 ), .B0(\us10/n24 ), 
        .B1(\us10/n96 ), .Y(\us10/n358 ) );
  AOI22XL \us10/U49  ( .A0(\us10/n43 ), .A1(\us10/n100 ), .B0(\us10/n24 ), 
        .B1(\us10/n125 ), .Y(\us10/n124 ) );
  AOI21XL \us10/U48  ( .A0(\us10/n159 ), .A1(\us10/n43 ), .B0(\us10/n40 ), .Y(
        \us10/n262 ) );
  AOI22XL \us10/U47  ( .A0(\us10/n40 ), .A1(\us10/n94 ), .B0(\us10/n43 ), .B1(
        \us10/n187 ), .Y(\us10/n244 ) );
  AOI22XL \us10/U46  ( .A0(\us10/n184 ), .A1(\us10/n5 ), .B0(\us10/n198 ), 
        .B1(\us10/n43 ), .Y(\us10/n197 ) );
  NOR2XL \us10/U45  ( .A(\us10/n33 ), .B(\us10/n2 ), .Y(\us10/n302 ) );
  MXI2XL \us10/U44  ( .A(\us10/n2 ), .B(\us10/n6 ), .S0(\us10/n28 ), .Y(
        \us10/n311 ) );
  INVXL \us10/U43  ( .A(\us10/n20 ), .Y(\us10/n2 ) );
  INVX4 \us10/U42  ( .A(\us10/n6 ), .Y(\us10/n18 ) );
  AOI21XL \us10/U41  ( .A0(\us10/n18 ), .A1(\us10/n162 ), .B0(\us10/n25 ), .Y(
        \us10/n161 ) );
  INVX4 \us10/U40  ( .A(sa10[2]), .Y(\us10/n69 ) );
  NOR2X4 \us10/U39  ( .A(\us10/n226 ), .B(\us10/n4 ), .Y(\us10/n40 ) );
  CLKINVX3 \us10/U38  ( .A(sa10[3]), .Y(\us10/n136 ) );
  NOR2X2 \us10/U37  ( .A(\us10/n136 ), .B(sa10[4]), .Y(\us10/n145 ) );
  CLKINVX3 \us10/U36  ( .A(sa10[4]), .Y(\us10/n58 ) );
  NOR2X2 \us10/U35  ( .A(\us10/n58 ), .B(sa10[3]), .Y(\us10/n159 ) );
  NOR2X2 \us10/U34  ( .A(\us10/n136 ), .B(\us10/n58 ), .Y(\us10/n259 ) );
  NOR2X2 \us10/U33  ( .A(sa10[4]), .B(sa10[3]), .Y(\us10/n278 ) );
  NOR2X2 \us10/U32  ( .A(\us10/n259 ), .B(\us10/n278 ), .Y(\us10/n47 ) );
  CLKINVX3 \us10/U31  ( .A(\us10/n259 ), .Y(\us10/n44 ) );
  NOR2X2 \us10/U30  ( .A(\us10/n44 ), .B(sa10[1]), .Y(\us10/n137 ) );
  AOI21XL \us10/U29  ( .A0(\us10/n44 ), .A1(\us10/n111 ), .B0(\us10/n4 ), .Y(
        \us10/n177 ) );
  AOI22XL \us10/U28  ( .A0(\us10/n23 ), .A1(\us10/n24 ), .B0(\us10/n25 ), .B1(
        sa10[2]), .Y(\us10/n22 ) );
  AOI22XL \us10/U27  ( .A0(\us10/n33 ), .A1(sa10[3]), .B0(\us10/n24 ), .B1(
        \us10/n58 ), .Y(\us10/n277 ) );
  NAND2XL \us10/U26  ( .A(\us10/n198 ), .B(\us10/n24 ), .Y(\us10/n132 ) );
  OAI2BB2XL \us10/U25  ( .B0(\us10/n20 ), .B1(\us10/n111 ), .A0N(\us10/n125 ), 
        .A1N(\us10/n24 ), .Y(\us10/n220 ) );
  NAND2XL \us10/U24  ( .A(\us10/n111 ), .B(\us10/n101 ), .Y(\us10/n21 ) );
  NAND2XL \us10/U23  ( .A(\us10/n111 ), .B(\us10/n300 ), .Y(\us10/n187 ) );
  NAND2XL \us10/U22  ( .A(\us10/n111 ), .B(\us10/n121 ), .Y(\us10/n303 ) );
  AOI221XL \us10/U21  ( .A0(\us10/n43 ), .A1(\us10/n151 ), .B0(\us10/n25 ), 
        .B1(\us10/n69 ), .C0(\us10/n275 ), .Y(\us10/n274 ) );
  NOR2BXL \us10/U20  ( .AN(\us10/n101 ), .B(\us10/n25 ), .Y(\us10/n172 ) );
  NAND2X2 \us10/U19  ( .A(\us10/n58 ), .B(\us10/n226 ), .Y(\us10/n34 ) );
  OAI222X1 \us10/U18  ( .A0(\us10/n27 ), .A1(\us10/n34 ), .B0(\us10/n69 ), 
        .B1(\us10/n205 ), .C0(\us10/n20 ), .C1(\us10/n79 ), .Y(\us10/n260 ) );
  OAI222X1 \us10/U17  ( .A0(\us10/n20 ), .A1(\us10/n99 ), .B0(\us10/n27 ), 
        .B1(\us10/n101 ), .C0(\us10/n184 ), .C1(\us10/n4 ), .Y(\us10/n250 ) );
  OAI222X1 \us10/U16  ( .A0(\us10/n4 ), .A1(\us10/n37 ), .B0(\us10/n38 ), .B1(
        \us10/n20 ), .C0(sa10[4]), .C1(\us10/n39 ), .Y(\us10/n35 ) );
  AOI221X1 \us10/U15  ( .A0(\us10/n5 ), .A1(\us10/n19 ), .B0(\us10/n33 ), .B1(
        \us10/n34 ), .C0(\us10/n35 ), .Y(\us10/n11 ) );
  OR2X2 \us10/U14  ( .A(sa10[2]), .B(sa10[7]), .Y(\us10/n1 ) );
  AOI221XL \us10/U13  ( .A0(\us10/n70 ), .A1(\us10/n43 ), .B0(\us10/n24 ), 
        .B1(\us10/n71 ), .C0(\us10/n72 ), .Y(\us10/n53 ) );
  AOI221XL \us10/U12  ( .A0(\us10/n59 ), .A1(\us10/n33 ), .B0(\us10/n43 ), 
        .B1(\us10/n126 ), .C0(\us10/n127 ), .Y(\us10/n113 ) );
  AOI222XL \us10/U11  ( .A0(\us10/n185 ), .A1(\us10/n43 ), .B0(\us10/n186 ), 
        .B1(\us10/n187 ), .C0(\us10/n6 ), .C1(\us10/n188 ), .Y(\us10/n164 ) );
  AOI221X1 \us10/U10  ( .A0(\us10/n313 ), .A1(\us10/n5 ), .B0(\us10/n23 ), 
        .B1(\us10/n2 ), .C0(\us10/n328 ), .Y(\us10/n320 ) );
  AOI221X1 \us10/U9  ( .A0(\us10/n40 ), .A1(\us10/n136 ), .B0(\us10/n33 ), 
        .B1(\us10/n178 ), .C0(\us10/n338 ), .Y(\us10/n337 ) );
  AOI222XL \us10/U8  ( .A0(\us10/n278 ), .A1(\us10/n24 ), .B0(\us10/n42 ), 
        .B1(\us10/n33 ), .C0(\us10/n43 ), .C1(\us10/n136 ), .Y(\us10/n351 ) );
  AOI31X1 \us10/U7  ( .A0(sa10[2]), .A1(\us10/n58 ), .A2(sa10[1]), .B0(
        \us10/n40 ), .Y(\us10/n350 ) );
  AOI31X1 \us10/U6  ( .A0(\us10/n44 ), .A1(\us10/n129 ), .A2(\us10/n130 ), 
        .B0(\us10/n131 ), .Y(\us10/n128 ) );
  AOI221X1 \us10/U5  ( .A0(\us10/n40 ), .A1(\us10/n136 ), .B0(\us10/n33 ), 
        .B1(\us10/n47 ), .C0(\us10/n156 ), .Y(\us10/n141 ) );
  OAI32X1 \us10/U4  ( .A0(\us10/n18 ), .A1(sa10[1]), .A2(\us10/n159 ), .B0(
        sa10[4]), .B1(\us10/n182 ), .Y(\us10/n318 ) );
  OAI32X1 \us10/U3  ( .A0(\us10/n210 ), .A1(\us10/n145 ), .A2(\us10/n18 ), 
        .B0(\us10/n27 ), .B1(\us10/n211 ), .Y(\us10/n209 ) );
  AOI221X1 \us10/U2  ( .A0(\us10/n278 ), .A1(\us10/n40 ), .B0(\us10/n185 ), 
        .B1(\us10/n2 ), .C0(\us10/n279 ), .Y(\us10/n273 ) );
  AOI31XL \us10/U1  ( .A0(\us10/n79 ), .A1(\us10/n44 ), .A2(\us10/n2 ), .B0(
        \us10/n280 ), .Y(\us10/n339 ) );
  NAND2X1 \us11/U366  ( .A(\us11/n47 ), .B(\us11/n226 ), .Y(\us11/n189 ) );
  NOR2X1 \us11/U365  ( .A(\us11/n226 ), .B(sa11[3]), .Y(\us11/n242 ) );
  INVX1 \us11/U364  ( .A(\us11/n242 ), .Y(\us11/n205 ) );
  AND2X1 \us11/U363  ( .A(\us11/n189 ), .B(\us11/n205 ), .Y(\us11/n65 ) );
  NOR2X1 \us11/U362  ( .A(\us11/n226 ), .B(\us11/n47 ), .Y(\us11/n45 ) );
  NOR2X1 \us11/U361  ( .A(\us11/n259 ), .B(\us11/n45 ), .Y(\us11/n73 ) );
  NAND2BX1 \us11/U360  ( .AN(\us11/n73 ), .B(\us11/n6 ), .Y(\us11/n158 ) );
  NOR2X1 \us11/U359  ( .A(\us11/n226 ), .B(\us11/n159 ), .Y(\us11/n95 ) );
  INVX1 \us11/U358  ( .A(\us11/n95 ), .Y(\us11/n111 ) );
  NOR2X1 \us11/U357  ( .A(\us11/n145 ), .B(sa11[1]), .Y(\us11/n42 ) );
  INVX1 \us11/U356  ( .A(\us11/n42 ), .Y(\us11/n121 ) );
  INVX1 \us11/U355  ( .A(\us11/n47 ), .Y(\us11/n96 ) );
  OAI211X1 \us11/U354  ( .A0(\us11/n65 ), .A1(\us11/n27 ), .B0(\us11/n158 ), 
        .C0(\us11/n358 ), .Y(\us11/n355 ) );
  NOR2X1 \us11/U353  ( .A(\us11/n226 ), .B(\us11/n145 ), .Y(\us11/n59 ) );
  NOR2X1 \us11/U352  ( .A(\us11/n96 ), .B(\us11/n59 ), .Y(\us11/n271 ) );
  NOR2X1 \us11/U351  ( .A(\us11/n226 ), .B(\us11/n278 ), .Y(\us11/n217 ) );
  INVX1 \us11/U350  ( .A(\us11/n217 ), .Y(\us11/n150 ) );
  NAND2X1 \us11/U349  ( .A(\us11/n44 ), .B(\us11/n150 ), .Y(\us11/n147 ) );
  NAND2X1 \us11/U348  ( .A(sa11[4]), .B(\us11/n226 ), .Y(\us11/n101 ) );
  INVX1 \us11/U347  ( .A(\us11/n159 ), .Y(\us11/n188 ) );
  NOR2X1 \us11/U346  ( .A(\us11/n188 ), .B(\us11/n226 ), .Y(\us11/n25 ) );
  INVX1 \us11/U345  ( .A(\us11/n172 ), .Y(\us11/n107 ) );
  AOI22X1 \us11/U344  ( .A0(\us11/n33 ), .A1(\us11/n147 ), .B0(\us11/n24 ), 
        .B1(\us11/n107 ), .Y(\us11/n357 ) );
  OAI221XL \us11/U343  ( .A0(\us11/n18 ), .A1(\us11/n121 ), .B0(\us11/n271 ), 
        .B1(\us11/n20 ), .C0(\us11/n357 ), .Y(\us11/n356 ) );
  MXI2X1 \us11/U342  ( .A(\us11/n355 ), .B(\us11/n356 ), .S0(\us11/n252 ), .Y(
        \us11/n331 ) );
  INVX1 \us11/U341  ( .A(\us11/n59 ), .Y(\us11/n79 ) );
  AND2X1 \us11/U340  ( .A(\us11/n101 ), .B(\us11/n79 ), .Y(\us11/n325 ) );
  XNOR2X1 \us11/U339  ( .A(sa11[5]), .B(\us11/n226 ), .Y(\us11/n352 ) );
  NOR2X1 \us11/U338  ( .A(\us11/n226 ), .B(\us11/n136 ), .Y(\us11/n281 ) );
  INVX1 \us11/U337  ( .A(\us11/n281 ), .Y(\us11/n19 ) );
  NAND2X1 \us11/U336  ( .A(\us11/n145 ), .B(\us11/n226 ), .Y(\us11/n223 ) );
  AOI21X1 \us11/U335  ( .A0(\us11/n19 ), .A1(\us11/n223 ), .B0(\us11/n27 ), 
        .Y(\us11/n354 ) );
  AOI31X1 \us11/U334  ( .A0(\us11/n6 ), .A1(\us11/n352 ), .A2(\us11/n259 ), 
        .B0(\us11/n354 ), .Y(\us11/n353 ) );
  OAI221XL \us11/U333  ( .A0(\us11/n20 ), .A1(\us11/n34 ), .B0(\us11/n325 ), 
        .B1(\us11/n4 ), .C0(\us11/n353 ), .Y(\us11/n347 ) );
  INVX1 \us11/U332  ( .A(\us11/n352 ), .Y(\us11/n349 ) );
  NAND2X1 \us11/U331  ( .A(\us11/n278 ), .B(\us11/n6 ), .Y(\us11/n74 ) );
  OAI211X1 \us11/U330  ( .A0(\us11/n349 ), .A1(\us11/n74 ), .B0(\us11/n350 ), 
        .C0(\us11/n351 ), .Y(\us11/n348 ) );
  MXI2X1 \us11/U329  ( .A(\us11/n347 ), .B(\us11/n348 ), .S0(\us11/n252 ), .Y(
        \us11/n332 ) );
  NOR2X1 \us11/U328  ( .A(\us11/n44 ), .B(\us11/n226 ), .Y(\us11/n157 ) );
  INVX1 \us11/U327  ( .A(\us11/n157 ), .Y(\us11/n240 ) );
  NAND2X1 \us11/U326  ( .A(\us11/n240 ), .B(\us11/n189 ), .Y(\us11/n68 ) );
  NOR2X1 \us11/U325  ( .A(\us11/n20 ), .B(\us11/n159 ), .Y(\us11/n225 ) );
  NOR2X1 \us11/U324  ( .A(\us11/n225 ), .B(\us11/n40 ), .Y(\us11/n345 ) );
  INVX1 \us11/U323  ( .A(\us11/n278 ), .Y(\us11/n94 ) );
  NAND2X1 \us11/U322  ( .A(\us11/n94 ), .B(\us11/n226 ), .Y(\us11/n199 ) );
  NAND2X1 \us11/U321  ( .A(\us11/n199 ), .B(\us11/n205 ), .Y(\us11/n82 ) );
  NAND2X1 \us11/U320  ( .A(\us11/n19 ), .B(\us11/n199 ), .Y(\us11/n295 ) );
  NOR2X1 \us11/U319  ( .A(\us11/n226 ), .B(\us11/n259 ), .Y(\us11/n210 ) );
  NOR2X1 \us11/U318  ( .A(\us11/n27 ), .B(\us11/n210 ), .Y(\us11/n173 ) );
  MXI2X1 \us11/U317  ( .A(\us11/n345 ), .B(\us11/n346 ), .S0(\us11/n252 ), .Y(
        \us11/n342 ) );
  NOR2X1 \us11/U316  ( .A(sa11[1]), .B(sa11[3]), .Y(\us11/n163 ) );
  INVX1 \us11/U315  ( .A(\us11/n163 ), .Y(\us11/n37 ) );
  INVX1 \us11/U314  ( .A(\us11/n173 ), .Y(\us11/n344 ) );
  AOI21X1 \us11/U313  ( .A0(\us11/n240 ), .A1(\us11/n37 ), .B0(\us11/n344 ), 
        .Y(\us11/n343 ) );
  AOI211X1 \us11/U312  ( .A0(\us11/n5 ), .A1(\us11/n68 ), .B0(\us11/n342 ), 
        .C0(\us11/n343 ), .Y(\us11/n333 ) );
  NOR2X1 \us11/U311  ( .A(\us11/n18 ), .B(\us11/n226 ), .Y(\us11/n258 ) );
  NAND2X1 \us11/U310  ( .A(\us11/n278 ), .B(sa11[1]), .Y(\us11/n204 ) );
  NOR2X1 \us11/U309  ( .A(\us11/n188 ), .B(sa11[1]), .Y(\us11/n179 ) );
  INVX1 \us11/U308  ( .A(\us11/n179 ), .Y(\us11/n330 ) );
  NAND2X1 \us11/U307  ( .A(\us11/n204 ), .B(\us11/n330 ), .Y(\us11/n239 ) );
  NOR2X1 \us11/U306  ( .A(\us11/n136 ), .B(sa11[1]), .Y(\us11/n299 ) );
  NOR2X1 \us11/U305  ( .A(\us11/n299 ), .B(\us11/n210 ), .Y(\us11/n341 ) );
  OAI32X1 \us11/U304  ( .A0(\us11/n27 ), .A1(\us11/n278 ), .A2(\us11/n95 ), 
        .B0(\us11/n341 ), .B1(\us11/n4 ), .Y(\us11/n340 ) );
  INVX1 \us11/U303  ( .A(\us11/n45 ), .Y(\us11/n126 ) );
  NAND2X1 \us11/U302  ( .A(\us11/n126 ), .B(\us11/n101 ), .Y(\us11/n178 ) );
  NOR2X1 \us11/U301  ( .A(\us11/n18 ), .B(\us11/n136 ), .Y(\us11/n280 ) );
  OAI21XL \us11/U300  ( .A0(\us11/n4 ), .A1(\us11/n121 ), .B0(\us11/n339 ), 
        .Y(\us11/n338 ) );
  MXI2X1 \us11/U299  ( .A(\us11/n336 ), .B(\us11/n337 ), .S0(\us11/n252 ), .Y(
        \us11/n335 ) );
  NOR2X1 \us11/U298  ( .A(\us11/n258 ), .B(\us11/n335 ), .Y(\us11/n334 ) );
  MX4X1 \us11/U297  ( .A(\us11/n331 ), .B(\us11/n332 ), .C(\us11/n333 ), .D(
        \us11/n334 ), .S0(sa11[6]), .S1(\us11/n234 ), .Y(sa10_sr[0]) );
  INVX1 \us11/U296  ( .A(\us11/n299 ), .Y(\us11/n80 ) );
  NOR2X1 \us11/U295  ( .A(\us11/n111 ), .B(\us11/n18 ), .Y(\us11/n269 ) );
  INVX1 \us11/U294  ( .A(\us11/n269 ), .Y(\us11/n75 ) );
  OAI221XL \us11/U293  ( .A0(\us11/n18 ), .A1(\us11/n330 ), .B0(\us11/n20 ), 
        .B1(\us11/n80 ), .C0(\us11/n75 ), .Y(\us11/n329 ) );
  AOI221X1 \us11/U292  ( .A0(\us11/n325 ), .A1(\us11/n33 ), .B0(\us11/n24 ), 
        .B1(\us11/n303 ), .C0(\us11/n329 ), .Y(\us11/n319 ) );
  NOR2X1 \us11/U291  ( .A(\us11/n234 ), .B(sa11[5]), .Y(\us11/n14 ) );
  NOR2X1 \us11/U290  ( .A(\us11/n25 ), .B(\us11/n299 ), .Y(\us11/n313 ) );
  NAND2X1 \us11/U289  ( .A(\us11/n44 ), .B(\us11/n226 ), .Y(\us11/n300 ) );
  AND2X1 \us11/U288  ( .A(\us11/n300 ), .B(\us11/n240 ), .Y(\us11/n23 ) );
  OAI32X1 \us11/U287  ( .A0(\us11/n4 ), .A1(\us11/n145 ), .A2(\us11/n210 ), 
        .B0(\us11/n137 ), .B1(\us11/n27 ), .Y(\us11/n328 ) );
  NOR2X1 \us11/U286  ( .A(sa11[0]), .B(sa11[5]), .Y(\us11/n16 ) );
  INVX1 \us11/U285  ( .A(\us11/n16 ), .Y(\us11/n114 ) );
  INVX1 \us11/U284  ( .A(\us11/n145 ), .Y(\us11/n149 ) );
  NOR2X1 \us11/U283  ( .A(\us11/n47 ), .B(sa11[1]), .Y(\us11/n98 ) );
  INVX1 \us11/U282  ( .A(\us11/n98 ), .Y(\us11/n284 ) );
  OAI21XL \us11/U281  ( .A0(\us11/n69 ), .A1(\us11/n284 ), .B0(\us11/n27 ), 
        .Y(\us11/n327 ) );
  AOI31X1 \us11/U280  ( .A0(\us11/n111 ), .A1(\us11/n149 ), .A2(\us11/n327 ), 
        .B0(\us11/n225 ), .Y(\us11/n326 ) );
  OAI21XL \us11/U279  ( .A0(\us11/n325 ), .A1(\us11/n18 ), .B0(\us11/n326 ), 
        .Y(\us11/n322 ) );
  NAND2X1 \us11/U278  ( .A(\us11/n19 ), .B(\us11/n189 ), .Y(\us11/n71 ) );
  NOR2X1 \us11/U277  ( .A(\us11/n71 ), .B(\us11/n18 ), .Y(\us11/n135 ) );
  AOI21X1 \us11/U276  ( .A0(\us11/n40 ), .A1(sa11[4]), .B0(\us11/n135 ), .Y(
        \us11/n324 ) );
  OAI221XL \us11/U275  ( .A0(\us11/n47 ), .A1(\us11/n27 ), .B0(\us11/n65 ), 
        .B1(\us11/n20 ), .C0(\us11/n324 ), .Y(\us11/n323 ) );
  AOI22X1 \us11/U274  ( .A0(\us11/n55 ), .A1(\us11/n322 ), .B0(\us11/n89 ), 
        .B1(\us11/n323 ), .Y(\us11/n321 ) );
  OAI221XL \us11/U273  ( .A0(\us11/n319 ), .A1(\us11/n52 ), .B0(\us11/n320 ), 
        .B1(\us11/n114 ), .C0(\us11/n321 ), .Y(\us11/n304 ) );
  NOR2X1 \us11/U272  ( .A(\us11/n226 ), .B(\us11/n58 ), .Y(\us11/n290 ) );
  INVX1 \us11/U271  ( .A(\us11/n290 ), .Y(\us11/n200 ) );
  NAND2X1 \us11/U270  ( .A(\us11/n34 ), .B(\us11/n200 ), .Y(\us11/n120 ) );
  INVX1 \us11/U269  ( .A(\us11/n210 ), .Y(\us11/n100 ) );
  OAI221XL \us11/U268  ( .A0(\us11/n20 ), .A1(\us11/n100 ), .B0(sa11[3]), .B1(
        \us11/n4 ), .C0(\us11/n262 ), .Y(\us11/n317 ) );
  INVX1 \us11/U267  ( .A(\us11/n258 ), .Y(\us11/n182 ) );
  AOI211X1 \us11/U266  ( .A0(\us11/n33 ), .A1(\us11/n120 ), .B0(\us11/n317 ), 
        .C0(\us11/n318 ), .Y(\us11/n306 ) );
  NAND2X1 \us11/U265  ( .A(\us11/n100 ), .B(\us11/n199 ), .Y(\us11/n151 ) );
  INVX1 \us11/U264  ( .A(\us11/n151 ), .Y(\us11/n314 ) );
  NOR2X1 \us11/U263  ( .A(\us11/n45 ), .B(\us11/n163 ), .Y(\us11/n160 ) );
  INVX1 \us11/U262  ( .A(\us11/n295 ), .Y(\us11/n92 ) );
  AOI21X1 \us11/U261  ( .A0(sa11[1]), .A1(\us11/n58 ), .B0(\us11/n98 ), .Y(
        \us11/n316 ) );
  OAI22X1 \us11/U260  ( .A0(\us11/n92 ), .A1(\us11/n18 ), .B0(\us11/n316 ), 
        .B1(\us11/n27 ), .Y(\us11/n315 ) );
  NOR2X1 \us11/U259  ( .A(\us11/n149 ), .B(\us11/n226 ), .Y(\us11/n41 ) );
  INVX1 \us11/U258  ( .A(\us11/n41 ), .Y(\us11/n105 ) );
  NAND2X1 \us11/U257  ( .A(\us11/n284 ), .B(\us11/n105 ), .Y(\us11/n227 ) );
  AOI21X1 \us11/U256  ( .A0(\us11/n313 ), .A1(\us11/n33 ), .B0(\us11/n269 ), 
        .Y(\us11/n312 ) );
  OAI221XL \us11/U255  ( .A0(\us11/n149 ), .A1(\us11/n20 ), .B0(\us11/n4 ), 
        .B1(\us11/n227 ), .C0(\us11/n312 ), .Y(\us11/n309 ) );
  AOI21X1 \us11/U254  ( .A0(\us11/n226 ), .A1(\us11/n188 ), .B0(\us11/n242 ), 
        .Y(\us11/n185 ) );
  INVX1 \us11/U253  ( .A(\us11/n185 ), .Y(\us11/n48 ) );
  AND2X1 \us11/U252  ( .A(\us11/n223 ), .B(\us11/n240 ), .Y(\us11/n28 ) );
  OAI221XL \us11/U251  ( .A0(\us11/n27 ), .A1(\us11/n44 ), .B0(\us11/n4 ), 
        .B1(\us11/n48 ), .C0(\us11/n311 ), .Y(\us11/n310 ) );
  AOI22X1 \us11/U250  ( .A0(\us11/n89 ), .A1(\us11/n309 ), .B0(\us11/n55 ), 
        .B1(\us11/n310 ), .Y(\us11/n308 ) );
  OAI221XL \us11/U249  ( .A0(\us11/n306 ), .A1(\us11/n52 ), .B0(\us11/n307 ), 
        .B1(\us11/n114 ), .C0(\us11/n308 ), .Y(\us11/n305 ) );
  MX2X1 \us11/U248  ( .A(\us11/n304 ), .B(\us11/n305 ), .S0(sa11[6]), .Y(
        sa10_sr[1]) );
  INVX1 \us11/U247  ( .A(\us11/n187 ), .Y(\us11/n61 ) );
  MXI2X1 \us11/U246  ( .A(\us11/n303 ), .B(\us11/n61 ), .S0(\us11/n69 ), .Y(
        \us11/n301 ) );
  MXI2X1 \us11/U245  ( .A(\us11/n301 ), .B(\us11/n147 ), .S0(\us11/n302 ), .Y(
        \us11/n285 ) );
  NAND2X1 \us11/U244  ( .A(\us11/n200 ), .B(\us11/n300 ), .Y(\us11/n99 ) );
  INVX1 \us11/U243  ( .A(\us11/n99 ), .Y(\us11/n296 ) );
  NOR2X1 \us11/U242  ( .A(\us11/n299 ), .B(\us11/n242 ), .Y(\us11/n298 ) );
  NAND2X1 \us11/U241  ( .A(sa11[1]), .B(\us11/n47 ), .Y(\us11/n122 ) );
  NOR2X1 \us11/U240  ( .A(\us11/n159 ), .B(\us11/n217 ), .Y(\us11/n198 ) );
  OAI221XL \us11/U239  ( .A0(\us11/n298 ), .A1(\us11/n27 ), .B0(\us11/n20 ), 
        .B1(\us11/n122 ), .C0(\us11/n132 ), .Y(\us11/n297 ) );
  AOI221X1 \us11/U238  ( .A0(\us11/n225 ), .A1(\us11/n226 ), .B0(\us11/n296 ), 
        .B1(\us11/n6 ), .C0(\us11/n297 ), .Y(\us11/n291 ) );
  OAI2BB2X1 \us11/U237  ( .B0(\us11/n27 ), .B1(\us11/n295 ), .A0N(\us11/n34 ), 
        .A1N(\us11/n24 ), .Y(\us11/n293 ) );
  AOI21X1 \us11/U236  ( .A0(\us11/n101 ), .A1(\us11/n150 ), .B0(\us11/n20 ), 
        .Y(\us11/n294 ) );
  AOI211X1 \us11/U235  ( .A0(\us11/n5 ), .A1(\us11/n79 ), .B0(\us11/n293 ), 
        .C0(\us11/n294 ), .Y(\us11/n292 ) );
  INVX1 \us11/U234  ( .A(\us11/n89 ), .Y(\us11/n10 ) );
  OAI22X1 \us11/U233  ( .A0(\us11/n291 ), .A1(\us11/n114 ), .B0(\us11/n292 ), 
        .B1(\us11/n10 ), .Y(\us11/n286 ) );
  INVX1 \us11/U232  ( .A(\us11/n225 ), .Y(\us11/n288 ) );
  NAND2X1 \us11/U231  ( .A(\us11/n200 ), .B(\us11/n284 ), .Y(\us11/n102 ) );
  NOR2X1 \us11/U230  ( .A(\us11/n290 ), .B(\us11/n163 ), .Y(\us11/n184 ) );
  AOI22X1 \us11/U229  ( .A0(\us11/n102 ), .A1(\us11/n69 ), .B0(\us11/n184 ), 
        .B1(\us11/n33 ), .Y(\us11/n289 ) );
  AOI31X1 \us11/U228  ( .A0(\us11/n132 ), .A1(\us11/n288 ), .A2(\us11/n289 ), 
        .B0(\us11/n52 ), .Y(\us11/n287 ) );
  AOI211X1 \us11/U227  ( .A0(\us11/n285 ), .A1(\us11/n55 ), .B0(\us11/n286 ), 
        .C0(\us11/n287 ), .Y(\us11/n263 ) );
  NAND2X1 \us11/U226  ( .A(\us11/n284 ), .B(\us11/n122 ), .Y(\us11/n125 ) );
  NOR2X1 \us11/U225  ( .A(\us11/n199 ), .B(\us11/n4 ), .Y(\us11/n50 ) );
  AOI21X1 \us11/U224  ( .A0(\us11/n200 ), .A1(\us11/n223 ), .B0(\us11/n20 ), 
        .Y(\us11/n283 ) );
  AOI211X1 \us11/U223  ( .A0(\us11/n5 ), .A1(\us11/n125 ), .B0(\us11/n50 ), 
        .C0(\us11/n283 ), .Y(\us11/n282 ) );
  OAI221XL \us11/U222  ( .A0(\us11/n281 ), .A1(\us11/n27 ), .B0(\us11/n4 ), 
        .B1(\us11/n111 ), .C0(\us11/n282 ), .Y(\us11/n265 ) );
  INVX1 \us11/U221  ( .A(\us11/n280 ), .Y(\us11/n247 ) );
  NAND2X1 \us11/U220  ( .A(\us11/n41 ), .B(\us11/n33 ), .Y(\us11/n272 ) );
  OAI221XL \us11/U219  ( .A0(sa11[1]), .A1(\us11/n247 ), .B0(\us11/n4 ), .B1(
        \us11/n189 ), .C0(\us11/n272 ), .Y(\us11/n279 ) );
  NAND2X1 \us11/U218  ( .A(sa11[2]), .B(\us11/n149 ), .Y(\us11/n276 ) );
  XNOR2X1 \us11/U217  ( .A(\us11/n129 ), .B(sa11[1]), .Y(\us11/n155 ) );
  MXI2X1 \us11/U216  ( .A(\us11/n276 ), .B(\us11/n277 ), .S0(\us11/n155 ), .Y(
        \us11/n275 ) );
  OAI22X1 \us11/U215  ( .A0(\us11/n273 ), .A1(\us11/n10 ), .B0(\us11/n274 ), 
        .B1(\us11/n52 ), .Y(\us11/n266 ) );
  NOR2X1 \us11/U214  ( .A(\us11/n20 ), .B(\us11/n226 ), .Y(\us11/n176 ) );
  OAI21XL \us11/U213  ( .A0(\us11/n4 ), .A1(\us11/n271 ), .B0(\us11/n272 ), 
        .Y(\us11/n270 ) );
  OAI31X1 \us11/U212  ( .A0(\us11/n176 ), .A1(\us11/n269 ), .A2(\us11/n270 ), 
        .B0(\us11/n16 ), .Y(\us11/n268 ) );
  INVX1 \us11/U211  ( .A(\us11/n268 ), .Y(\us11/n267 ) );
  AOI211X1 \us11/U210  ( .A0(\us11/n55 ), .A1(\us11/n265 ), .B0(\us11/n266 ), 
        .C0(\us11/n267 ), .Y(\us11/n264 ) );
  MXI2X1 \us11/U209  ( .A(\us11/n263 ), .B(\us11/n264 ), .S0(sa11[6]), .Y(
        sa10_sr[2]) );
  NOR2X1 \us11/U208  ( .A(\us11/n94 ), .B(sa11[1]), .Y(\us11/n211 ) );
  INVX1 \us11/U207  ( .A(\us11/n262 ), .Y(\us11/n261 ) );
  AOI211X1 \us11/U206  ( .A0(\us11/n259 ), .A1(\us11/n24 ), .B0(\us11/n260 ), 
        .C0(\us11/n261 ), .Y(\us11/n255 ) );
  OAI22X1 \us11/U205  ( .A0(\us11/n20 ), .A1(\us11/n68 ), .B0(\us11/n27 ), 
        .B1(\us11/n37 ), .Y(\us11/n257 ) );
  NOR3X1 \us11/U204  ( .A(\us11/n257 ), .B(\us11/n258 ), .C(\us11/n50 ), .Y(
        \us11/n256 ) );
  MXI2X1 \us11/U203  ( .A(\us11/n255 ), .B(\us11/n256 ), .S0(\us11/n252 ), .Y(
        \us11/n254 ) );
  AOI221X1 \us11/U202  ( .A0(\us11/n211 ), .A1(\us11/n5 ), .B0(\us11/n40 ), 
        .B1(sa11[4]), .C0(\us11/n254 ), .Y(\us11/n248 ) );
  INVX1 \us11/U201  ( .A(\us11/n211 ), .Y(\us11/n106 ) );
  NAND2X1 \us11/U200  ( .A(\us11/n200 ), .B(\us11/n106 ), .Y(\us11/n83 ) );
  NAND2X1 \us11/U199  ( .A(\us11/n199 ), .B(\us11/n204 ), .Y(\us11/n169 ) );
  AOI2BB2X1 \us11/U198  ( .B0(\us11/n65 ), .B1(\us11/n24 ), .A0N(\us11/n169 ), 
        .A1N(\us11/n20 ), .Y(\us11/n253 ) );
  OAI221XL \us11/U197  ( .A0(\us11/n172 ), .A1(\us11/n18 ), .B0(\us11/n27 ), 
        .B1(\us11/n83 ), .C0(\us11/n253 ), .Y(\us11/n251 ) );
  MXI2X1 \us11/U196  ( .A(\us11/n250 ), .B(\us11/n251 ), .S0(\us11/n252 ), .Y(
        \us11/n249 ) );
  MXI2X1 \us11/U195  ( .A(\us11/n248 ), .B(\us11/n249 ), .S0(\us11/n234 ), .Y(
        \us11/n228 ) );
  OAI21XL \us11/U194  ( .A0(\us11/n58 ), .A1(\us11/n27 ), .B0(\us11/n247 ), 
        .Y(\us11/n245 ) );
  NOR2X1 \us11/U193  ( .A(sa11[7]), .B(\us11/n145 ), .Y(\us11/n246 ) );
  XNOR2X1 \us11/U192  ( .A(\us11/n69 ), .B(sa11[1]), .Y(\us11/n130 ) );
  MXI2X1 \us11/U191  ( .A(\us11/n245 ), .B(\us11/n246 ), .S0(\us11/n130 ), .Y(
        \us11/n243 ) );
  OAI211X1 \us11/U190  ( .A0(\us11/n4 ), .A1(\us11/n149 ), .B0(\us11/n243 ), 
        .C0(\us11/n244 ), .Y(\us11/n230 ) );
  NOR2X1 \us11/U189  ( .A(\us11/n242 ), .B(\us11/n137 ), .Y(\us11/n70 ) );
  OAI221XL \us11/U188  ( .A0(\us11/n159 ), .A1(\us11/n27 ), .B0(\us11/n20 ), 
        .B1(\us11/n34 ), .C0(\us11/n241 ), .Y(\us11/n231 ) );
  NAND2X1 \us11/U187  ( .A(\us11/n101 ), .B(\us11/n240 ), .Y(\us11/n76 ) );
  AOI21X1 \us11/U186  ( .A0(\us11/n122 ), .A1(\us11/n106 ), .B0(\us11/n129 ), 
        .Y(\us11/n237 ) );
  INVX1 \us11/U185  ( .A(\us11/n239 ), .Y(\us11/n238 ) );
  OAI21XL \us11/U184  ( .A0(\us11/n237 ), .A1(\us11/n43 ), .B0(\us11/n238 ), 
        .Y(\us11/n236 ) );
  OAI221XL \us11/U183  ( .A0(\us11/n18 ), .A1(\us11/n76 ), .B0(\us11/n59 ), 
        .B1(\us11/n27 ), .C0(\us11/n236 ), .Y(\us11/n232 ) );
  AOI2BB2X1 \us11/U182  ( .B0(\us11/n24 ), .B1(\us11/n187 ), .A0N(\us11/n227 ), 
        .A1N(\us11/n20 ), .Y(\us11/n235 ) );
  OAI211X1 \us11/U181  ( .A0(\us11/n27 ), .A1(\us11/n122 ), .B0(\us11/n158 ), 
        .C0(\us11/n235 ), .Y(\us11/n233 ) );
  MX4X1 \us11/U180  ( .A(\us11/n230 ), .B(\us11/n231 ), .C(\us11/n232 ), .D(
        \us11/n233 ), .S0(\us11/n234 ), .S1(sa11[5]), .Y(\us11/n229 ) );
  MX2X1 \us11/U179  ( .A(\us11/n228 ), .B(\us11/n229 ), .S0(sa11[6]), .Y(
        sa10_sr[3]) );
  NOR2BX1 \us11/U178  ( .AN(\us11/n204 ), .B(\us11/n137 ), .Y(\us11/n110 ) );
  INVX1 \us11/U177  ( .A(\us11/n110 ), .Y(\us11/n64 ) );
  AOI22X1 \us11/U176  ( .A0(\us11/n225 ), .A1(\us11/n226 ), .B0(\us11/n6 ), 
        .B1(\us11/n227 ), .Y(\us11/n224 ) );
  OAI221XL \us11/U175  ( .A0(\us11/n27 ), .A1(\us11/n64 ), .B0(\us11/n4 ), 
        .B1(\us11/n83 ), .C0(\us11/n224 ), .Y(\us11/n212 ) );
  NAND2X1 \us11/U174  ( .A(\us11/n34 ), .B(\us11/n204 ), .Y(\us11/n221 ) );
  OAI21XL \us11/U173  ( .A0(\us11/n69 ), .A1(\us11/n223 ), .B0(\us11/n27 ), 
        .Y(\us11/n222 ) );
  NOR2X1 \us11/U172  ( .A(\us11/n217 ), .B(\us11/n42 ), .Y(\us11/n208 ) );
  AOI211X1 \us11/U171  ( .A0(\us11/n208 ), .A1(\us11/n5 ), .B0(\us11/n220 ), 
        .C0(\us11/n173 ), .Y(\us11/n219 ) );
  OAI22X1 \us11/U170  ( .A0(\us11/n218 ), .A1(\us11/n10 ), .B0(\us11/n219 ), 
        .B1(\us11/n114 ), .Y(\us11/n213 ) );
  INVX1 \us11/U169  ( .A(\us11/n135 ), .Y(\us11/n215 ) );
  NOR2X1 \us11/U168  ( .A(\us11/n4 ), .B(\us11/n159 ), .Y(\us11/n31 ) );
  INVX1 \us11/U167  ( .A(\us11/n31 ), .Y(\us11/n196 ) );
  AOI31X1 \us11/U166  ( .A0(\us11/n215 ), .A1(\us11/n196 ), .A2(\us11/n216 ), 
        .B0(\us11/n52 ), .Y(\us11/n214 ) );
  AOI211X1 \us11/U165  ( .A0(\us11/n55 ), .A1(\us11/n212 ), .B0(\us11/n213 ), 
        .C0(\us11/n214 ), .Y(\us11/n190 ) );
  INVX1 \us11/U164  ( .A(\us11/n207 ), .Y(\us11/n192 ) );
  NOR2X1 \us11/U163  ( .A(\us11/n25 ), .B(\us11/n98 ), .Y(\us11/n32 ) );
  OAI22X1 \us11/U162  ( .A0(\us11/n28 ), .A1(\us11/n4 ), .B0(\us11/n188 ), 
        .B1(\us11/n27 ), .Y(\us11/n206 ) );
  NAND2X1 \us11/U161  ( .A(\us11/n204 ), .B(\us11/n80 ), .Y(\us11/n118 ) );
  INVX1 \us11/U160  ( .A(\us11/n118 ), .Y(\us11/n123 ) );
  NAND2X1 \us11/U159  ( .A(\us11/n94 ), .B(\us11/n79 ), .Y(\us11/n203 ) );
  OAI2BB1X1 \us11/U158  ( .A0N(\us11/n199 ), .A1N(\us11/n200 ), .B0(\us11/n33 ), .Y(\us11/n195 ) );
  INVX1 \us11/U157  ( .A(\us11/n55 ), .Y(\us11/n12 ) );
  AOI31X1 \us11/U156  ( .A0(\us11/n195 ), .A1(\us11/n196 ), .A2(\us11/n197 ), 
        .B0(\us11/n12 ), .Y(\us11/n194 ) );
  AOI211X1 \us11/U155  ( .A0(\us11/n89 ), .A1(\us11/n192 ), .B0(\us11/n193 ), 
        .C0(\us11/n194 ), .Y(\us11/n191 ) );
  MXI2X1 \us11/U154  ( .A(\us11/n190 ), .B(\us11/n191 ), .S0(sa11[6]), .Y(
        sa10_sr[4]) );
  OAI21XL \us11/U153  ( .A0(\us11/n69 ), .A1(\us11/n189 ), .B0(\us11/n27 ), 
        .Y(\us11/n186 ) );
  INVX1 \us11/U152  ( .A(\us11/n183 ), .Y(\us11/n180 ) );
  NAND2X1 \us11/U151  ( .A(\us11/n74 ), .B(\us11/n182 ), .Y(\us11/n181 ) );
  AOI211X1 \us11/U150  ( .A0(\us11/n179 ), .A1(\us11/n24 ), .B0(\us11/n180 ), 
        .C0(\us11/n181 ), .Y(\us11/n165 ) );
  INVX1 \us11/U149  ( .A(\us11/n178 ), .Y(\us11/n175 ) );
  AOI211X1 \us11/U148  ( .A0(\us11/n175 ), .A1(\us11/n5 ), .B0(\us11/n176 ), 
        .C0(\us11/n177 ), .Y(\us11/n174 ) );
  OAI221XL \us11/U147  ( .A0(\us11/n159 ), .A1(\us11/n27 ), .B0(\us11/n145 ), 
        .B1(\us11/n20 ), .C0(\us11/n174 ), .Y(\us11/n167 ) );
  MXI2X1 \us11/U146  ( .A(\us11/n40 ), .B(\us11/n173 ), .S0(\us11/n96 ), .Y(
        \us11/n170 ) );
  AOI22X1 \us11/U145  ( .A0(\us11/n137 ), .A1(\us11/n24 ), .B0(\us11/n172 ), 
        .B1(\us11/n6 ), .Y(\us11/n171 ) );
  OAI211X1 \us11/U144  ( .A0(\us11/n20 ), .A1(\us11/n169 ), .B0(\us11/n170 ), 
        .C0(\us11/n171 ), .Y(\us11/n168 ) );
  AOI22X1 \us11/U143  ( .A0(\us11/n89 ), .A1(\us11/n167 ), .B0(\us11/n55 ), 
        .B1(\us11/n168 ), .Y(\us11/n166 ) );
  OAI221XL \us11/U142  ( .A0(\us11/n164 ), .A1(\us11/n114 ), .B0(\us11/n165 ), 
        .B1(\us11/n52 ), .C0(\us11/n166 ), .Y(\us11/n138 ) );
  OAI21XL \us11/U141  ( .A0(\us11/n41 ), .A1(\us11/n163 ), .B0(\us11/n69 ), 
        .Y(\us11/n162 ) );
  AOI221X1 \us11/U140  ( .A0(\us11/n159 ), .A1(\us11/n24 ), .B0(\us11/n160 ), 
        .B1(\us11/n33 ), .C0(\us11/n161 ), .Y(\us11/n140 ) );
  OAI21XL \us11/U139  ( .A0(\us11/n157 ), .A1(\us11/n20 ), .B0(\us11/n158 ), 
        .Y(\us11/n156 ) );
  NOR2X1 \us11/U138  ( .A(\us11/n4 ), .B(\us11/n136 ), .Y(\us11/n153 ) );
  NOR2X1 \us11/U137  ( .A(\us11/n145 ), .B(\us11/n69 ), .Y(\us11/n154 ) );
  MXI2X1 \us11/U136  ( .A(\us11/n153 ), .B(\us11/n154 ), .S0(\us11/n155 ), .Y(
        \us11/n152 ) );
  OAI221XL \us11/U135  ( .A0(\us11/n110 ), .A1(\us11/n18 ), .B0(\us11/n20 ), 
        .B1(\us11/n151 ), .C0(\us11/n152 ), .Y(\us11/n143 ) );
  AOI21X1 \us11/U134  ( .A0(\us11/n149 ), .A1(\us11/n150 ), .B0(\us11/n18 ), 
        .Y(\us11/n148 ) );
  AOI2BB1X1 \us11/U133  ( .A0N(\us11/n147 ), .A1N(\us11/n27 ), .B0(\us11/n148 ), .Y(\us11/n146 ) );
  OAI221XL \us11/U132  ( .A0(\us11/n145 ), .A1(\us11/n20 ), .B0(\us11/n4 ), 
        .B1(\us11/n34 ), .C0(\us11/n146 ), .Y(\us11/n144 ) );
  AOI22X1 \us11/U131  ( .A0(\us11/n89 ), .A1(\us11/n143 ), .B0(\us11/n14 ), 
        .B1(\us11/n144 ), .Y(\us11/n142 ) );
  OAI221XL \us11/U130  ( .A0(\us11/n140 ), .A1(\us11/n12 ), .B0(\us11/n141 ), 
        .B1(\us11/n114 ), .C0(\us11/n142 ), .Y(\us11/n139 ) );
  MX2X1 \us11/U129  ( .A(\us11/n138 ), .B(\us11/n139 ), .S0(sa11[6]), .Y(
        sa10_sr[5]) );
  INVX1 \us11/U128  ( .A(\us11/n70 ), .Y(\us11/n133 ) );
  OAI22X1 \us11/U127  ( .A0(\us11/n4 ), .A1(\us11/n136 ), .B0(\us11/n137 ), 
        .B1(\us11/n27 ), .Y(\us11/n134 ) );
  AOI211X1 \us11/U126  ( .A0(\us11/n133 ), .A1(\us11/n69 ), .B0(\us11/n134 ), 
        .C0(\us11/n135 ), .Y(\us11/n112 ) );
  INVX1 \us11/U125  ( .A(\us11/n132 ), .Y(\us11/n131 ) );
  OAI21XL \us11/U124  ( .A0(\us11/n18 ), .A1(\us11/n37 ), .B0(\us11/n128 ), 
        .Y(\us11/n127 ) );
  OAI221XL \us11/U123  ( .A0(\us11/n18 ), .A1(\us11/n105 ), .B0(\us11/n123 ), 
        .B1(\us11/n27 ), .C0(\us11/n124 ), .Y(\us11/n116 ) );
  NAND2X1 \us11/U122  ( .A(\us11/n121 ), .B(\us11/n122 ), .Y(\us11/n30 ) );
  OAI221XL \us11/U121  ( .A0(\us11/n18 ), .A1(\us11/n118 ), .B0(\us11/n27 ), 
        .B1(\us11/n30 ), .C0(\us11/n119 ), .Y(\us11/n117 ) );
  AOI22X1 \us11/U120  ( .A0(\us11/n89 ), .A1(\us11/n116 ), .B0(\us11/n55 ), 
        .B1(\us11/n117 ), .Y(\us11/n115 ) );
  OAI221XL \us11/U119  ( .A0(\us11/n112 ), .A1(\us11/n52 ), .B0(\us11/n113 ), 
        .B1(\us11/n114 ), .C0(\us11/n115 ), .Y(\us11/n84 ) );
  OAI22X1 \us11/U118  ( .A0(\us11/n110 ), .A1(\us11/n4 ), .B0(\us11/n20 ), 
        .B1(\us11/n21 ), .Y(\us11/n108 ) );
  AOI21X1 \us11/U117  ( .A0(sa11[1]), .A1(\us11/n58 ), .B0(\us11/n27 ), .Y(
        \us11/n109 ) );
  AOI211X1 \us11/U116  ( .A0(\us11/n5 ), .A1(\us11/n107 ), .B0(\us11/n108 ), 
        .C0(\us11/n109 ), .Y(\us11/n86 ) );
  OAI22X1 \us11/U115  ( .A0(\us11/n45 ), .A1(\us11/n4 ), .B0(sa11[4]), .B1(
        \us11/n18 ), .Y(\us11/n103 ) );
  AOI21X1 \us11/U114  ( .A0(\us11/n105 ), .A1(\us11/n106 ), .B0(\us11/n20 ), 
        .Y(\us11/n104 ) );
  AOI211X1 \us11/U113  ( .A0(\us11/n33 ), .A1(\us11/n102 ), .B0(\us11/n103 ), 
        .C0(\us11/n104 ), .Y(\us11/n87 ) );
  NAND2X1 \us11/U112  ( .A(\us11/n100 ), .B(\us11/n101 ), .Y(\us11/n62 ) );
  OAI221XL \us11/U111  ( .A0(\us11/n27 ), .A1(\us11/n62 ), .B0(\us11/n4 ), 
        .B1(\us11/n21 ), .C0(\us11/n97 ), .Y(\us11/n90 ) );
  NOR3X1 \us11/U110  ( .A(\us11/n4 ), .B(\us11/n95 ), .C(\us11/n96 ), .Y(
        \us11/n67 ) );
  AOI31X1 \us11/U109  ( .A0(\us11/n79 ), .A1(\us11/n94 ), .A2(\us11/n6 ), .B0(
        \us11/n67 ), .Y(\us11/n93 ) );
  OAI221XL \us11/U108  ( .A0(\us11/n73 ), .A1(\us11/n27 ), .B0(\us11/n92 ), 
        .B1(\us11/n20 ), .C0(\us11/n93 ), .Y(\us11/n91 ) );
  AOI22X1 \us11/U107  ( .A0(\us11/n89 ), .A1(\us11/n90 ), .B0(\us11/n16 ), 
        .B1(\us11/n91 ), .Y(\us11/n88 ) );
  OAI221XL \us11/U106  ( .A0(\us11/n86 ), .A1(\us11/n52 ), .B0(\us11/n87 ), 
        .B1(\us11/n12 ), .C0(\us11/n88 ), .Y(\us11/n85 ) );
  MX2X1 \us11/U105  ( .A(\us11/n84 ), .B(\us11/n85 ), .S0(sa11[6]), .Y(
        sa10_sr[6]) );
  INVX1 \us11/U104  ( .A(\us11/n81 ), .Y(\us11/n77 ) );
  AOI21X1 \us11/U103  ( .A0(\us11/n79 ), .A1(\us11/n80 ), .B0(\us11/n27 ), .Y(
        \us11/n78 ) );
  AOI211X1 \us11/U102  ( .A0(\us11/n5 ), .A1(\us11/n76 ), .B0(\us11/n77 ), 
        .C0(\us11/n78 ), .Y(\us11/n51 ) );
  OAI211X1 \us11/U101  ( .A0(\us11/n73 ), .A1(\us11/n27 ), .B0(\us11/n74 ), 
        .C0(\us11/n75 ), .Y(\us11/n72 ) );
  AOI21X1 \us11/U100  ( .A0(\us11/n68 ), .A1(\us11/n69 ), .B0(\us11/n6 ), .Y(
        \us11/n63 ) );
  INVX1 \us11/U99  ( .A(\us11/n67 ), .Y(\us11/n66 ) );
  OAI221XL \us11/U98  ( .A0(\us11/n63 ), .A1(\us11/n64 ), .B0(\us11/n65 ), 
        .B1(\us11/n27 ), .C0(\us11/n66 ), .Y(\us11/n56 ) );
  AOI2BB2X1 \us11/U97  ( .B0(\us11/n61 ), .B1(\us11/n24 ), .A0N(\us11/n62 ), 
        .A1N(\us11/n20 ), .Y(\us11/n60 ) );
  OAI221XL \us11/U96  ( .A0(\us11/n58 ), .A1(\us11/n18 ), .B0(\us11/n59 ), 
        .B1(\us11/n27 ), .C0(\us11/n60 ), .Y(\us11/n57 ) );
  AOI22X1 \us11/U95  ( .A0(\us11/n55 ), .A1(\us11/n56 ), .B0(\us11/n16 ), .B1(
        \us11/n57 ), .Y(\us11/n54 ) );
  OAI221XL \us11/U94  ( .A0(\us11/n51 ), .A1(\us11/n52 ), .B0(\us11/n53 ), 
        .B1(\us11/n10 ), .C0(\us11/n54 ), .Y(\us11/n7 ) );
  INVX1 \us11/U93  ( .A(\us11/n50 ), .Y(\us11/n49 ) );
  OAI221XL \us11/U92  ( .A0(\us11/n47 ), .A1(\us11/n18 ), .B0(\us11/n27 ), 
        .B1(\us11/n48 ), .C0(\us11/n49 ), .Y(\us11/n46 ) );
  NOR2X1 \us11/U91  ( .A(\us11/n41 ), .B(\us11/n42 ), .Y(\us11/n38 ) );
  INVX1 \us11/U90  ( .A(\us11/n40 ), .Y(\us11/n39 ) );
  INVX1 \us11/U89  ( .A(\us11/n32 ), .Y(\us11/n26 ) );
  AOI21X1 \us11/U88  ( .A0(\us11/n5 ), .A1(\us11/n30 ), .B0(\us11/n31 ), .Y(
        \us11/n29 ) );
  OAI221XL \us11/U87  ( .A0(\us11/n26 ), .A1(\us11/n27 ), .B0(\us11/n28 ), 
        .B1(\us11/n20 ), .C0(\us11/n29 ), .Y(\us11/n15 ) );
  OAI221XL \us11/U86  ( .A0(\us11/n18 ), .A1(\us11/n19 ), .B0(\us11/n20 ), 
        .B1(\us11/n21 ), .C0(\us11/n22 ), .Y(\us11/n17 ) );
  AOI22X1 \us11/U85  ( .A0(\us11/n14 ), .A1(\us11/n15 ), .B0(\us11/n16 ), .B1(
        \us11/n17 ), .Y(\us11/n13 ) );
  OAI221XL \us11/U84  ( .A0(\us11/n9 ), .A1(\us11/n10 ), .B0(\us11/n11 ), .B1(
        \us11/n12 ), .C0(\us11/n13 ), .Y(\us11/n8 ) );
  MX2X1 \us11/U83  ( .A(\us11/n7 ), .B(\us11/n8 ), .S0(sa11[6]), .Y(sa10_sr[7]) );
  NOR2X4 \us11/U82  ( .A(\us11/n129 ), .B(sa11[2]), .Y(\us11/n43 ) );
  CLKINVX3 \us11/U81  ( .A(\us11/n14 ), .Y(\us11/n52 ) );
  OAI22XL \us11/U80  ( .A0(\us11/n201 ), .A1(\us11/n52 ), .B0(\us11/n202 ), 
        .B1(\us11/n114 ), .Y(\us11/n193 ) );
  CLKINVX3 \us11/U79  ( .A(sa11[5]), .Y(\us11/n252 ) );
  NOR2X2 \us11/U78  ( .A(\us11/n252 ), .B(\us11/n234 ), .Y(\us11/n55 ) );
  CLKINVX3 \us11/U77  ( .A(sa11[7]), .Y(\us11/n129 ) );
  NOR2X4 \us11/U76  ( .A(\us11/n129 ), .B(\us11/n69 ), .Y(\us11/n24 ) );
  AOI22XL \us11/U75  ( .A0(\us11/n70 ), .A1(\us11/n24 ), .B0(\us11/n96 ), .B1(
        \us11/n129 ), .Y(\us11/n241 ) );
  NOR2X2 \us11/U74  ( .A(\us11/n252 ), .B(sa11[0]), .Y(\us11/n89 ) );
  CLKINVX3 \us11/U73  ( .A(sa11[0]), .Y(\us11/n234 ) );
  NOR2X4 \us11/U72  ( .A(\us11/n69 ), .B(sa11[7]), .Y(\us11/n33 ) );
  INVX12 \us11/U71  ( .A(\us11/n33 ), .Y(\us11/n27 ) );
  CLKINVX3 \us11/U70  ( .A(\us11/n1 ), .Y(\us11/n6 ) );
  CLKINVX3 \us11/U69  ( .A(\us11/n1 ), .Y(\us11/n5 ) );
  INVXL \us11/U68  ( .A(\us11/n24 ), .Y(\us11/n36 ) );
  INVX4 \us11/U67  ( .A(\us11/n3 ), .Y(\us11/n4 ) );
  INVXL \us11/U66  ( .A(\us11/n36 ), .Y(\us11/n3 ) );
  INVX4 \us11/U65  ( .A(sa11[1]), .Y(\us11/n226 ) );
  INVX4 \us11/U64  ( .A(\us11/n43 ), .Y(\us11/n20 ) );
  AOI221X4 \us11/U63  ( .A0(\us11/n24 ), .A1(\us11/n82 ), .B0(\us11/n43 ), 
        .B1(\us11/n295 ), .C0(\us11/n173 ), .Y(\us11/n346 ) );
  AOI221X4 \us11/U62  ( .A0(\us11/n5 ), .A1(\us11/n96 ), .B0(\us11/n43 ), .B1(
        \us11/n239 ), .C0(\us11/n340 ), .Y(\us11/n336 ) );
  AOI222X4 \us11/U61  ( .A0(\us11/n59 ), .A1(\us11/n43 ), .B0(\us11/n6 ), .B1(
        \us11/n221 ), .C0(\us11/n222 ), .C1(\us11/n187 ), .Y(\us11/n218 ) );
  AOI222X4 \us11/U60  ( .A0(\us11/n123 ), .A1(\us11/n43 ), .B0(sa11[2]), .B1(
        \us11/n203 ), .C0(\us11/n6 ), .C1(\us11/n71 ), .Y(\us11/n202 ) );
  AOI221X4 \us11/U59  ( .A0(\us11/n314 ), .A1(\us11/n43 ), .B0(\us11/n160 ), 
        .B1(\us11/n24 ), .C0(\us11/n315 ), .Y(\us11/n307 ) );
  AOI221X4 \us11/U58  ( .A0(\us11/n43 ), .A1(\us11/n208 ), .B0(\us11/n76 ), 
        .B1(\us11/n24 ), .C0(\us11/n209 ), .Y(\us11/n207 ) );
  AOI221X4 \us11/U57  ( .A0(\us11/n43 ), .A1(\us11/n205 ), .B0(\us11/n32 ), 
        .B1(\us11/n6 ), .C0(\us11/n206 ), .Y(\us11/n201 ) );
  AOI221X4 \us11/U56  ( .A0(\us11/n43 ), .A1(\us11/n44 ), .B0(\us11/n45 ), 
        .B1(\us11/n24 ), .C0(\us11/n46 ), .Y(\us11/n9 ) );
  AOI22XL \us11/U55  ( .A0(\us11/n217 ), .A1(\us11/n43 ), .B0(\us11/n33 ), 
        .B1(\us11/n47 ), .Y(\us11/n216 ) );
  AOI22XL \us11/U54  ( .A0(\us11/n98 ), .A1(\us11/n43 ), .B0(\us11/n6 ), .B1(
        \us11/n99 ), .Y(\us11/n97 ) );
  AOI22XL \us11/U53  ( .A0(\us11/n82 ), .A1(\us11/n43 ), .B0(\us11/n83 ), .B1(
        \us11/n24 ), .Y(\us11/n81 ) );
  AOI2BB2XL \us11/U52  ( .B0(\us11/n43 ), .B1(\us11/n94 ), .A0N(\us11/n120 ), 
        .A1N(\us11/n4 ), .Y(\us11/n119 ) );
  AOI222X4 \us11/U51  ( .A0(\us11/n125 ), .A1(\us11/n33 ), .B0(\us11/n145 ), 
        .B1(\us11/n40 ), .C0(\us11/n43 ), .C1(\us11/n184 ), .Y(\us11/n183 ) );
  AOI22XL \us11/U50  ( .A0(\us11/n43 ), .A1(\us11/n303 ), .B0(\us11/n24 ), 
        .B1(\us11/n96 ), .Y(\us11/n358 ) );
  AOI22XL \us11/U49  ( .A0(\us11/n43 ), .A1(\us11/n100 ), .B0(\us11/n24 ), 
        .B1(\us11/n125 ), .Y(\us11/n124 ) );
  AOI21XL \us11/U48  ( .A0(\us11/n159 ), .A1(\us11/n43 ), .B0(\us11/n40 ), .Y(
        \us11/n262 ) );
  AOI22XL \us11/U47  ( .A0(\us11/n40 ), .A1(\us11/n94 ), .B0(\us11/n43 ), .B1(
        \us11/n187 ), .Y(\us11/n244 ) );
  AOI22XL \us11/U46  ( .A0(\us11/n184 ), .A1(\us11/n5 ), .B0(\us11/n198 ), 
        .B1(\us11/n43 ), .Y(\us11/n197 ) );
  NOR2XL \us11/U45  ( .A(\us11/n33 ), .B(\us11/n2 ), .Y(\us11/n302 ) );
  MXI2XL \us11/U44  ( .A(\us11/n2 ), .B(\us11/n6 ), .S0(\us11/n28 ), .Y(
        \us11/n311 ) );
  INVXL \us11/U43  ( .A(\us11/n20 ), .Y(\us11/n2 ) );
  INVX4 \us11/U42  ( .A(\us11/n6 ), .Y(\us11/n18 ) );
  AOI21XL \us11/U41  ( .A0(\us11/n18 ), .A1(\us11/n162 ), .B0(\us11/n25 ), .Y(
        \us11/n161 ) );
  INVX4 \us11/U40  ( .A(sa11[2]), .Y(\us11/n69 ) );
  NOR2X4 \us11/U39  ( .A(\us11/n226 ), .B(\us11/n4 ), .Y(\us11/n40 ) );
  CLKINVX3 \us11/U38  ( .A(sa11[3]), .Y(\us11/n136 ) );
  NOR2X2 \us11/U37  ( .A(\us11/n136 ), .B(sa11[4]), .Y(\us11/n145 ) );
  CLKINVX3 \us11/U36  ( .A(sa11[4]), .Y(\us11/n58 ) );
  NOR2X2 \us11/U35  ( .A(\us11/n58 ), .B(sa11[3]), .Y(\us11/n159 ) );
  NOR2X2 \us11/U34  ( .A(\us11/n136 ), .B(\us11/n58 ), .Y(\us11/n259 ) );
  NOR2X2 \us11/U33  ( .A(sa11[4]), .B(sa11[3]), .Y(\us11/n278 ) );
  NOR2X2 \us11/U32  ( .A(\us11/n259 ), .B(\us11/n278 ), .Y(\us11/n47 ) );
  CLKINVX3 \us11/U31  ( .A(\us11/n259 ), .Y(\us11/n44 ) );
  NOR2X2 \us11/U30  ( .A(\us11/n44 ), .B(sa11[1]), .Y(\us11/n137 ) );
  AOI21XL \us11/U29  ( .A0(\us11/n44 ), .A1(\us11/n111 ), .B0(\us11/n4 ), .Y(
        \us11/n177 ) );
  AOI22XL \us11/U28  ( .A0(\us11/n23 ), .A1(\us11/n24 ), .B0(\us11/n25 ), .B1(
        sa11[2]), .Y(\us11/n22 ) );
  AOI22XL \us11/U27  ( .A0(\us11/n33 ), .A1(sa11[3]), .B0(\us11/n24 ), .B1(
        \us11/n58 ), .Y(\us11/n277 ) );
  NAND2XL \us11/U26  ( .A(\us11/n198 ), .B(\us11/n24 ), .Y(\us11/n132 ) );
  OAI2BB2XL \us11/U25  ( .B0(\us11/n20 ), .B1(\us11/n111 ), .A0N(\us11/n125 ), 
        .A1N(\us11/n24 ), .Y(\us11/n220 ) );
  NAND2XL \us11/U24  ( .A(\us11/n111 ), .B(\us11/n101 ), .Y(\us11/n21 ) );
  NAND2XL \us11/U23  ( .A(\us11/n111 ), .B(\us11/n300 ), .Y(\us11/n187 ) );
  NAND2XL \us11/U22  ( .A(\us11/n111 ), .B(\us11/n121 ), .Y(\us11/n303 ) );
  AOI221XL \us11/U21  ( .A0(\us11/n43 ), .A1(\us11/n151 ), .B0(\us11/n25 ), 
        .B1(\us11/n69 ), .C0(\us11/n275 ), .Y(\us11/n274 ) );
  NOR2BXL \us11/U20  ( .AN(\us11/n101 ), .B(\us11/n25 ), .Y(\us11/n172 ) );
  NAND2X2 \us11/U19  ( .A(\us11/n58 ), .B(\us11/n226 ), .Y(\us11/n34 ) );
  OAI222X1 \us11/U18  ( .A0(\us11/n27 ), .A1(\us11/n34 ), .B0(\us11/n69 ), 
        .B1(\us11/n205 ), .C0(\us11/n20 ), .C1(\us11/n79 ), .Y(\us11/n260 ) );
  OAI222X1 \us11/U17  ( .A0(\us11/n20 ), .A1(\us11/n99 ), .B0(\us11/n27 ), 
        .B1(\us11/n101 ), .C0(\us11/n184 ), .C1(\us11/n4 ), .Y(\us11/n250 ) );
  OAI222X1 \us11/U16  ( .A0(\us11/n4 ), .A1(\us11/n37 ), .B0(\us11/n38 ), .B1(
        \us11/n20 ), .C0(sa11[4]), .C1(\us11/n39 ), .Y(\us11/n35 ) );
  AOI221X1 \us11/U15  ( .A0(\us11/n5 ), .A1(\us11/n19 ), .B0(\us11/n33 ), .B1(
        \us11/n34 ), .C0(\us11/n35 ), .Y(\us11/n11 ) );
  OR2X2 \us11/U14  ( .A(sa11[2]), .B(sa11[7]), .Y(\us11/n1 ) );
  AOI221XL \us11/U13  ( .A0(\us11/n70 ), .A1(\us11/n43 ), .B0(\us11/n24 ), 
        .B1(\us11/n71 ), .C0(\us11/n72 ), .Y(\us11/n53 ) );
  AOI221XL \us11/U12  ( .A0(\us11/n59 ), .A1(\us11/n33 ), .B0(\us11/n43 ), 
        .B1(\us11/n126 ), .C0(\us11/n127 ), .Y(\us11/n113 ) );
  AOI222XL \us11/U11  ( .A0(\us11/n185 ), .A1(\us11/n43 ), .B0(\us11/n186 ), 
        .B1(\us11/n187 ), .C0(\us11/n6 ), .C1(\us11/n188 ), .Y(\us11/n164 ) );
  AOI221X1 \us11/U10  ( .A0(\us11/n313 ), .A1(\us11/n5 ), .B0(\us11/n23 ), 
        .B1(\us11/n2 ), .C0(\us11/n328 ), .Y(\us11/n320 ) );
  AOI221X1 \us11/U9  ( .A0(\us11/n40 ), .A1(\us11/n136 ), .B0(\us11/n33 ), 
        .B1(\us11/n178 ), .C0(\us11/n338 ), .Y(\us11/n337 ) );
  AOI222XL \us11/U8  ( .A0(\us11/n278 ), .A1(\us11/n24 ), .B0(\us11/n42 ), 
        .B1(\us11/n33 ), .C0(\us11/n43 ), .C1(\us11/n136 ), .Y(\us11/n351 ) );
  AOI31X1 \us11/U7  ( .A0(sa11[2]), .A1(\us11/n58 ), .A2(sa11[1]), .B0(
        \us11/n40 ), .Y(\us11/n350 ) );
  AOI31X1 \us11/U6  ( .A0(\us11/n44 ), .A1(\us11/n129 ), .A2(\us11/n130 ), 
        .B0(\us11/n131 ), .Y(\us11/n128 ) );
  AOI221X1 \us11/U5  ( .A0(\us11/n40 ), .A1(\us11/n136 ), .B0(\us11/n33 ), 
        .B1(\us11/n47 ), .C0(\us11/n156 ), .Y(\us11/n141 ) );
  OAI32X1 \us11/U4  ( .A0(\us11/n18 ), .A1(sa11[1]), .A2(\us11/n159 ), .B0(
        sa11[4]), .B1(\us11/n182 ), .Y(\us11/n318 ) );
  OAI32X1 \us11/U3  ( .A0(\us11/n210 ), .A1(\us11/n145 ), .A2(\us11/n18 ), 
        .B0(\us11/n27 ), .B1(\us11/n211 ), .Y(\us11/n209 ) );
  AOI221X1 \us11/U2  ( .A0(\us11/n278 ), .A1(\us11/n40 ), .B0(\us11/n185 ), 
        .B1(\us11/n2 ), .C0(\us11/n279 ), .Y(\us11/n273 ) );
  AOI31XL \us11/U1  ( .A0(\us11/n79 ), .A1(\us11/n44 ), .A2(\us11/n2 ), .B0(
        \us11/n280 ), .Y(\us11/n339 ) );
  NAND2X1 \us12/U366  ( .A(\us12/n47 ), .B(\us12/n226 ), .Y(\us12/n189 ) );
  NOR2X1 \us12/U365  ( .A(\us12/n226 ), .B(sa12[3]), .Y(\us12/n242 ) );
  INVX1 \us12/U364  ( .A(\us12/n242 ), .Y(\us12/n205 ) );
  AND2X1 \us12/U363  ( .A(\us12/n189 ), .B(\us12/n205 ), .Y(\us12/n65 ) );
  NOR2X1 \us12/U362  ( .A(\us12/n226 ), .B(\us12/n47 ), .Y(\us12/n45 ) );
  NOR2X1 \us12/U361  ( .A(\us12/n259 ), .B(\us12/n45 ), .Y(\us12/n73 ) );
  NAND2BX1 \us12/U360  ( .AN(\us12/n73 ), .B(\us12/n6 ), .Y(\us12/n158 ) );
  NOR2X1 \us12/U359  ( .A(\us12/n226 ), .B(\us12/n159 ), .Y(\us12/n95 ) );
  INVX1 \us12/U358  ( .A(\us12/n95 ), .Y(\us12/n111 ) );
  NOR2X1 \us12/U357  ( .A(\us12/n145 ), .B(sa12[1]), .Y(\us12/n42 ) );
  INVX1 \us12/U356  ( .A(\us12/n42 ), .Y(\us12/n121 ) );
  INVX1 \us12/U355  ( .A(\us12/n47 ), .Y(\us12/n96 ) );
  OAI211X1 \us12/U354  ( .A0(\us12/n65 ), .A1(\us12/n27 ), .B0(\us12/n158 ), 
        .C0(\us12/n358 ), .Y(\us12/n355 ) );
  NOR2X1 \us12/U353  ( .A(\us12/n226 ), .B(\us12/n145 ), .Y(\us12/n59 ) );
  NOR2X1 \us12/U352  ( .A(\us12/n96 ), .B(\us12/n59 ), .Y(\us12/n271 ) );
  NOR2X1 \us12/U351  ( .A(\us12/n226 ), .B(\us12/n278 ), .Y(\us12/n217 ) );
  INVX1 \us12/U350  ( .A(\us12/n217 ), .Y(\us12/n150 ) );
  NAND2X1 \us12/U349  ( .A(\us12/n44 ), .B(\us12/n150 ), .Y(\us12/n147 ) );
  NAND2X1 \us12/U348  ( .A(sa12[4]), .B(\us12/n226 ), .Y(\us12/n101 ) );
  INVX1 \us12/U347  ( .A(\us12/n159 ), .Y(\us12/n188 ) );
  NOR2X1 \us12/U346  ( .A(\us12/n188 ), .B(\us12/n226 ), .Y(\us12/n25 ) );
  INVX1 \us12/U345  ( .A(\us12/n172 ), .Y(\us12/n107 ) );
  AOI22X1 \us12/U344  ( .A0(\us12/n33 ), .A1(\us12/n147 ), .B0(\us12/n24 ), 
        .B1(\us12/n107 ), .Y(\us12/n357 ) );
  OAI221XL \us12/U343  ( .A0(\us12/n18 ), .A1(\us12/n121 ), .B0(\us12/n271 ), 
        .B1(\us12/n20 ), .C0(\us12/n357 ), .Y(\us12/n356 ) );
  MXI2X1 \us12/U342  ( .A(\us12/n355 ), .B(\us12/n356 ), .S0(\us12/n252 ), .Y(
        \us12/n331 ) );
  INVX1 \us12/U341  ( .A(\us12/n59 ), .Y(\us12/n79 ) );
  AND2X1 \us12/U340  ( .A(\us12/n101 ), .B(\us12/n79 ), .Y(\us12/n325 ) );
  XNOR2X1 \us12/U339  ( .A(sa12[5]), .B(\us12/n226 ), .Y(\us12/n352 ) );
  NOR2X1 \us12/U338  ( .A(\us12/n226 ), .B(\us12/n136 ), .Y(\us12/n281 ) );
  INVX1 \us12/U337  ( .A(\us12/n281 ), .Y(\us12/n19 ) );
  NAND2X1 \us12/U336  ( .A(\us12/n145 ), .B(\us12/n226 ), .Y(\us12/n223 ) );
  AOI21X1 \us12/U335  ( .A0(\us12/n19 ), .A1(\us12/n223 ), .B0(\us12/n27 ), 
        .Y(\us12/n354 ) );
  AOI31X1 \us12/U334  ( .A0(\us12/n6 ), .A1(\us12/n352 ), .A2(\us12/n259 ), 
        .B0(\us12/n354 ), .Y(\us12/n353 ) );
  OAI221XL \us12/U333  ( .A0(\us12/n20 ), .A1(\us12/n34 ), .B0(\us12/n325 ), 
        .B1(\us12/n4 ), .C0(\us12/n353 ), .Y(\us12/n347 ) );
  INVX1 \us12/U332  ( .A(\us12/n352 ), .Y(\us12/n349 ) );
  NAND2X1 \us12/U331  ( .A(\us12/n278 ), .B(\us12/n6 ), .Y(\us12/n74 ) );
  OAI211X1 \us12/U330  ( .A0(\us12/n349 ), .A1(\us12/n74 ), .B0(\us12/n350 ), 
        .C0(\us12/n351 ), .Y(\us12/n348 ) );
  MXI2X1 \us12/U329  ( .A(\us12/n347 ), .B(\us12/n348 ), .S0(\us12/n252 ), .Y(
        \us12/n332 ) );
  NOR2X1 \us12/U328  ( .A(\us12/n44 ), .B(\us12/n226 ), .Y(\us12/n157 ) );
  INVX1 \us12/U327  ( .A(\us12/n157 ), .Y(\us12/n240 ) );
  NAND2X1 \us12/U326  ( .A(\us12/n240 ), .B(\us12/n189 ), .Y(\us12/n68 ) );
  NOR2X1 \us12/U325  ( .A(\us12/n20 ), .B(\us12/n159 ), .Y(\us12/n225 ) );
  NOR2X1 \us12/U324  ( .A(\us12/n225 ), .B(\us12/n40 ), .Y(\us12/n345 ) );
  INVX1 \us12/U323  ( .A(\us12/n278 ), .Y(\us12/n94 ) );
  NAND2X1 \us12/U322  ( .A(\us12/n94 ), .B(\us12/n226 ), .Y(\us12/n199 ) );
  NAND2X1 \us12/U321  ( .A(\us12/n199 ), .B(\us12/n205 ), .Y(\us12/n82 ) );
  NAND2X1 \us12/U320  ( .A(\us12/n19 ), .B(\us12/n199 ), .Y(\us12/n295 ) );
  NOR2X1 \us12/U319  ( .A(\us12/n226 ), .B(\us12/n259 ), .Y(\us12/n210 ) );
  NOR2X1 \us12/U318  ( .A(\us12/n27 ), .B(\us12/n210 ), .Y(\us12/n173 ) );
  MXI2X1 \us12/U317  ( .A(\us12/n345 ), .B(\us12/n346 ), .S0(\us12/n252 ), .Y(
        \us12/n342 ) );
  NOR2X1 \us12/U316  ( .A(sa12[1]), .B(sa12[3]), .Y(\us12/n163 ) );
  INVX1 \us12/U315  ( .A(\us12/n163 ), .Y(\us12/n37 ) );
  INVX1 \us12/U314  ( .A(\us12/n173 ), .Y(\us12/n344 ) );
  AOI21X1 \us12/U313  ( .A0(\us12/n240 ), .A1(\us12/n37 ), .B0(\us12/n344 ), 
        .Y(\us12/n343 ) );
  AOI211X1 \us12/U312  ( .A0(\us12/n5 ), .A1(\us12/n68 ), .B0(\us12/n342 ), 
        .C0(\us12/n343 ), .Y(\us12/n333 ) );
  NOR2X1 \us12/U311  ( .A(\us12/n18 ), .B(\us12/n226 ), .Y(\us12/n258 ) );
  NAND2X1 \us12/U310  ( .A(\us12/n278 ), .B(sa12[1]), .Y(\us12/n204 ) );
  NOR2X1 \us12/U309  ( .A(\us12/n188 ), .B(sa12[1]), .Y(\us12/n179 ) );
  INVX1 \us12/U308  ( .A(\us12/n179 ), .Y(\us12/n330 ) );
  NAND2X1 \us12/U307  ( .A(\us12/n204 ), .B(\us12/n330 ), .Y(\us12/n239 ) );
  NOR2X1 \us12/U306  ( .A(\us12/n136 ), .B(sa12[1]), .Y(\us12/n299 ) );
  NOR2X1 \us12/U305  ( .A(\us12/n299 ), .B(\us12/n210 ), .Y(\us12/n341 ) );
  OAI32X1 \us12/U304  ( .A0(\us12/n27 ), .A1(\us12/n278 ), .A2(\us12/n95 ), 
        .B0(\us12/n341 ), .B1(\us12/n4 ), .Y(\us12/n340 ) );
  INVX1 \us12/U303  ( .A(\us12/n45 ), .Y(\us12/n126 ) );
  NAND2X1 \us12/U302  ( .A(\us12/n126 ), .B(\us12/n101 ), .Y(\us12/n178 ) );
  NOR2X1 \us12/U301  ( .A(\us12/n18 ), .B(\us12/n136 ), .Y(\us12/n280 ) );
  OAI21XL \us12/U300  ( .A0(\us12/n4 ), .A1(\us12/n121 ), .B0(\us12/n339 ), 
        .Y(\us12/n338 ) );
  MXI2X1 \us12/U299  ( .A(\us12/n336 ), .B(\us12/n337 ), .S0(\us12/n252 ), .Y(
        \us12/n335 ) );
  NOR2X1 \us12/U298  ( .A(\us12/n258 ), .B(\us12/n335 ), .Y(\us12/n334 ) );
  MX4X1 \us12/U297  ( .A(\us12/n331 ), .B(\us12/n332 ), .C(\us12/n333 ), .D(
        \us12/n334 ), .S0(sa12[6]), .S1(\us12/n234 ), .Y(sa11_sr[0]) );
  INVX1 \us12/U296  ( .A(\us12/n299 ), .Y(\us12/n80 ) );
  NOR2X1 \us12/U295  ( .A(\us12/n111 ), .B(\us12/n18 ), .Y(\us12/n269 ) );
  INVX1 \us12/U294  ( .A(\us12/n269 ), .Y(\us12/n75 ) );
  OAI221XL \us12/U293  ( .A0(\us12/n18 ), .A1(\us12/n330 ), .B0(\us12/n20 ), 
        .B1(\us12/n80 ), .C0(\us12/n75 ), .Y(\us12/n329 ) );
  AOI221X1 \us12/U292  ( .A0(\us12/n325 ), .A1(\us12/n33 ), .B0(\us12/n24 ), 
        .B1(\us12/n303 ), .C0(\us12/n329 ), .Y(\us12/n319 ) );
  NOR2X1 \us12/U291  ( .A(\us12/n234 ), .B(sa12[5]), .Y(\us12/n14 ) );
  NOR2X1 \us12/U290  ( .A(\us12/n25 ), .B(\us12/n299 ), .Y(\us12/n313 ) );
  NAND2X1 \us12/U289  ( .A(\us12/n44 ), .B(\us12/n226 ), .Y(\us12/n300 ) );
  AND2X1 \us12/U288  ( .A(\us12/n300 ), .B(\us12/n240 ), .Y(\us12/n23 ) );
  OAI32X1 \us12/U287  ( .A0(\us12/n4 ), .A1(\us12/n145 ), .A2(\us12/n210 ), 
        .B0(\us12/n137 ), .B1(\us12/n27 ), .Y(\us12/n328 ) );
  NOR2X1 \us12/U286  ( .A(sa12[0]), .B(sa12[5]), .Y(\us12/n16 ) );
  INVX1 \us12/U285  ( .A(\us12/n16 ), .Y(\us12/n114 ) );
  INVX1 \us12/U284  ( .A(\us12/n145 ), .Y(\us12/n149 ) );
  NOR2X1 \us12/U283  ( .A(\us12/n47 ), .B(sa12[1]), .Y(\us12/n98 ) );
  INVX1 \us12/U282  ( .A(\us12/n98 ), .Y(\us12/n284 ) );
  OAI21XL \us12/U281  ( .A0(\us12/n69 ), .A1(\us12/n284 ), .B0(\us12/n27 ), 
        .Y(\us12/n327 ) );
  AOI31X1 \us12/U280  ( .A0(\us12/n111 ), .A1(\us12/n149 ), .A2(\us12/n327 ), 
        .B0(\us12/n225 ), .Y(\us12/n326 ) );
  OAI21XL \us12/U279  ( .A0(\us12/n325 ), .A1(\us12/n18 ), .B0(\us12/n326 ), 
        .Y(\us12/n322 ) );
  NAND2X1 \us12/U278  ( .A(\us12/n19 ), .B(\us12/n189 ), .Y(\us12/n71 ) );
  NOR2X1 \us12/U277  ( .A(\us12/n71 ), .B(\us12/n18 ), .Y(\us12/n135 ) );
  AOI21X1 \us12/U276  ( .A0(\us12/n40 ), .A1(sa12[4]), .B0(\us12/n135 ), .Y(
        \us12/n324 ) );
  OAI221XL \us12/U275  ( .A0(\us12/n47 ), .A1(\us12/n27 ), .B0(\us12/n65 ), 
        .B1(\us12/n20 ), .C0(\us12/n324 ), .Y(\us12/n323 ) );
  AOI22X1 \us12/U274  ( .A0(\us12/n55 ), .A1(\us12/n322 ), .B0(\us12/n89 ), 
        .B1(\us12/n323 ), .Y(\us12/n321 ) );
  OAI221XL \us12/U273  ( .A0(\us12/n319 ), .A1(\us12/n52 ), .B0(\us12/n320 ), 
        .B1(\us12/n114 ), .C0(\us12/n321 ), .Y(\us12/n304 ) );
  NOR2X1 \us12/U272  ( .A(\us12/n226 ), .B(\us12/n58 ), .Y(\us12/n290 ) );
  INVX1 \us12/U271  ( .A(\us12/n290 ), .Y(\us12/n200 ) );
  NAND2X1 \us12/U270  ( .A(\us12/n34 ), .B(\us12/n200 ), .Y(\us12/n120 ) );
  INVX1 \us12/U269  ( .A(\us12/n210 ), .Y(\us12/n100 ) );
  OAI221XL \us12/U268  ( .A0(\us12/n20 ), .A1(\us12/n100 ), .B0(sa12[3]), .B1(
        \us12/n4 ), .C0(\us12/n262 ), .Y(\us12/n317 ) );
  INVX1 \us12/U267  ( .A(\us12/n258 ), .Y(\us12/n182 ) );
  AOI211X1 \us12/U266  ( .A0(\us12/n33 ), .A1(\us12/n120 ), .B0(\us12/n317 ), 
        .C0(\us12/n318 ), .Y(\us12/n306 ) );
  NAND2X1 \us12/U265  ( .A(\us12/n100 ), .B(\us12/n199 ), .Y(\us12/n151 ) );
  INVX1 \us12/U264  ( .A(\us12/n151 ), .Y(\us12/n314 ) );
  NOR2X1 \us12/U263  ( .A(\us12/n45 ), .B(\us12/n163 ), .Y(\us12/n160 ) );
  INVX1 \us12/U262  ( .A(\us12/n295 ), .Y(\us12/n92 ) );
  AOI21X1 \us12/U261  ( .A0(sa12[1]), .A1(\us12/n58 ), .B0(\us12/n98 ), .Y(
        \us12/n316 ) );
  OAI22X1 \us12/U260  ( .A0(\us12/n92 ), .A1(\us12/n18 ), .B0(\us12/n316 ), 
        .B1(\us12/n27 ), .Y(\us12/n315 ) );
  NOR2X1 \us12/U259  ( .A(\us12/n149 ), .B(\us12/n226 ), .Y(\us12/n41 ) );
  INVX1 \us12/U258  ( .A(\us12/n41 ), .Y(\us12/n105 ) );
  NAND2X1 \us12/U257  ( .A(\us12/n284 ), .B(\us12/n105 ), .Y(\us12/n227 ) );
  AOI21X1 \us12/U256  ( .A0(\us12/n313 ), .A1(\us12/n33 ), .B0(\us12/n269 ), 
        .Y(\us12/n312 ) );
  OAI221XL \us12/U255  ( .A0(\us12/n149 ), .A1(\us12/n20 ), .B0(\us12/n4 ), 
        .B1(\us12/n227 ), .C0(\us12/n312 ), .Y(\us12/n309 ) );
  AOI21X1 \us12/U254  ( .A0(\us12/n226 ), .A1(\us12/n188 ), .B0(\us12/n242 ), 
        .Y(\us12/n185 ) );
  INVX1 \us12/U253  ( .A(\us12/n185 ), .Y(\us12/n48 ) );
  AND2X1 \us12/U252  ( .A(\us12/n223 ), .B(\us12/n240 ), .Y(\us12/n28 ) );
  OAI221XL \us12/U251  ( .A0(\us12/n27 ), .A1(\us12/n44 ), .B0(\us12/n4 ), 
        .B1(\us12/n48 ), .C0(\us12/n311 ), .Y(\us12/n310 ) );
  AOI22X1 \us12/U250  ( .A0(\us12/n89 ), .A1(\us12/n309 ), .B0(\us12/n55 ), 
        .B1(\us12/n310 ), .Y(\us12/n308 ) );
  OAI221XL \us12/U249  ( .A0(\us12/n306 ), .A1(\us12/n52 ), .B0(\us12/n307 ), 
        .B1(\us12/n114 ), .C0(\us12/n308 ), .Y(\us12/n305 ) );
  MX2X1 \us12/U248  ( .A(\us12/n304 ), .B(\us12/n305 ), .S0(sa12[6]), .Y(
        sa11_sr[1]) );
  INVX1 \us12/U247  ( .A(\us12/n187 ), .Y(\us12/n61 ) );
  MXI2X1 \us12/U246  ( .A(\us12/n303 ), .B(\us12/n61 ), .S0(\us12/n69 ), .Y(
        \us12/n301 ) );
  MXI2X1 \us12/U245  ( .A(\us12/n301 ), .B(\us12/n147 ), .S0(\us12/n302 ), .Y(
        \us12/n285 ) );
  NAND2X1 \us12/U244  ( .A(\us12/n200 ), .B(\us12/n300 ), .Y(\us12/n99 ) );
  INVX1 \us12/U243  ( .A(\us12/n99 ), .Y(\us12/n296 ) );
  NOR2X1 \us12/U242  ( .A(\us12/n299 ), .B(\us12/n242 ), .Y(\us12/n298 ) );
  NAND2X1 \us12/U241  ( .A(sa12[1]), .B(\us12/n47 ), .Y(\us12/n122 ) );
  NOR2X1 \us12/U240  ( .A(\us12/n159 ), .B(\us12/n217 ), .Y(\us12/n198 ) );
  OAI221XL \us12/U239  ( .A0(\us12/n298 ), .A1(\us12/n27 ), .B0(\us12/n20 ), 
        .B1(\us12/n122 ), .C0(\us12/n132 ), .Y(\us12/n297 ) );
  AOI221X1 \us12/U238  ( .A0(\us12/n225 ), .A1(\us12/n226 ), .B0(\us12/n296 ), 
        .B1(\us12/n6 ), .C0(\us12/n297 ), .Y(\us12/n291 ) );
  OAI2BB2X1 \us12/U237  ( .B0(\us12/n27 ), .B1(\us12/n295 ), .A0N(\us12/n34 ), 
        .A1N(\us12/n24 ), .Y(\us12/n293 ) );
  AOI21X1 \us12/U236  ( .A0(\us12/n101 ), .A1(\us12/n150 ), .B0(\us12/n20 ), 
        .Y(\us12/n294 ) );
  AOI211X1 \us12/U235  ( .A0(\us12/n5 ), .A1(\us12/n79 ), .B0(\us12/n293 ), 
        .C0(\us12/n294 ), .Y(\us12/n292 ) );
  INVX1 \us12/U234  ( .A(\us12/n89 ), .Y(\us12/n10 ) );
  OAI22X1 \us12/U233  ( .A0(\us12/n291 ), .A1(\us12/n114 ), .B0(\us12/n292 ), 
        .B1(\us12/n10 ), .Y(\us12/n286 ) );
  INVX1 \us12/U232  ( .A(\us12/n225 ), .Y(\us12/n288 ) );
  NAND2X1 \us12/U231  ( .A(\us12/n200 ), .B(\us12/n284 ), .Y(\us12/n102 ) );
  NOR2X1 \us12/U230  ( .A(\us12/n290 ), .B(\us12/n163 ), .Y(\us12/n184 ) );
  AOI22X1 \us12/U229  ( .A0(\us12/n102 ), .A1(\us12/n69 ), .B0(\us12/n184 ), 
        .B1(\us12/n33 ), .Y(\us12/n289 ) );
  AOI31X1 \us12/U228  ( .A0(\us12/n132 ), .A1(\us12/n288 ), .A2(\us12/n289 ), 
        .B0(\us12/n52 ), .Y(\us12/n287 ) );
  AOI211X1 \us12/U227  ( .A0(\us12/n285 ), .A1(\us12/n55 ), .B0(\us12/n286 ), 
        .C0(\us12/n287 ), .Y(\us12/n263 ) );
  NAND2X1 \us12/U226  ( .A(\us12/n284 ), .B(\us12/n122 ), .Y(\us12/n125 ) );
  NOR2X1 \us12/U225  ( .A(\us12/n199 ), .B(\us12/n4 ), .Y(\us12/n50 ) );
  AOI21X1 \us12/U224  ( .A0(\us12/n200 ), .A1(\us12/n223 ), .B0(\us12/n20 ), 
        .Y(\us12/n283 ) );
  AOI211X1 \us12/U223  ( .A0(\us12/n5 ), .A1(\us12/n125 ), .B0(\us12/n50 ), 
        .C0(\us12/n283 ), .Y(\us12/n282 ) );
  OAI221XL \us12/U222  ( .A0(\us12/n281 ), .A1(\us12/n27 ), .B0(\us12/n4 ), 
        .B1(\us12/n111 ), .C0(\us12/n282 ), .Y(\us12/n265 ) );
  INVX1 \us12/U221  ( .A(\us12/n280 ), .Y(\us12/n247 ) );
  NAND2X1 \us12/U220  ( .A(\us12/n41 ), .B(\us12/n33 ), .Y(\us12/n272 ) );
  OAI221XL \us12/U219  ( .A0(sa12[1]), .A1(\us12/n247 ), .B0(\us12/n4 ), .B1(
        \us12/n189 ), .C0(\us12/n272 ), .Y(\us12/n279 ) );
  NAND2X1 \us12/U218  ( .A(sa12[2]), .B(\us12/n149 ), .Y(\us12/n276 ) );
  XNOR2X1 \us12/U217  ( .A(\us12/n129 ), .B(sa12[1]), .Y(\us12/n155 ) );
  MXI2X1 \us12/U216  ( .A(\us12/n276 ), .B(\us12/n277 ), .S0(\us12/n155 ), .Y(
        \us12/n275 ) );
  OAI22X1 \us12/U215  ( .A0(\us12/n273 ), .A1(\us12/n10 ), .B0(\us12/n274 ), 
        .B1(\us12/n52 ), .Y(\us12/n266 ) );
  NOR2X1 \us12/U214  ( .A(\us12/n20 ), .B(\us12/n226 ), .Y(\us12/n176 ) );
  OAI21XL \us12/U213  ( .A0(\us12/n4 ), .A1(\us12/n271 ), .B0(\us12/n272 ), 
        .Y(\us12/n270 ) );
  OAI31X1 \us12/U212  ( .A0(\us12/n176 ), .A1(\us12/n269 ), .A2(\us12/n270 ), 
        .B0(\us12/n16 ), .Y(\us12/n268 ) );
  INVX1 \us12/U211  ( .A(\us12/n268 ), .Y(\us12/n267 ) );
  AOI211X1 \us12/U210  ( .A0(\us12/n55 ), .A1(\us12/n265 ), .B0(\us12/n266 ), 
        .C0(\us12/n267 ), .Y(\us12/n264 ) );
  MXI2X1 \us12/U209  ( .A(\us12/n263 ), .B(\us12/n264 ), .S0(sa12[6]), .Y(
        sa11_sr[2]) );
  NOR2X1 \us12/U208  ( .A(\us12/n94 ), .B(sa12[1]), .Y(\us12/n211 ) );
  INVX1 \us12/U207  ( .A(\us12/n262 ), .Y(\us12/n261 ) );
  AOI211X1 \us12/U206  ( .A0(\us12/n259 ), .A1(\us12/n24 ), .B0(\us12/n260 ), 
        .C0(\us12/n261 ), .Y(\us12/n255 ) );
  OAI22X1 \us12/U205  ( .A0(\us12/n20 ), .A1(\us12/n68 ), .B0(\us12/n27 ), 
        .B1(\us12/n37 ), .Y(\us12/n257 ) );
  NOR3X1 \us12/U204  ( .A(\us12/n257 ), .B(\us12/n258 ), .C(\us12/n50 ), .Y(
        \us12/n256 ) );
  MXI2X1 \us12/U203  ( .A(\us12/n255 ), .B(\us12/n256 ), .S0(\us12/n252 ), .Y(
        \us12/n254 ) );
  AOI221X1 \us12/U202  ( .A0(\us12/n211 ), .A1(\us12/n5 ), .B0(\us12/n40 ), 
        .B1(sa12[4]), .C0(\us12/n254 ), .Y(\us12/n248 ) );
  INVX1 \us12/U201  ( .A(\us12/n211 ), .Y(\us12/n106 ) );
  NAND2X1 \us12/U200  ( .A(\us12/n200 ), .B(\us12/n106 ), .Y(\us12/n83 ) );
  NAND2X1 \us12/U199  ( .A(\us12/n199 ), .B(\us12/n204 ), .Y(\us12/n169 ) );
  AOI2BB2X1 \us12/U198  ( .B0(\us12/n65 ), .B1(\us12/n24 ), .A0N(\us12/n169 ), 
        .A1N(\us12/n20 ), .Y(\us12/n253 ) );
  OAI221XL \us12/U197  ( .A0(\us12/n172 ), .A1(\us12/n18 ), .B0(\us12/n27 ), 
        .B1(\us12/n83 ), .C0(\us12/n253 ), .Y(\us12/n251 ) );
  MXI2X1 \us12/U196  ( .A(\us12/n250 ), .B(\us12/n251 ), .S0(\us12/n252 ), .Y(
        \us12/n249 ) );
  MXI2X1 \us12/U195  ( .A(\us12/n248 ), .B(\us12/n249 ), .S0(\us12/n234 ), .Y(
        \us12/n228 ) );
  OAI21XL \us12/U194  ( .A0(\us12/n58 ), .A1(\us12/n27 ), .B0(\us12/n247 ), 
        .Y(\us12/n245 ) );
  NOR2X1 \us12/U193  ( .A(sa12[7]), .B(\us12/n145 ), .Y(\us12/n246 ) );
  XNOR2X1 \us12/U192  ( .A(\us12/n69 ), .B(sa12[1]), .Y(\us12/n130 ) );
  MXI2X1 \us12/U191  ( .A(\us12/n245 ), .B(\us12/n246 ), .S0(\us12/n130 ), .Y(
        \us12/n243 ) );
  OAI211X1 \us12/U190  ( .A0(\us12/n4 ), .A1(\us12/n149 ), .B0(\us12/n243 ), 
        .C0(\us12/n244 ), .Y(\us12/n230 ) );
  NOR2X1 \us12/U189  ( .A(\us12/n242 ), .B(\us12/n137 ), .Y(\us12/n70 ) );
  OAI221XL \us12/U188  ( .A0(\us12/n159 ), .A1(\us12/n27 ), .B0(\us12/n20 ), 
        .B1(\us12/n34 ), .C0(\us12/n241 ), .Y(\us12/n231 ) );
  NAND2X1 \us12/U187  ( .A(\us12/n101 ), .B(\us12/n240 ), .Y(\us12/n76 ) );
  AOI21X1 \us12/U186  ( .A0(\us12/n122 ), .A1(\us12/n106 ), .B0(\us12/n129 ), 
        .Y(\us12/n237 ) );
  INVX1 \us12/U185  ( .A(\us12/n239 ), .Y(\us12/n238 ) );
  OAI21XL \us12/U184  ( .A0(\us12/n237 ), .A1(\us12/n43 ), .B0(\us12/n238 ), 
        .Y(\us12/n236 ) );
  OAI221XL \us12/U183  ( .A0(\us12/n18 ), .A1(\us12/n76 ), .B0(\us12/n59 ), 
        .B1(\us12/n27 ), .C0(\us12/n236 ), .Y(\us12/n232 ) );
  AOI2BB2X1 \us12/U182  ( .B0(\us12/n24 ), .B1(\us12/n187 ), .A0N(\us12/n227 ), 
        .A1N(\us12/n20 ), .Y(\us12/n235 ) );
  OAI211X1 \us12/U181  ( .A0(\us12/n27 ), .A1(\us12/n122 ), .B0(\us12/n158 ), 
        .C0(\us12/n235 ), .Y(\us12/n233 ) );
  MX4X1 \us12/U180  ( .A(\us12/n230 ), .B(\us12/n231 ), .C(\us12/n232 ), .D(
        \us12/n233 ), .S0(\us12/n234 ), .S1(sa12[5]), .Y(\us12/n229 ) );
  MX2X1 \us12/U179  ( .A(\us12/n228 ), .B(\us12/n229 ), .S0(sa12[6]), .Y(
        sa11_sr[3]) );
  NOR2BX1 \us12/U178  ( .AN(\us12/n204 ), .B(\us12/n137 ), .Y(\us12/n110 ) );
  INVX1 \us12/U177  ( .A(\us12/n110 ), .Y(\us12/n64 ) );
  AOI22X1 \us12/U176  ( .A0(\us12/n225 ), .A1(\us12/n226 ), .B0(\us12/n6 ), 
        .B1(\us12/n227 ), .Y(\us12/n224 ) );
  OAI221XL \us12/U175  ( .A0(\us12/n27 ), .A1(\us12/n64 ), .B0(\us12/n4 ), 
        .B1(\us12/n83 ), .C0(\us12/n224 ), .Y(\us12/n212 ) );
  NAND2X1 \us12/U174  ( .A(\us12/n34 ), .B(\us12/n204 ), .Y(\us12/n221 ) );
  OAI21XL \us12/U173  ( .A0(\us12/n69 ), .A1(\us12/n223 ), .B0(\us12/n27 ), 
        .Y(\us12/n222 ) );
  NOR2X1 \us12/U172  ( .A(\us12/n217 ), .B(\us12/n42 ), .Y(\us12/n208 ) );
  AOI211X1 \us12/U171  ( .A0(\us12/n208 ), .A1(\us12/n5 ), .B0(\us12/n220 ), 
        .C0(\us12/n173 ), .Y(\us12/n219 ) );
  OAI22X1 \us12/U170  ( .A0(\us12/n218 ), .A1(\us12/n10 ), .B0(\us12/n219 ), 
        .B1(\us12/n114 ), .Y(\us12/n213 ) );
  INVX1 \us12/U169  ( .A(\us12/n135 ), .Y(\us12/n215 ) );
  NOR2X1 \us12/U168  ( .A(\us12/n4 ), .B(\us12/n159 ), .Y(\us12/n31 ) );
  INVX1 \us12/U167  ( .A(\us12/n31 ), .Y(\us12/n196 ) );
  AOI31X1 \us12/U166  ( .A0(\us12/n215 ), .A1(\us12/n196 ), .A2(\us12/n216 ), 
        .B0(\us12/n52 ), .Y(\us12/n214 ) );
  AOI211X1 \us12/U165  ( .A0(\us12/n55 ), .A1(\us12/n212 ), .B0(\us12/n213 ), 
        .C0(\us12/n214 ), .Y(\us12/n190 ) );
  INVX1 \us12/U164  ( .A(\us12/n207 ), .Y(\us12/n192 ) );
  NOR2X1 \us12/U163  ( .A(\us12/n25 ), .B(\us12/n98 ), .Y(\us12/n32 ) );
  OAI22X1 \us12/U162  ( .A0(\us12/n28 ), .A1(\us12/n4 ), .B0(\us12/n188 ), 
        .B1(\us12/n27 ), .Y(\us12/n206 ) );
  NAND2X1 \us12/U161  ( .A(\us12/n204 ), .B(\us12/n80 ), .Y(\us12/n118 ) );
  INVX1 \us12/U160  ( .A(\us12/n118 ), .Y(\us12/n123 ) );
  NAND2X1 \us12/U159  ( .A(\us12/n94 ), .B(\us12/n79 ), .Y(\us12/n203 ) );
  OAI2BB1X1 \us12/U158  ( .A0N(\us12/n199 ), .A1N(\us12/n200 ), .B0(\us12/n33 ), .Y(\us12/n195 ) );
  INVX1 \us12/U157  ( .A(\us12/n55 ), .Y(\us12/n12 ) );
  AOI31X1 \us12/U156  ( .A0(\us12/n195 ), .A1(\us12/n196 ), .A2(\us12/n197 ), 
        .B0(\us12/n12 ), .Y(\us12/n194 ) );
  AOI211X1 \us12/U155  ( .A0(\us12/n89 ), .A1(\us12/n192 ), .B0(\us12/n193 ), 
        .C0(\us12/n194 ), .Y(\us12/n191 ) );
  MXI2X1 \us12/U154  ( .A(\us12/n190 ), .B(\us12/n191 ), .S0(sa12[6]), .Y(
        sa11_sr[4]) );
  OAI21XL \us12/U153  ( .A0(\us12/n69 ), .A1(\us12/n189 ), .B0(\us12/n27 ), 
        .Y(\us12/n186 ) );
  INVX1 \us12/U152  ( .A(\us12/n183 ), .Y(\us12/n180 ) );
  NAND2X1 \us12/U151  ( .A(\us12/n74 ), .B(\us12/n182 ), .Y(\us12/n181 ) );
  AOI211X1 \us12/U150  ( .A0(\us12/n179 ), .A1(\us12/n24 ), .B0(\us12/n180 ), 
        .C0(\us12/n181 ), .Y(\us12/n165 ) );
  INVX1 \us12/U149  ( .A(\us12/n178 ), .Y(\us12/n175 ) );
  AOI211X1 \us12/U148  ( .A0(\us12/n175 ), .A1(\us12/n5 ), .B0(\us12/n176 ), 
        .C0(\us12/n177 ), .Y(\us12/n174 ) );
  OAI221XL \us12/U147  ( .A0(\us12/n159 ), .A1(\us12/n27 ), .B0(\us12/n145 ), 
        .B1(\us12/n20 ), .C0(\us12/n174 ), .Y(\us12/n167 ) );
  MXI2X1 \us12/U146  ( .A(\us12/n40 ), .B(\us12/n173 ), .S0(\us12/n96 ), .Y(
        \us12/n170 ) );
  AOI22X1 \us12/U145  ( .A0(\us12/n137 ), .A1(\us12/n24 ), .B0(\us12/n172 ), 
        .B1(\us12/n6 ), .Y(\us12/n171 ) );
  OAI211X1 \us12/U144  ( .A0(\us12/n20 ), .A1(\us12/n169 ), .B0(\us12/n170 ), 
        .C0(\us12/n171 ), .Y(\us12/n168 ) );
  AOI22X1 \us12/U143  ( .A0(\us12/n89 ), .A1(\us12/n167 ), .B0(\us12/n55 ), 
        .B1(\us12/n168 ), .Y(\us12/n166 ) );
  OAI221XL \us12/U142  ( .A0(\us12/n164 ), .A1(\us12/n114 ), .B0(\us12/n165 ), 
        .B1(\us12/n52 ), .C0(\us12/n166 ), .Y(\us12/n138 ) );
  OAI21XL \us12/U141  ( .A0(\us12/n41 ), .A1(\us12/n163 ), .B0(\us12/n69 ), 
        .Y(\us12/n162 ) );
  AOI221X1 \us12/U140  ( .A0(\us12/n159 ), .A1(\us12/n24 ), .B0(\us12/n160 ), 
        .B1(\us12/n33 ), .C0(\us12/n161 ), .Y(\us12/n140 ) );
  OAI21XL \us12/U139  ( .A0(\us12/n157 ), .A1(\us12/n20 ), .B0(\us12/n158 ), 
        .Y(\us12/n156 ) );
  NOR2X1 \us12/U138  ( .A(\us12/n4 ), .B(\us12/n136 ), .Y(\us12/n153 ) );
  NOR2X1 \us12/U137  ( .A(\us12/n145 ), .B(\us12/n69 ), .Y(\us12/n154 ) );
  MXI2X1 \us12/U136  ( .A(\us12/n153 ), .B(\us12/n154 ), .S0(\us12/n155 ), .Y(
        \us12/n152 ) );
  OAI221XL \us12/U135  ( .A0(\us12/n110 ), .A1(\us12/n18 ), .B0(\us12/n20 ), 
        .B1(\us12/n151 ), .C0(\us12/n152 ), .Y(\us12/n143 ) );
  AOI21X1 \us12/U134  ( .A0(\us12/n149 ), .A1(\us12/n150 ), .B0(\us12/n18 ), 
        .Y(\us12/n148 ) );
  AOI2BB1X1 \us12/U133  ( .A0N(\us12/n147 ), .A1N(\us12/n27 ), .B0(\us12/n148 ), .Y(\us12/n146 ) );
  OAI221XL \us12/U132  ( .A0(\us12/n145 ), .A1(\us12/n20 ), .B0(\us12/n4 ), 
        .B1(\us12/n34 ), .C0(\us12/n146 ), .Y(\us12/n144 ) );
  AOI22X1 \us12/U131  ( .A0(\us12/n89 ), .A1(\us12/n143 ), .B0(\us12/n14 ), 
        .B1(\us12/n144 ), .Y(\us12/n142 ) );
  OAI221XL \us12/U130  ( .A0(\us12/n140 ), .A1(\us12/n12 ), .B0(\us12/n141 ), 
        .B1(\us12/n114 ), .C0(\us12/n142 ), .Y(\us12/n139 ) );
  MX2X1 \us12/U129  ( .A(\us12/n138 ), .B(\us12/n139 ), .S0(sa12[6]), .Y(
        sa11_sr[5]) );
  INVX1 \us12/U128  ( .A(\us12/n70 ), .Y(\us12/n133 ) );
  OAI22X1 \us12/U127  ( .A0(\us12/n4 ), .A1(\us12/n136 ), .B0(\us12/n137 ), 
        .B1(\us12/n27 ), .Y(\us12/n134 ) );
  AOI211X1 \us12/U126  ( .A0(\us12/n133 ), .A1(\us12/n69 ), .B0(\us12/n134 ), 
        .C0(\us12/n135 ), .Y(\us12/n112 ) );
  INVX1 \us12/U125  ( .A(\us12/n132 ), .Y(\us12/n131 ) );
  OAI21XL \us12/U124  ( .A0(\us12/n18 ), .A1(\us12/n37 ), .B0(\us12/n128 ), 
        .Y(\us12/n127 ) );
  OAI221XL \us12/U123  ( .A0(\us12/n18 ), .A1(\us12/n105 ), .B0(\us12/n123 ), 
        .B1(\us12/n27 ), .C0(\us12/n124 ), .Y(\us12/n116 ) );
  NAND2X1 \us12/U122  ( .A(\us12/n121 ), .B(\us12/n122 ), .Y(\us12/n30 ) );
  OAI221XL \us12/U121  ( .A0(\us12/n18 ), .A1(\us12/n118 ), .B0(\us12/n27 ), 
        .B1(\us12/n30 ), .C0(\us12/n119 ), .Y(\us12/n117 ) );
  AOI22X1 \us12/U120  ( .A0(\us12/n89 ), .A1(\us12/n116 ), .B0(\us12/n55 ), 
        .B1(\us12/n117 ), .Y(\us12/n115 ) );
  OAI221XL \us12/U119  ( .A0(\us12/n112 ), .A1(\us12/n52 ), .B0(\us12/n113 ), 
        .B1(\us12/n114 ), .C0(\us12/n115 ), .Y(\us12/n84 ) );
  OAI22X1 \us12/U118  ( .A0(\us12/n110 ), .A1(\us12/n4 ), .B0(\us12/n20 ), 
        .B1(\us12/n21 ), .Y(\us12/n108 ) );
  AOI21X1 \us12/U117  ( .A0(sa12[1]), .A1(\us12/n58 ), .B0(\us12/n27 ), .Y(
        \us12/n109 ) );
  AOI211X1 \us12/U116  ( .A0(\us12/n5 ), .A1(\us12/n107 ), .B0(\us12/n108 ), 
        .C0(\us12/n109 ), .Y(\us12/n86 ) );
  OAI22X1 \us12/U115  ( .A0(\us12/n45 ), .A1(\us12/n4 ), .B0(sa12[4]), .B1(
        \us12/n18 ), .Y(\us12/n103 ) );
  AOI21X1 \us12/U114  ( .A0(\us12/n105 ), .A1(\us12/n106 ), .B0(\us12/n20 ), 
        .Y(\us12/n104 ) );
  AOI211X1 \us12/U113  ( .A0(\us12/n33 ), .A1(\us12/n102 ), .B0(\us12/n103 ), 
        .C0(\us12/n104 ), .Y(\us12/n87 ) );
  NAND2X1 \us12/U112  ( .A(\us12/n100 ), .B(\us12/n101 ), .Y(\us12/n62 ) );
  OAI221XL \us12/U111  ( .A0(\us12/n27 ), .A1(\us12/n62 ), .B0(\us12/n4 ), 
        .B1(\us12/n21 ), .C0(\us12/n97 ), .Y(\us12/n90 ) );
  NOR3X1 \us12/U110  ( .A(\us12/n4 ), .B(\us12/n95 ), .C(\us12/n96 ), .Y(
        \us12/n67 ) );
  AOI31X1 \us12/U109  ( .A0(\us12/n79 ), .A1(\us12/n94 ), .A2(\us12/n6 ), .B0(
        \us12/n67 ), .Y(\us12/n93 ) );
  OAI221XL \us12/U108  ( .A0(\us12/n73 ), .A1(\us12/n27 ), .B0(\us12/n92 ), 
        .B1(\us12/n20 ), .C0(\us12/n93 ), .Y(\us12/n91 ) );
  AOI22X1 \us12/U107  ( .A0(\us12/n89 ), .A1(\us12/n90 ), .B0(\us12/n16 ), 
        .B1(\us12/n91 ), .Y(\us12/n88 ) );
  OAI221XL \us12/U106  ( .A0(\us12/n86 ), .A1(\us12/n52 ), .B0(\us12/n87 ), 
        .B1(\us12/n12 ), .C0(\us12/n88 ), .Y(\us12/n85 ) );
  MX2X1 \us12/U105  ( .A(\us12/n84 ), .B(\us12/n85 ), .S0(sa12[6]), .Y(
        sa11_sr[6]) );
  INVX1 \us12/U104  ( .A(\us12/n81 ), .Y(\us12/n77 ) );
  AOI21X1 \us12/U103  ( .A0(\us12/n79 ), .A1(\us12/n80 ), .B0(\us12/n27 ), .Y(
        \us12/n78 ) );
  AOI211X1 \us12/U102  ( .A0(\us12/n5 ), .A1(\us12/n76 ), .B0(\us12/n77 ), 
        .C0(\us12/n78 ), .Y(\us12/n51 ) );
  OAI211X1 \us12/U101  ( .A0(\us12/n73 ), .A1(\us12/n27 ), .B0(\us12/n74 ), 
        .C0(\us12/n75 ), .Y(\us12/n72 ) );
  AOI21X1 \us12/U100  ( .A0(\us12/n68 ), .A1(\us12/n69 ), .B0(\us12/n6 ), .Y(
        \us12/n63 ) );
  INVX1 \us12/U99  ( .A(\us12/n67 ), .Y(\us12/n66 ) );
  OAI221XL \us12/U98  ( .A0(\us12/n63 ), .A1(\us12/n64 ), .B0(\us12/n65 ), 
        .B1(\us12/n27 ), .C0(\us12/n66 ), .Y(\us12/n56 ) );
  AOI2BB2X1 \us12/U97  ( .B0(\us12/n61 ), .B1(\us12/n24 ), .A0N(\us12/n62 ), 
        .A1N(\us12/n20 ), .Y(\us12/n60 ) );
  OAI221XL \us12/U96  ( .A0(\us12/n58 ), .A1(\us12/n18 ), .B0(\us12/n59 ), 
        .B1(\us12/n27 ), .C0(\us12/n60 ), .Y(\us12/n57 ) );
  AOI22X1 \us12/U95  ( .A0(\us12/n55 ), .A1(\us12/n56 ), .B0(\us12/n16 ), .B1(
        \us12/n57 ), .Y(\us12/n54 ) );
  OAI221XL \us12/U94  ( .A0(\us12/n51 ), .A1(\us12/n52 ), .B0(\us12/n53 ), 
        .B1(\us12/n10 ), .C0(\us12/n54 ), .Y(\us12/n7 ) );
  INVX1 \us12/U93  ( .A(\us12/n50 ), .Y(\us12/n49 ) );
  OAI221XL \us12/U92  ( .A0(\us12/n47 ), .A1(\us12/n18 ), .B0(\us12/n27 ), 
        .B1(\us12/n48 ), .C0(\us12/n49 ), .Y(\us12/n46 ) );
  NOR2X1 \us12/U91  ( .A(\us12/n41 ), .B(\us12/n42 ), .Y(\us12/n38 ) );
  INVX1 \us12/U90  ( .A(\us12/n40 ), .Y(\us12/n39 ) );
  INVX1 \us12/U89  ( .A(\us12/n32 ), .Y(\us12/n26 ) );
  AOI21X1 \us12/U88  ( .A0(\us12/n5 ), .A1(\us12/n30 ), .B0(\us12/n31 ), .Y(
        \us12/n29 ) );
  OAI221XL \us12/U87  ( .A0(\us12/n26 ), .A1(\us12/n27 ), .B0(\us12/n28 ), 
        .B1(\us12/n20 ), .C0(\us12/n29 ), .Y(\us12/n15 ) );
  OAI221XL \us12/U86  ( .A0(\us12/n18 ), .A1(\us12/n19 ), .B0(\us12/n20 ), 
        .B1(\us12/n21 ), .C0(\us12/n22 ), .Y(\us12/n17 ) );
  AOI22X1 \us12/U85  ( .A0(\us12/n14 ), .A1(\us12/n15 ), .B0(\us12/n16 ), .B1(
        \us12/n17 ), .Y(\us12/n13 ) );
  OAI221XL \us12/U84  ( .A0(\us12/n9 ), .A1(\us12/n10 ), .B0(\us12/n11 ), .B1(
        \us12/n12 ), .C0(\us12/n13 ), .Y(\us12/n8 ) );
  MX2X1 \us12/U83  ( .A(\us12/n7 ), .B(\us12/n8 ), .S0(sa12[6]), .Y(sa11_sr[7]) );
  NOR2X4 \us12/U82  ( .A(\us12/n129 ), .B(sa12[2]), .Y(\us12/n43 ) );
  CLKINVX3 \us12/U81  ( .A(\us12/n14 ), .Y(\us12/n52 ) );
  OAI22XL \us12/U80  ( .A0(\us12/n201 ), .A1(\us12/n52 ), .B0(\us12/n202 ), 
        .B1(\us12/n114 ), .Y(\us12/n193 ) );
  CLKINVX3 \us12/U79  ( .A(sa12[5]), .Y(\us12/n252 ) );
  NOR2X2 \us12/U78  ( .A(\us12/n252 ), .B(\us12/n234 ), .Y(\us12/n55 ) );
  CLKINVX3 \us12/U77  ( .A(sa12[7]), .Y(\us12/n129 ) );
  NOR2X4 \us12/U76  ( .A(\us12/n129 ), .B(\us12/n69 ), .Y(\us12/n24 ) );
  AOI22XL \us12/U75  ( .A0(\us12/n70 ), .A1(\us12/n24 ), .B0(\us12/n96 ), .B1(
        \us12/n129 ), .Y(\us12/n241 ) );
  NOR2X2 \us12/U74  ( .A(\us12/n252 ), .B(sa12[0]), .Y(\us12/n89 ) );
  CLKINVX3 \us12/U73  ( .A(sa12[0]), .Y(\us12/n234 ) );
  NOR2X4 \us12/U72  ( .A(\us12/n69 ), .B(sa12[7]), .Y(\us12/n33 ) );
  INVX12 \us12/U71  ( .A(\us12/n33 ), .Y(\us12/n27 ) );
  CLKINVX3 \us12/U70  ( .A(\us12/n1 ), .Y(\us12/n6 ) );
  CLKINVX3 \us12/U69  ( .A(\us12/n1 ), .Y(\us12/n5 ) );
  INVXL \us12/U68  ( .A(\us12/n24 ), .Y(\us12/n36 ) );
  INVX4 \us12/U67  ( .A(\us12/n3 ), .Y(\us12/n4 ) );
  INVXL \us12/U66  ( .A(\us12/n36 ), .Y(\us12/n3 ) );
  INVX4 \us12/U65  ( .A(sa12[1]), .Y(\us12/n226 ) );
  INVX4 \us12/U64  ( .A(\us12/n43 ), .Y(\us12/n20 ) );
  AOI221X4 \us12/U63  ( .A0(\us12/n24 ), .A1(\us12/n82 ), .B0(\us12/n43 ), 
        .B1(\us12/n295 ), .C0(\us12/n173 ), .Y(\us12/n346 ) );
  AOI221X4 \us12/U62  ( .A0(\us12/n5 ), .A1(\us12/n96 ), .B0(\us12/n43 ), .B1(
        \us12/n239 ), .C0(\us12/n340 ), .Y(\us12/n336 ) );
  AOI222X4 \us12/U61  ( .A0(\us12/n59 ), .A1(\us12/n43 ), .B0(\us12/n6 ), .B1(
        \us12/n221 ), .C0(\us12/n222 ), .C1(\us12/n187 ), .Y(\us12/n218 ) );
  AOI222X4 \us12/U60  ( .A0(\us12/n123 ), .A1(\us12/n43 ), .B0(sa12[2]), .B1(
        \us12/n203 ), .C0(\us12/n6 ), .C1(\us12/n71 ), .Y(\us12/n202 ) );
  AOI221X4 \us12/U59  ( .A0(\us12/n314 ), .A1(\us12/n43 ), .B0(\us12/n160 ), 
        .B1(\us12/n24 ), .C0(\us12/n315 ), .Y(\us12/n307 ) );
  AOI221X4 \us12/U58  ( .A0(\us12/n43 ), .A1(\us12/n208 ), .B0(\us12/n76 ), 
        .B1(\us12/n24 ), .C0(\us12/n209 ), .Y(\us12/n207 ) );
  AOI221X4 \us12/U57  ( .A0(\us12/n43 ), .A1(\us12/n205 ), .B0(\us12/n32 ), 
        .B1(\us12/n6 ), .C0(\us12/n206 ), .Y(\us12/n201 ) );
  AOI221X4 \us12/U56  ( .A0(\us12/n43 ), .A1(\us12/n44 ), .B0(\us12/n45 ), 
        .B1(\us12/n24 ), .C0(\us12/n46 ), .Y(\us12/n9 ) );
  AOI22XL \us12/U55  ( .A0(\us12/n217 ), .A1(\us12/n43 ), .B0(\us12/n33 ), 
        .B1(\us12/n47 ), .Y(\us12/n216 ) );
  AOI22XL \us12/U54  ( .A0(\us12/n98 ), .A1(\us12/n43 ), .B0(\us12/n6 ), .B1(
        \us12/n99 ), .Y(\us12/n97 ) );
  AOI22XL \us12/U53  ( .A0(\us12/n82 ), .A1(\us12/n43 ), .B0(\us12/n83 ), .B1(
        \us12/n24 ), .Y(\us12/n81 ) );
  AOI2BB2XL \us12/U52  ( .B0(\us12/n43 ), .B1(\us12/n94 ), .A0N(\us12/n120 ), 
        .A1N(\us12/n4 ), .Y(\us12/n119 ) );
  AOI222X4 \us12/U51  ( .A0(\us12/n125 ), .A1(\us12/n33 ), .B0(\us12/n145 ), 
        .B1(\us12/n40 ), .C0(\us12/n43 ), .C1(\us12/n184 ), .Y(\us12/n183 ) );
  AOI22XL \us12/U50  ( .A0(\us12/n43 ), .A1(\us12/n303 ), .B0(\us12/n24 ), 
        .B1(\us12/n96 ), .Y(\us12/n358 ) );
  AOI22XL \us12/U49  ( .A0(\us12/n43 ), .A1(\us12/n100 ), .B0(\us12/n24 ), 
        .B1(\us12/n125 ), .Y(\us12/n124 ) );
  AOI21XL \us12/U48  ( .A0(\us12/n159 ), .A1(\us12/n43 ), .B0(\us12/n40 ), .Y(
        \us12/n262 ) );
  AOI22XL \us12/U47  ( .A0(\us12/n40 ), .A1(\us12/n94 ), .B0(\us12/n43 ), .B1(
        \us12/n187 ), .Y(\us12/n244 ) );
  AOI22XL \us12/U46  ( .A0(\us12/n184 ), .A1(\us12/n5 ), .B0(\us12/n198 ), 
        .B1(\us12/n43 ), .Y(\us12/n197 ) );
  NOR2XL \us12/U45  ( .A(\us12/n33 ), .B(\us12/n2 ), .Y(\us12/n302 ) );
  MXI2XL \us12/U44  ( .A(\us12/n2 ), .B(\us12/n6 ), .S0(\us12/n28 ), .Y(
        \us12/n311 ) );
  INVXL \us12/U43  ( .A(\us12/n20 ), .Y(\us12/n2 ) );
  INVX4 \us12/U42  ( .A(\us12/n6 ), .Y(\us12/n18 ) );
  AOI21XL \us12/U41  ( .A0(\us12/n18 ), .A1(\us12/n162 ), .B0(\us12/n25 ), .Y(
        \us12/n161 ) );
  INVX4 \us12/U40  ( .A(sa12[2]), .Y(\us12/n69 ) );
  NOR2X4 \us12/U39  ( .A(\us12/n226 ), .B(\us12/n4 ), .Y(\us12/n40 ) );
  CLKINVX3 \us12/U38  ( .A(sa12[3]), .Y(\us12/n136 ) );
  NOR2X2 \us12/U37  ( .A(\us12/n136 ), .B(sa12[4]), .Y(\us12/n145 ) );
  CLKINVX3 \us12/U36  ( .A(sa12[4]), .Y(\us12/n58 ) );
  NOR2X2 \us12/U35  ( .A(\us12/n58 ), .B(sa12[3]), .Y(\us12/n159 ) );
  NOR2X2 \us12/U34  ( .A(\us12/n136 ), .B(\us12/n58 ), .Y(\us12/n259 ) );
  NOR2X2 \us12/U33  ( .A(sa12[4]), .B(sa12[3]), .Y(\us12/n278 ) );
  NOR2X2 \us12/U32  ( .A(\us12/n259 ), .B(\us12/n278 ), .Y(\us12/n47 ) );
  CLKINVX3 \us12/U31  ( .A(\us12/n259 ), .Y(\us12/n44 ) );
  NOR2X2 \us12/U30  ( .A(\us12/n44 ), .B(sa12[1]), .Y(\us12/n137 ) );
  AOI21XL \us12/U29  ( .A0(\us12/n44 ), .A1(\us12/n111 ), .B0(\us12/n4 ), .Y(
        \us12/n177 ) );
  AOI22XL \us12/U28  ( .A0(\us12/n23 ), .A1(\us12/n24 ), .B0(\us12/n25 ), .B1(
        sa12[2]), .Y(\us12/n22 ) );
  AOI22XL \us12/U27  ( .A0(\us12/n33 ), .A1(sa12[3]), .B0(\us12/n24 ), .B1(
        \us12/n58 ), .Y(\us12/n277 ) );
  NAND2XL \us12/U26  ( .A(\us12/n198 ), .B(\us12/n24 ), .Y(\us12/n132 ) );
  OAI2BB2XL \us12/U25  ( .B0(\us12/n20 ), .B1(\us12/n111 ), .A0N(\us12/n125 ), 
        .A1N(\us12/n24 ), .Y(\us12/n220 ) );
  NAND2XL \us12/U24  ( .A(\us12/n111 ), .B(\us12/n101 ), .Y(\us12/n21 ) );
  NAND2XL \us12/U23  ( .A(\us12/n111 ), .B(\us12/n300 ), .Y(\us12/n187 ) );
  NAND2XL \us12/U22  ( .A(\us12/n111 ), .B(\us12/n121 ), .Y(\us12/n303 ) );
  AOI221XL \us12/U21  ( .A0(\us12/n43 ), .A1(\us12/n151 ), .B0(\us12/n25 ), 
        .B1(\us12/n69 ), .C0(\us12/n275 ), .Y(\us12/n274 ) );
  NOR2BXL \us12/U20  ( .AN(\us12/n101 ), .B(\us12/n25 ), .Y(\us12/n172 ) );
  NAND2X2 \us12/U19  ( .A(\us12/n58 ), .B(\us12/n226 ), .Y(\us12/n34 ) );
  OAI222X1 \us12/U18  ( .A0(\us12/n27 ), .A1(\us12/n34 ), .B0(\us12/n69 ), 
        .B1(\us12/n205 ), .C0(\us12/n20 ), .C1(\us12/n79 ), .Y(\us12/n260 ) );
  OAI222X1 \us12/U17  ( .A0(\us12/n20 ), .A1(\us12/n99 ), .B0(\us12/n27 ), 
        .B1(\us12/n101 ), .C0(\us12/n184 ), .C1(\us12/n4 ), .Y(\us12/n250 ) );
  OAI222X1 \us12/U16  ( .A0(\us12/n4 ), .A1(\us12/n37 ), .B0(\us12/n38 ), .B1(
        \us12/n20 ), .C0(sa12[4]), .C1(\us12/n39 ), .Y(\us12/n35 ) );
  AOI221X1 \us12/U15  ( .A0(\us12/n5 ), .A1(\us12/n19 ), .B0(\us12/n33 ), .B1(
        \us12/n34 ), .C0(\us12/n35 ), .Y(\us12/n11 ) );
  OR2X2 \us12/U14  ( .A(sa12[2]), .B(sa12[7]), .Y(\us12/n1 ) );
  AOI221XL \us12/U13  ( .A0(\us12/n70 ), .A1(\us12/n43 ), .B0(\us12/n24 ), 
        .B1(\us12/n71 ), .C0(\us12/n72 ), .Y(\us12/n53 ) );
  AOI221XL \us12/U12  ( .A0(\us12/n59 ), .A1(\us12/n33 ), .B0(\us12/n43 ), 
        .B1(\us12/n126 ), .C0(\us12/n127 ), .Y(\us12/n113 ) );
  AOI222XL \us12/U11  ( .A0(\us12/n185 ), .A1(\us12/n43 ), .B0(\us12/n186 ), 
        .B1(\us12/n187 ), .C0(\us12/n6 ), .C1(\us12/n188 ), .Y(\us12/n164 ) );
  AOI221X1 \us12/U10  ( .A0(\us12/n313 ), .A1(\us12/n5 ), .B0(\us12/n23 ), 
        .B1(\us12/n2 ), .C0(\us12/n328 ), .Y(\us12/n320 ) );
  AOI221X1 \us12/U9  ( .A0(\us12/n40 ), .A1(\us12/n136 ), .B0(\us12/n33 ), 
        .B1(\us12/n178 ), .C0(\us12/n338 ), .Y(\us12/n337 ) );
  AOI222XL \us12/U8  ( .A0(\us12/n278 ), .A1(\us12/n24 ), .B0(\us12/n42 ), 
        .B1(\us12/n33 ), .C0(\us12/n43 ), .C1(\us12/n136 ), .Y(\us12/n351 ) );
  AOI31X1 \us12/U7  ( .A0(sa12[2]), .A1(\us12/n58 ), .A2(sa12[1]), .B0(
        \us12/n40 ), .Y(\us12/n350 ) );
  AOI31X1 \us12/U6  ( .A0(\us12/n44 ), .A1(\us12/n129 ), .A2(\us12/n130 ), 
        .B0(\us12/n131 ), .Y(\us12/n128 ) );
  AOI221X1 \us12/U5  ( .A0(\us12/n40 ), .A1(\us12/n136 ), .B0(\us12/n33 ), 
        .B1(\us12/n47 ), .C0(\us12/n156 ), .Y(\us12/n141 ) );
  OAI32X1 \us12/U4  ( .A0(\us12/n18 ), .A1(sa12[1]), .A2(\us12/n159 ), .B0(
        sa12[4]), .B1(\us12/n182 ), .Y(\us12/n318 ) );
  OAI32X1 \us12/U3  ( .A0(\us12/n210 ), .A1(\us12/n145 ), .A2(\us12/n18 ), 
        .B0(\us12/n27 ), .B1(\us12/n211 ), .Y(\us12/n209 ) );
  AOI221X1 \us12/U2  ( .A0(\us12/n278 ), .A1(\us12/n40 ), .B0(\us12/n185 ), 
        .B1(\us12/n2 ), .C0(\us12/n279 ), .Y(\us12/n273 ) );
  AOI31XL \us12/U1  ( .A0(\us12/n79 ), .A1(\us12/n44 ), .A2(\us12/n2 ), .B0(
        \us12/n280 ), .Y(\us12/n339 ) );
  NAND2X1 \us13/U366  ( .A(\us13/n47 ), .B(\us13/n226 ), .Y(\us13/n189 ) );
  NOR2X1 \us13/U365  ( .A(\us13/n226 ), .B(sa13[3]), .Y(\us13/n242 ) );
  INVX1 \us13/U364  ( .A(\us13/n242 ), .Y(\us13/n205 ) );
  AND2X1 \us13/U363  ( .A(\us13/n189 ), .B(\us13/n205 ), .Y(\us13/n65 ) );
  NOR2X1 \us13/U362  ( .A(\us13/n226 ), .B(\us13/n47 ), .Y(\us13/n45 ) );
  NOR2X1 \us13/U361  ( .A(\us13/n259 ), .B(\us13/n45 ), .Y(\us13/n73 ) );
  NAND2BX1 \us13/U360  ( .AN(\us13/n73 ), .B(\us13/n6 ), .Y(\us13/n158 ) );
  NOR2X1 \us13/U359  ( .A(\us13/n226 ), .B(\us13/n159 ), .Y(\us13/n95 ) );
  INVX1 \us13/U358  ( .A(\us13/n95 ), .Y(\us13/n111 ) );
  NOR2X1 \us13/U357  ( .A(\us13/n145 ), .B(sa13[1]), .Y(\us13/n42 ) );
  INVX1 \us13/U356  ( .A(\us13/n42 ), .Y(\us13/n121 ) );
  INVX1 \us13/U355  ( .A(\us13/n47 ), .Y(\us13/n96 ) );
  OAI211X1 \us13/U354  ( .A0(\us13/n65 ), .A1(\us13/n27 ), .B0(\us13/n158 ), 
        .C0(\us13/n358 ), .Y(\us13/n355 ) );
  NOR2X1 \us13/U353  ( .A(\us13/n226 ), .B(\us13/n145 ), .Y(\us13/n59 ) );
  NOR2X1 \us13/U352  ( .A(\us13/n96 ), .B(\us13/n59 ), .Y(\us13/n271 ) );
  NOR2X1 \us13/U351  ( .A(\us13/n226 ), .B(\us13/n278 ), .Y(\us13/n217 ) );
  INVX1 \us13/U350  ( .A(\us13/n217 ), .Y(\us13/n150 ) );
  NAND2X1 \us13/U349  ( .A(\us13/n44 ), .B(\us13/n150 ), .Y(\us13/n147 ) );
  NAND2X1 \us13/U348  ( .A(sa13[4]), .B(\us13/n226 ), .Y(\us13/n101 ) );
  INVX1 \us13/U347  ( .A(\us13/n159 ), .Y(\us13/n188 ) );
  NOR2X1 \us13/U346  ( .A(\us13/n188 ), .B(\us13/n226 ), .Y(\us13/n25 ) );
  INVX1 \us13/U345  ( .A(\us13/n172 ), .Y(\us13/n107 ) );
  AOI22X1 \us13/U344  ( .A0(\us13/n33 ), .A1(\us13/n147 ), .B0(\us13/n24 ), 
        .B1(\us13/n107 ), .Y(\us13/n357 ) );
  OAI221XL \us13/U343  ( .A0(\us13/n18 ), .A1(\us13/n121 ), .B0(\us13/n271 ), 
        .B1(\us13/n20 ), .C0(\us13/n357 ), .Y(\us13/n356 ) );
  MXI2X1 \us13/U342  ( .A(\us13/n355 ), .B(\us13/n356 ), .S0(\us13/n252 ), .Y(
        \us13/n331 ) );
  INVX1 \us13/U341  ( .A(\us13/n59 ), .Y(\us13/n79 ) );
  AND2X1 \us13/U340  ( .A(\us13/n101 ), .B(\us13/n79 ), .Y(\us13/n325 ) );
  XNOR2X1 \us13/U339  ( .A(sa13[5]), .B(\us13/n226 ), .Y(\us13/n352 ) );
  NOR2X1 \us13/U338  ( .A(\us13/n226 ), .B(\us13/n136 ), .Y(\us13/n281 ) );
  INVX1 \us13/U337  ( .A(\us13/n281 ), .Y(\us13/n19 ) );
  NAND2X1 \us13/U336  ( .A(\us13/n145 ), .B(\us13/n226 ), .Y(\us13/n223 ) );
  AOI21X1 \us13/U335  ( .A0(\us13/n19 ), .A1(\us13/n223 ), .B0(\us13/n27 ), 
        .Y(\us13/n354 ) );
  AOI31X1 \us13/U334  ( .A0(\us13/n6 ), .A1(\us13/n352 ), .A2(\us13/n259 ), 
        .B0(\us13/n354 ), .Y(\us13/n353 ) );
  OAI221XL \us13/U333  ( .A0(\us13/n20 ), .A1(\us13/n34 ), .B0(\us13/n325 ), 
        .B1(\us13/n4 ), .C0(\us13/n353 ), .Y(\us13/n347 ) );
  INVX1 \us13/U332  ( .A(\us13/n352 ), .Y(\us13/n349 ) );
  NAND2X1 \us13/U331  ( .A(\us13/n278 ), .B(\us13/n6 ), .Y(\us13/n74 ) );
  OAI211X1 \us13/U330  ( .A0(\us13/n349 ), .A1(\us13/n74 ), .B0(\us13/n350 ), 
        .C0(\us13/n351 ), .Y(\us13/n348 ) );
  MXI2X1 \us13/U329  ( .A(\us13/n347 ), .B(\us13/n348 ), .S0(\us13/n252 ), .Y(
        \us13/n332 ) );
  NOR2X1 \us13/U328  ( .A(\us13/n44 ), .B(\us13/n226 ), .Y(\us13/n157 ) );
  INVX1 \us13/U327  ( .A(\us13/n157 ), .Y(\us13/n240 ) );
  NAND2X1 \us13/U326  ( .A(\us13/n240 ), .B(\us13/n189 ), .Y(\us13/n68 ) );
  NOR2X1 \us13/U325  ( .A(\us13/n20 ), .B(\us13/n159 ), .Y(\us13/n225 ) );
  NOR2X1 \us13/U324  ( .A(\us13/n225 ), .B(\us13/n40 ), .Y(\us13/n345 ) );
  INVX1 \us13/U323  ( .A(\us13/n278 ), .Y(\us13/n94 ) );
  NAND2X1 \us13/U322  ( .A(\us13/n94 ), .B(\us13/n226 ), .Y(\us13/n199 ) );
  NAND2X1 \us13/U321  ( .A(\us13/n199 ), .B(\us13/n205 ), .Y(\us13/n82 ) );
  NAND2X1 \us13/U320  ( .A(\us13/n19 ), .B(\us13/n199 ), .Y(\us13/n295 ) );
  NOR2X1 \us13/U319  ( .A(\us13/n226 ), .B(\us13/n259 ), .Y(\us13/n210 ) );
  NOR2X1 \us13/U318  ( .A(\us13/n27 ), .B(\us13/n210 ), .Y(\us13/n173 ) );
  MXI2X1 \us13/U317  ( .A(\us13/n345 ), .B(\us13/n346 ), .S0(\us13/n252 ), .Y(
        \us13/n342 ) );
  NOR2X1 \us13/U316  ( .A(sa13[1]), .B(sa13[3]), .Y(\us13/n163 ) );
  INVX1 \us13/U315  ( .A(\us13/n163 ), .Y(\us13/n37 ) );
  INVX1 \us13/U314  ( .A(\us13/n173 ), .Y(\us13/n344 ) );
  AOI21X1 \us13/U313  ( .A0(\us13/n240 ), .A1(\us13/n37 ), .B0(\us13/n344 ), 
        .Y(\us13/n343 ) );
  AOI211X1 \us13/U312  ( .A0(\us13/n5 ), .A1(\us13/n68 ), .B0(\us13/n342 ), 
        .C0(\us13/n343 ), .Y(\us13/n333 ) );
  NOR2X1 \us13/U311  ( .A(\us13/n18 ), .B(\us13/n226 ), .Y(\us13/n258 ) );
  NAND2X1 \us13/U310  ( .A(\us13/n278 ), .B(sa13[1]), .Y(\us13/n204 ) );
  NOR2X1 \us13/U309  ( .A(\us13/n188 ), .B(sa13[1]), .Y(\us13/n179 ) );
  INVX1 \us13/U308  ( .A(\us13/n179 ), .Y(\us13/n330 ) );
  NAND2X1 \us13/U307  ( .A(\us13/n204 ), .B(\us13/n330 ), .Y(\us13/n239 ) );
  NOR2X1 \us13/U306  ( .A(\us13/n136 ), .B(sa13[1]), .Y(\us13/n299 ) );
  NOR2X1 \us13/U305  ( .A(\us13/n299 ), .B(\us13/n210 ), .Y(\us13/n341 ) );
  OAI32X1 \us13/U304  ( .A0(\us13/n27 ), .A1(\us13/n278 ), .A2(\us13/n95 ), 
        .B0(\us13/n341 ), .B1(\us13/n4 ), .Y(\us13/n340 ) );
  INVX1 \us13/U303  ( .A(\us13/n45 ), .Y(\us13/n126 ) );
  NAND2X1 \us13/U302  ( .A(\us13/n126 ), .B(\us13/n101 ), .Y(\us13/n178 ) );
  NOR2X1 \us13/U301  ( .A(\us13/n18 ), .B(\us13/n136 ), .Y(\us13/n280 ) );
  OAI21XL \us13/U300  ( .A0(\us13/n4 ), .A1(\us13/n121 ), .B0(\us13/n339 ), 
        .Y(\us13/n338 ) );
  MXI2X1 \us13/U299  ( .A(\us13/n336 ), .B(\us13/n337 ), .S0(\us13/n252 ), .Y(
        \us13/n335 ) );
  NOR2X1 \us13/U298  ( .A(\us13/n258 ), .B(\us13/n335 ), .Y(\us13/n334 ) );
  MX4X1 \us13/U297  ( .A(\us13/n331 ), .B(\us13/n332 ), .C(\us13/n333 ), .D(
        \us13/n334 ), .S0(sa13[6]), .S1(\us13/n234 ), .Y(sa12_sr[0]) );
  INVX1 \us13/U296  ( .A(\us13/n299 ), .Y(\us13/n80 ) );
  NOR2X1 \us13/U295  ( .A(\us13/n111 ), .B(\us13/n18 ), .Y(\us13/n269 ) );
  INVX1 \us13/U294  ( .A(\us13/n269 ), .Y(\us13/n75 ) );
  OAI221XL \us13/U293  ( .A0(\us13/n18 ), .A1(\us13/n330 ), .B0(\us13/n20 ), 
        .B1(\us13/n80 ), .C0(\us13/n75 ), .Y(\us13/n329 ) );
  AOI221X1 \us13/U292  ( .A0(\us13/n325 ), .A1(\us13/n33 ), .B0(\us13/n24 ), 
        .B1(\us13/n303 ), .C0(\us13/n329 ), .Y(\us13/n319 ) );
  NOR2X1 \us13/U291  ( .A(\us13/n234 ), .B(sa13[5]), .Y(\us13/n14 ) );
  NOR2X1 \us13/U290  ( .A(\us13/n25 ), .B(\us13/n299 ), .Y(\us13/n313 ) );
  NAND2X1 \us13/U289  ( .A(\us13/n44 ), .B(\us13/n226 ), .Y(\us13/n300 ) );
  AND2X1 \us13/U288  ( .A(\us13/n300 ), .B(\us13/n240 ), .Y(\us13/n23 ) );
  OAI32X1 \us13/U287  ( .A0(\us13/n4 ), .A1(\us13/n145 ), .A2(\us13/n210 ), 
        .B0(\us13/n137 ), .B1(\us13/n27 ), .Y(\us13/n328 ) );
  NOR2X1 \us13/U286  ( .A(sa13[0]), .B(sa13[5]), .Y(\us13/n16 ) );
  INVX1 \us13/U285  ( .A(\us13/n16 ), .Y(\us13/n114 ) );
  INVX1 \us13/U284  ( .A(\us13/n145 ), .Y(\us13/n149 ) );
  NOR2X1 \us13/U283  ( .A(\us13/n47 ), .B(sa13[1]), .Y(\us13/n98 ) );
  INVX1 \us13/U282  ( .A(\us13/n98 ), .Y(\us13/n284 ) );
  OAI21XL \us13/U281  ( .A0(\us13/n69 ), .A1(\us13/n284 ), .B0(\us13/n27 ), 
        .Y(\us13/n327 ) );
  AOI31X1 \us13/U280  ( .A0(\us13/n111 ), .A1(\us13/n149 ), .A2(\us13/n327 ), 
        .B0(\us13/n225 ), .Y(\us13/n326 ) );
  OAI21XL \us13/U279  ( .A0(\us13/n325 ), .A1(\us13/n18 ), .B0(\us13/n326 ), 
        .Y(\us13/n322 ) );
  NAND2X1 \us13/U278  ( .A(\us13/n19 ), .B(\us13/n189 ), .Y(\us13/n71 ) );
  NOR2X1 \us13/U277  ( .A(\us13/n71 ), .B(\us13/n18 ), .Y(\us13/n135 ) );
  AOI21X1 \us13/U276  ( .A0(\us13/n40 ), .A1(sa13[4]), .B0(\us13/n135 ), .Y(
        \us13/n324 ) );
  OAI221XL \us13/U275  ( .A0(\us13/n47 ), .A1(\us13/n27 ), .B0(\us13/n65 ), 
        .B1(\us13/n20 ), .C0(\us13/n324 ), .Y(\us13/n323 ) );
  AOI22X1 \us13/U274  ( .A0(\us13/n55 ), .A1(\us13/n322 ), .B0(\us13/n89 ), 
        .B1(\us13/n323 ), .Y(\us13/n321 ) );
  OAI221XL \us13/U273  ( .A0(\us13/n319 ), .A1(\us13/n52 ), .B0(\us13/n320 ), 
        .B1(\us13/n114 ), .C0(\us13/n321 ), .Y(\us13/n304 ) );
  NOR2X1 \us13/U272  ( .A(\us13/n226 ), .B(\us13/n58 ), .Y(\us13/n290 ) );
  INVX1 \us13/U271  ( .A(\us13/n290 ), .Y(\us13/n200 ) );
  NAND2X1 \us13/U270  ( .A(\us13/n34 ), .B(\us13/n200 ), .Y(\us13/n120 ) );
  INVX1 \us13/U269  ( .A(\us13/n210 ), .Y(\us13/n100 ) );
  OAI221XL \us13/U268  ( .A0(\us13/n20 ), .A1(\us13/n100 ), .B0(sa13[3]), .B1(
        \us13/n4 ), .C0(\us13/n262 ), .Y(\us13/n317 ) );
  INVX1 \us13/U267  ( .A(\us13/n258 ), .Y(\us13/n182 ) );
  AOI211X1 \us13/U266  ( .A0(\us13/n33 ), .A1(\us13/n120 ), .B0(\us13/n317 ), 
        .C0(\us13/n318 ), .Y(\us13/n306 ) );
  NAND2X1 \us13/U265  ( .A(\us13/n100 ), .B(\us13/n199 ), .Y(\us13/n151 ) );
  INVX1 \us13/U264  ( .A(\us13/n151 ), .Y(\us13/n314 ) );
  NOR2X1 \us13/U263  ( .A(\us13/n45 ), .B(\us13/n163 ), .Y(\us13/n160 ) );
  INVX1 \us13/U262  ( .A(\us13/n295 ), .Y(\us13/n92 ) );
  AOI21X1 \us13/U261  ( .A0(sa13[1]), .A1(\us13/n58 ), .B0(\us13/n98 ), .Y(
        \us13/n316 ) );
  OAI22X1 \us13/U260  ( .A0(\us13/n92 ), .A1(\us13/n18 ), .B0(\us13/n316 ), 
        .B1(\us13/n27 ), .Y(\us13/n315 ) );
  NOR2X1 \us13/U259  ( .A(\us13/n149 ), .B(\us13/n226 ), .Y(\us13/n41 ) );
  INVX1 \us13/U258  ( .A(\us13/n41 ), .Y(\us13/n105 ) );
  NAND2X1 \us13/U257  ( .A(\us13/n284 ), .B(\us13/n105 ), .Y(\us13/n227 ) );
  AOI21X1 \us13/U256  ( .A0(\us13/n313 ), .A1(\us13/n33 ), .B0(\us13/n269 ), 
        .Y(\us13/n312 ) );
  OAI221XL \us13/U255  ( .A0(\us13/n149 ), .A1(\us13/n20 ), .B0(\us13/n4 ), 
        .B1(\us13/n227 ), .C0(\us13/n312 ), .Y(\us13/n309 ) );
  AOI21X1 \us13/U254  ( .A0(\us13/n226 ), .A1(\us13/n188 ), .B0(\us13/n242 ), 
        .Y(\us13/n185 ) );
  INVX1 \us13/U253  ( .A(\us13/n185 ), .Y(\us13/n48 ) );
  AND2X1 \us13/U252  ( .A(\us13/n223 ), .B(\us13/n240 ), .Y(\us13/n28 ) );
  OAI221XL \us13/U251  ( .A0(\us13/n27 ), .A1(\us13/n44 ), .B0(\us13/n4 ), 
        .B1(\us13/n48 ), .C0(\us13/n311 ), .Y(\us13/n310 ) );
  AOI22X1 \us13/U250  ( .A0(\us13/n89 ), .A1(\us13/n309 ), .B0(\us13/n55 ), 
        .B1(\us13/n310 ), .Y(\us13/n308 ) );
  OAI221XL \us13/U249  ( .A0(\us13/n306 ), .A1(\us13/n52 ), .B0(\us13/n307 ), 
        .B1(\us13/n114 ), .C0(\us13/n308 ), .Y(\us13/n305 ) );
  MX2X1 \us13/U248  ( .A(\us13/n304 ), .B(\us13/n305 ), .S0(sa13[6]), .Y(
        sa12_sr[1]) );
  INVX1 \us13/U247  ( .A(\us13/n187 ), .Y(\us13/n61 ) );
  MXI2X1 \us13/U246  ( .A(\us13/n303 ), .B(\us13/n61 ), .S0(\us13/n69 ), .Y(
        \us13/n301 ) );
  MXI2X1 \us13/U245  ( .A(\us13/n301 ), .B(\us13/n147 ), .S0(\us13/n302 ), .Y(
        \us13/n285 ) );
  NAND2X1 \us13/U244  ( .A(\us13/n200 ), .B(\us13/n300 ), .Y(\us13/n99 ) );
  INVX1 \us13/U243  ( .A(\us13/n99 ), .Y(\us13/n296 ) );
  NOR2X1 \us13/U242  ( .A(\us13/n299 ), .B(\us13/n242 ), .Y(\us13/n298 ) );
  NAND2X1 \us13/U241  ( .A(sa13[1]), .B(\us13/n47 ), .Y(\us13/n122 ) );
  NOR2X1 \us13/U240  ( .A(\us13/n159 ), .B(\us13/n217 ), .Y(\us13/n198 ) );
  OAI221XL \us13/U239  ( .A0(\us13/n298 ), .A1(\us13/n27 ), .B0(\us13/n20 ), 
        .B1(\us13/n122 ), .C0(\us13/n132 ), .Y(\us13/n297 ) );
  AOI221X1 \us13/U238  ( .A0(\us13/n225 ), .A1(\us13/n226 ), .B0(\us13/n296 ), 
        .B1(\us13/n6 ), .C0(\us13/n297 ), .Y(\us13/n291 ) );
  OAI2BB2X1 \us13/U237  ( .B0(\us13/n27 ), .B1(\us13/n295 ), .A0N(\us13/n34 ), 
        .A1N(\us13/n24 ), .Y(\us13/n293 ) );
  AOI21X1 \us13/U236  ( .A0(\us13/n101 ), .A1(\us13/n150 ), .B0(\us13/n20 ), 
        .Y(\us13/n294 ) );
  AOI211X1 \us13/U235  ( .A0(\us13/n5 ), .A1(\us13/n79 ), .B0(\us13/n293 ), 
        .C0(\us13/n294 ), .Y(\us13/n292 ) );
  INVX1 \us13/U234  ( .A(\us13/n89 ), .Y(\us13/n10 ) );
  OAI22X1 \us13/U233  ( .A0(\us13/n291 ), .A1(\us13/n114 ), .B0(\us13/n292 ), 
        .B1(\us13/n10 ), .Y(\us13/n286 ) );
  INVX1 \us13/U232  ( .A(\us13/n225 ), .Y(\us13/n288 ) );
  NAND2X1 \us13/U231  ( .A(\us13/n200 ), .B(\us13/n284 ), .Y(\us13/n102 ) );
  NOR2X1 \us13/U230  ( .A(\us13/n290 ), .B(\us13/n163 ), .Y(\us13/n184 ) );
  AOI22X1 \us13/U229  ( .A0(\us13/n102 ), .A1(\us13/n69 ), .B0(\us13/n184 ), 
        .B1(\us13/n33 ), .Y(\us13/n289 ) );
  AOI31X1 \us13/U228  ( .A0(\us13/n132 ), .A1(\us13/n288 ), .A2(\us13/n289 ), 
        .B0(\us13/n52 ), .Y(\us13/n287 ) );
  AOI211X1 \us13/U227  ( .A0(\us13/n285 ), .A1(\us13/n55 ), .B0(\us13/n286 ), 
        .C0(\us13/n287 ), .Y(\us13/n263 ) );
  NAND2X1 \us13/U226  ( .A(\us13/n284 ), .B(\us13/n122 ), .Y(\us13/n125 ) );
  NOR2X1 \us13/U225  ( .A(\us13/n199 ), .B(\us13/n4 ), .Y(\us13/n50 ) );
  AOI21X1 \us13/U224  ( .A0(\us13/n200 ), .A1(\us13/n223 ), .B0(\us13/n20 ), 
        .Y(\us13/n283 ) );
  AOI211X1 \us13/U223  ( .A0(\us13/n5 ), .A1(\us13/n125 ), .B0(\us13/n50 ), 
        .C0(\us13/n283 ), .Y(\us13/n282 ) );
  OAI221XL \us13/U222  ( .A0(\us13/n281 ), .A1(\us13/n27 ), .B0(\us13/n4 ), 
        .B1(\us13/n111 ), .C0(\us13/n282 ), .Y(\us13/n265 ) );
  INVX1 \us13/U221  ( .A(\us13/n280 ), .Y(\us13/n247 ) );
  NAND2X1 \us13/U220  ( .A(\us13/n41 ), .B(\us13/n33 ), .Y(\us13/n272 ) );
  OAI221XL \us13/U219  ( .A0(sa13[1]), .A1(\us13/n247 ), .B0(\us13/n4 ), .B1(
        \us13/n189 ), .C0(\us13/n272 ), .Y(\us13/n279 ) );
  NAND2X1 \us13/U218  ( .A(sa13[2]), .B(\us13/n149 ), .Y(\us13/n276 ) );
  XNOR2X1 \us13/U217  ( .A(\us13/n129 ), .B(sa13[1]), .Y(\us13/n155 ) );
  MXI2X1 \us13/U216  ( .A(\us13/n276 ), .B(\us13/n277 ), .S0(\us13/n155 ), .Y(
        \us13/n275 ) );
  OAI22X1 \us13/U215  ( .A0(\us13/n273 ), .A1(\us13/n10 ), .B0(\us13/n274 ), 
        .B1(\us13/n52 ), .Y(\us13/n266 ) );
  NOR2X1 \us13/U214  ( .A(\us13/n20 ), .B(\us13/n226 ), .Y(\us13/n176 ) );
  OAI21XL \us13/U213  ( .A0(\us13/n4 ), .A1(\us13/n271 ), .B0(\us13/n272 ), 
        .Y(\us13/n270 ) );
  OAI31X1 \us13/U212  ( .A0(\us13/n176 ), .A1(\us13/n269 ), .A2(\us13/n270 ), 
        .B0(\us13/n16 ), .Y(\us13/n268 ) );
  INVX1 \us13/U211  ( .A(\us13/n268 ), .Y(\us13/n267 ) );
  AOI211X1 \us13/U210  ( .A0(\us13/n55 ), .A1(\us13/n265 ), .B0(\us13/n266 ), 
        .C0(\us13/n267 ), .Y(\us13/n264 ) );
  MXI2X1 \us13/U209  ( .A(\us13/n263 ), .B(\us13/n264 ), .S0(sa13[6]), .Y(
        sa12_sr[2]) );
  NOR2X1 \us13/U208  ( .A(\us13/n94 ), .B(sa13[1]), .Y(\us13/n211 ) );
  INVX1 \us13/U207  ( .A(\us13/n262 ), .Y(\us13/n261 ) );
  AOI211X1 \us13/U206  ( .A0(\us13/n259 ), .A1(\us13/n24 ), .B0(\us13/n260 ), 
        .C0(\us13/n261 ), .Y(\us13/n255 ) );
  OAI22X1 \us13/U205  ( .A0(\us13/n20 ), .A1(\us13/n68 ), .B0(\us13/n27 ), 
        .B1(\us13/n37 ), .Y(\us13/n257 ) );
  NOR3X1 \us13/U204  ( .A(\us13/n257 ), .B(\us13/n258 ), .C(\us13/n50 ), .Y(
        \us13/n256 ) );
  MXI2X1 \us13/U203  ( .A(\us13/n255 ), .B(\us13/n256 ), .S0(\us13/n252 ), .Y(
        \us13/n254 ) );
  AOI221X1 \us13/U202  ( .A0(\us13/n211 ), .A1(\us13/n5 ), .B0(\us13/n40 ), 
        .B1(sa13[4]), .C0(\us13/n254 ), .Y(\us13/n248 ) );
  INVX1 \us13/U201  ( .A(\us13/n211 ), .Y(\us13/n106 ) );
  NAND2X1 \us13/U200  ( .A(\us13/n200 ), .B(\us13/n106 ), .Y(\us13/n83 ) );
  NAND2X1 \us13/U199  ( .A(\us13/n199 ), .B(\us13/n204 ), .Y(\us13/n169 ) );
  AOI2BB2X1 \us13/U198  ( .B0(\us13/n65 ), .B1(\us13/n24 ), .A0N(\us13/n169 ), 
        .A1N(\us13/n20 ), .Y(\us13/n253 ) );
  OAI221XL \us13/U197  ( .A0(\us13/n172 ), .A1(\us13/n18 ), .B0(\us13/n27 ), 
        .B1(\us13/n83 ), .C0(\us13/n253 ), .Y(\us13/n251 ) );
  MXI2X1 \us13/U196  ( .A(\us13/n250 ), .B(\us13/n251 ), .S0(\us13/n252 ), .Y(
        \us13/n249 ) );
  MXI2X1 \us13/U195  ( .A(\us13/n248 ), .B(\us13/n249 ), .S0(\us13/n234 ), .Y(
        \us13/n228 ) );
  OAI21XL \us13/U194  ( .A0(\us13/n58 ), .A1(\us13/n27 ), .B0(\us13/n247 ), 
        .Y(\us13/n245 ) );
  NOR2X1 \us13/U193  ( .A(sa13[7]), .B(\us13/n145 ), .Y(\us13/n246 ) );
  XNOR2X1 \us13/U192  ( .A(\us13/n69 ), .B(sa13[1]), .Y(\us13/n130 ) );
  MXI2X1 \us13/U191  ( .A(\us13/n245 ), .B(\us13/n246 ), .S0(\us13/n130 ), .Y(
        \us13/n243 ) );
  OAI211X1 \us13/U190  ( .A0(\us13/n4 ), .A1(\us13/n149 ), .B0(\us13/n243 ), 
        .C0(\us13/n244 ), .Y(\us13/n230 ) );
  NOR2X1 \us13/U189  ( .A(\us13/n242 ), .B(\us13/n137 ), .Y(\us13/n70 ) );
  OAI221XL \us13/U188  ( .A0(\us13/n159 ), .A1(\us13/n27 ), .B0(\us13/n20 ), 
        .B1(\us13/n34 ), .C0(\us13/n241 ), .Y(\us13/n231 ) );
  NAND2X1 \us13/U187  ( .A(\us13/n101 ), .B(\us13/n240 ), .Y(\us13/n76 ) );
  AOI21X1 \us13/U186  ( .A0(\us13/n122 ), .A1(\us13/n106 ), .B0(\us13/n129 ), 
        .Y(\us13/n237 ) );
  INVX1 \us13/U185  ( .A(\us13/n239 ), .Y(\us13/n238 ) );
  OAI21XL \us13/U184  ( .A0(\us13/n237 ), .A1(\us13/n43 ), .B0(\us13/n238 ), 
        .Y(\us13/n236 ) );
  OAI221XL \us13/U183  ( .A0(\us13/n18 ), .A1(\us13/n76 ), .B0(\us13/n59 ), 
        .B1(\us13/n27 ), .C0(\us13/n236 ), .Y(\us13/n232 ) );
  AOI2BB2X1 \us13/U182  ( .B0(\us13/n24 ), .B1(\us13/n187 ), .A0N(\us13/n227 ), 
        .A1N(\us13/n20 ), .Y(\us13/n235 ) );
  OAI211X1 \us13/U181  ( .A0(\us13/n27 ), .A1(\us13/n122 ), .B0(\us13/n158 ), 
        .C0(\us13/n235 ), .Y(\us13/n233 ) );
  MX4X1 \us13/U180  ( .A(\us13/n230 ), .B(\us13/n231 ), .C(\us13/n232 ), .D(
        \us13/n233 ), .S0(\us13/n234 ), .S1(sa13[5]), .Y(\us13/n229 ) );
  MX2X1 \us13/U179  ( .A(\us13/n228 ), .B(\us13/n229 ), .S0(sa13[6]), .Y(
        sa12_sr[3]) );
  NOR2BX1 \us13/U178  ( .AN(\us13/n204 ), .B(\us13/n137 ), .Y(\us13/n110 ) );
  INVX1 \us13/U177  ( .A(\us13/n110 ), .Y(\us13/n64 ) );
  AOI22X1 \us13/U176  ( .A0(\us13/n225 ), .A1(\us13/n226 ), .B0(\us13/n6 ), 
        .B1(\us13/n227 ), .Y(\us13/n224 ) );
  OAI221XL \us13/U175  ( .A0(\us13/n27 ), .A1(\us13/n64 ), .B0(\us13/n4 ), 
        .B1(\us13/n83 ), .C0(\us13/n224 ), .Y(\us13/n212 ) );
  NAND2X1 \us13/U174  ( .A(\us13/n34 ), .B(\us13/n204 ), .Y(\us13/n221 ) );
  OAI21XL \us13/U173  ( .A0(\us13/n69 ), .A1(\us13/n223 ), .B0(\us13/n27 ), 
        .Y(\us13/n222 ) );
  NOR2X1 \us13/U172  ( .A(\us13/n217 ), .B(\us13/n42 ), .Y(\us13/n208 ) );
  AOI211X1 \us13/U171  ( .A0(\us13/n208 ), .A1(\us13/n5 ), .B0(\us13/n220 ), 
        .C0(\us13/n173 ), .Y(\us13/n219 ) );
  OAI22X1 \us13/U170  ( .A0(\us13/n218 ), .A1(\us13/n10 ), .B0(\us13/n219 ), 
        .B1(\us13/n114 ), .Y(\us13/n213 ) );
  INVX1 \us13/U169  ( .A(\us13/n135 ), .Y(\us13/n215 ) );
  NOR2X1 \us13/U168  ( .A(\us13/n4 ), .B(\us13/n159 ), .Y(\us13/n31 ) );
  INVX1 \us13/U167  ( .A(\us13/n31 ), .Y(\us13/n196 ) );
  AOI31X1 \us13/U166  ( .A0(\us13/n215 ), .A1(\us13/n196 ), .A2(\us13/n216 ), 
        .B0(\us13/n52 ), .Y(\us13/n214 ) );
  AOI211X1 \us13/U165  ( .A0(\us13/n55 ), .A1(\us13/n212 ), .B0(\us13/n213 ), 
        .C0(\us13/n214 ), .Y(\us13/n190 ) );
  INVX1 \us13/U164  ( .A(\us13/n207 ), .Y(\us13/n192 ) );
  NOR2X1 \us13/U163  ( .A(\us13/n25 ), .B(\us13/n98 ), .Y(\us13/n32 ) );
  OAI22X1 \us13/U162  ( .A0(\us13/n28 ), .A1(\us13/n4 ), .B0(\us13/n188 ), 
        .B1(\us13/n27 ), .Y(\us13/n206 ) );
  NAND2X1 \us13/U161  ( .A(\us13/n204 ), .B(\us13/n80 ), .Y(\us13/n118 ) );
  INVX1 \us13/U160  ( .A(\us13/n118 ), .Y(\us13/n123 ) );
  NAND2X1 \us13/U159  ( .A(\us13/n94 ), .B(\us13/n79 ), .Y(\us13/n203 ) );
  OAI2BB1X1 \us13/U158  ( .A0N(\us13/n199 ), .A1N(\us13/n200 ), .B0(\us13/n33 ), .Y(\us13/n195 ) );
  INVX1 \us13/U157  ( .A(\us13/n55 ), .Y(\us13/n12 ) );
  AOI31X1 \us13/U156  ( .A0(\us13/n195 ), .A1(\us13/n196 ), .A2(\us13/n197 ), 
        .B0(\us13/n12 ), .Y(\us13/n194 ) );
  AOI211X1 \us13/U155  ( .A0(\us13/n89 ), .A1(\us13/n192 ), .B0(\us13/n193 ), 
        .C0(\us13/n194 ), .Y(\us13/n191 ) );
  MXI2X1 \us13/U154  ( .A(\us13/n190 ), .B(\us13/n191 ), .S0(sa13[6]), .Y(
        sa12_sr[4]) );
  OAI21XL \us13/U153  ( .A0(\us13/n69 ), .A1(\us13/n189 ), .B0(\us13/n27 ), 
        .Y(\us13/n186 ) );
  INVX1 \us13/U152  ( .A(\us13/n183 ), .Y(\us13/n180 ) );
  NAND2X1 \us13/U151  ( .A(\us13/n74 ), .B(\us13/n182 ), .Y(\us13/n181 ) );
  AOI211X1 \us13/U150  ( .A0(\us13/n179 ), .A1(\us13/n24 ), .B0(\us13/n180 ), 
        .C0(\us13/n181 ), .Y(\us13/n165 ) );
  INVX1 \us13/U149  ( .A(\us13/n178 ), .Y(\us13/n175 ) );
  AOI211X1 \us13/U148  ( .A0(\us13/n175 ), .A1(\us13/n5 ), .B0(\us13/n176 ), 
        .C0(\us13/n177 ), .Y(\us13/n174 ) );
  OAI221XL \us13/U147  ( .A0(\us13/n159 ), .A1(\us13/n27 ), .B0(\us13/n145 ), 
        .B1(\us13/n20 ), .C0(\us13/n174 ), .Y(\us13/n167 ) );
  MXI2X1 \us13/U146  ( .A(\us13/n40 ), .B(\us13/n173 ), .S0(\us13/n96 ), .Y(
        \us13/n170 ) );
  AOI22X1 \us13/U145  ( .A0(\us13/n137 ), .A1(\us13/n24 ), .B0(\us13/n172 ), 
        .B1(\us13/n6 ), .Y(\us13/n171 ) );
  OAI211X1 \us13/U144  ( .A0(\us13/n20 ), .A1(\us13/n169 ), .B0(\us13/n170 ), 
        .C0(\us13/n171 ), .Y(\us13/n168 ) );
  AOI22X1 \us13/U143  ( .A0(\us13/n89 ), .A1(\us13/n167 ), .B0(\us13/n55 ), 
        .B1(\us13/n168 ), .Y(\us13/n166 ) );
  OAI221XL \us13/U142  ( .A0(\us13/n164 ), .A1(\us13/n114 ), .B0(\us13/n165 ), 
        .B1(\us13/n52 ), .C0(\us13/n166 ), .Y(\us13/n138 ) );
  OAI21XL \us13/U141  ( .A0(\us13/n41 ), .A1(\us13/n163 ), .B0(\us13/n69 ), 
        .Y(\us13/n162 ) );
  AOI221X1 \us13/U140  ( .A0(\us13/n159 ), .A1(\us13/n24 ), .B0(\us13/n160 ), 
        .B1(\us13/n33 ), .C0(\us13/n161 ), .Y(\us13/n140 ) );
  OAI21XL \us13/U139  ( .A0(\us13/n157 ), .A1(\us13/n20 ), .B0(\us13/n158 ), 
        .Y(\us13/n156 ) );
  NOR2X1 \us13/U138  ( .A(\us13/n4 ), .B(\us13/n136 ), .Y(\us13/n153 ) );
  NOR2X1 \us13/U137  ( .A(\us13/n145 ), .B(\us13/n69 ), .Y(\us13/n154 ) );
  MXI2X1 \us13/U136  ( .A(\us13/n153 ), .B(\us13/n154 ), .S0(\us13/n155 ), .Y(
        \us13/n152 ) );
  OAI221XL \us13/U135  ( .A0(\us13/n110 ), .A1(\us13/n18 ), .B0(\us13/n20 ), 
        .B1(\us13/n151 ), .C0(\us13/n152 ), .Y(\us13/n143 ) );
  AOI21X1 \us13/U134  ( .A0(\us13/n149 ), .A1(\us13/n150 ), .B0(\us13/n18 ), 
        .Y(\us13/n148 ) );
  AOI2BB1X1 \us13/U133  ( .A0N(\us13/n147 ), .A1N(\us13/n27 ), .B0(\us13/n148 ), .Y(\us13/n146 ) );
  OAI221XL \us13/U132  ( .A0(\us13/n145 ), .A1(\us13/n20 ), .B0(\us13/n4 ), 
        .B1(\us13/n34 ), .C0(\us13/n146 ), .Y(\us13/n144 ) );
  AOI22X1 \us13/U131  ( .A0(\us13/n89 ), .A1(\us13/n143 ), .B0(\us13/n14 ), 
        .B1(\us13/n144 ), .Y(\us13/n142 ) );
  OAI221XL \us13/U130  ( .A0(\us13/n140 ), .A1(\us13/n12 ), .B0(\us13/n141 ), 
        .B1(\us13/n114 ), .C0(\us13/n142 ), .Y(\us13/n139 ) );
  MX2X1 \us13/U129  ( .A(\us13/n138 ), .B(\us13/n139 ), .S0(sa13[6]), .Y(
        sa12_sr[5]) );
  INVX1 \us13/U128  ( .A(\us13/n70 ), .Y(\us13/n133 ) );
  OAI22X1 \us13/U127  ( .A0(\us13/n4 ), .A1(\us13/n136 ), .B0(\us13/n137 ), 
        .B1(\us13/n27 ), .Y(\us13/n134 ) );
  AOI211X1 \us13/U126  ( .A0(\us13/n133 ), .A1(\us13/n69 ), .B0(\us13/n134 ), 
        .C0(\us13/n135 ), .Y(\us13/n112 ) );
  INVX1 \us13/U125  ( .A(\us13/n132 ), .Y(\us13/n131 ) );
  OAI21XL \us13/U124  ( .A0(\us13/n18 ), .A1(\us13/n37 ), .B0(\us13/n128 ), 
        .Y(\us13/n127 ) );
  OAI221XL \us13/U123  ( .A0(\us13/n18 ), .A1(\us13/n105 ), .B0(\us13/n123 ), 
        .B1(\us13/n27 ), .C0(\us13/n124 ), .Y(\us13/n116 ) );
  NAND2X1 \us13/U122  ( .A(\us13/n121 ), .B(\us13/n122 ), .Y(\us13/n30 ) );
  OAI221XL \us13/U121  ( .A0(\us13/n18 ), .A1(\us13/n118 ), .B0(\us13/n27 ), 
        .B1(\us13/n30 ), .C0(\us13/n119 ), .Y(\us13/n117 ) );
  AOI22X1 \us13/U120  ( .A0(\us13/n89 ), .A1(\us13/n116 ), .B0(\us13/n55 ), 
        .B1(\us13/n117 ), .Y(\us13/n115 ) );
  OAI221XL \us13/U119  ( .A0(\us13/n112 ), .A1(\us13/n52 ), .B0(\us13/n113 ), 
        .B1(\us13/n114 ), .C0(\us13/n115 ), .Y(\us13/n84 ) );
  OAI22X1 \us13/U118  ( .A0(\us13/n110 ), .A1(\us13/n4 ), .B0(\us13/n20 ), 
        .B1(\us13/n21 ), .Y(\us13/n108 ) );
  AOI21X1 \us13/U117  ( .A0(sa13[1]), .A1(\us13/n58 ), .B0(\us13/n27 ), .Y(
        \us13/n109 ) );
  AOI211X1 \us13/U116  ( .A0(\us13/n5 ), .A1(\us13/n107 ), .B0(\us13/n108 ), 
        .C0(\us13/n109 ), .Y(\us13/n86 ) );
  OAI22X1 \us13/U115  ( .A0(\us13/n45 ), .A1(\us13/n4 ), .B0(sa13[4]), .B1(
        \us13/n18 ), .Y(\us13/n103 ) );
  AOI21X1 \us13/U114  ( .A0(\us13/n105 ), .A1(\us13/n106 ), .B0(\us13/n20 ), 
        .Y(\us13/n104 ) );
  AOI211X1 \us13/U113  ( .A0(\us13/n33 ), .A1(\us13/n102 ), .B0(\us13/n103 ), 
        .C0(\us13/n104 ), .Y(\us13/n87 ) );
  NAND2X1 \us13/U112  ( .A(\us13/n100 ), .B(\us13/n101 ), .Y(\us13/n62 ) );
  OAI221XL \us13/U111  ( .A0(\us13/n27 ), .A1(\us13/n62 ), .B0(\us13/n4 ), 
        .B1(\us13/n21 ), .C0(\us13/n97 ), .Y(\us13/n90 ) );
  NOR3X1 \us13/U110  ( .A(\us13/n4 ), .B(\us13/n95 ), .C(\us13/n96 ), .Y(
        \us13/n67 ) );
  AOI31X1 \us13/U109  ( .A0(\us13/n79 ), .A1(\us13/n94 ), .A2(\us13/n6 ), .B0(
        \us13/n67 ), .Y(\us13/n93 ) );
  OAI221XL \us13/U108  ( .A0(\us13/n73 ), .A1(\us13/n27 ), .B0(\us13/n92 ), 
        .B1(\us13/n20 ), .C0(\us13/n93 ), .Y(\us13/n91 ) );
  AOI22X1 \us13/U107  ( .A0(\us13/n89 ), .A1(\us13/n90 ), .B0(\us13/n16 ), 
        .B1(\us13/n91 ), .Y(\us13/n88 ) );
  OAI221XL \us13/U106  ( .A0(\us13/n86 ), .A1(\us13/n52 ), .B0(\us13/n87 ), 
        .B1(\us13/n12 ), .C0(\us13/n88 ), .Y(\us13/n85 ) );
  MX2X1 \us13/U105  ( .A(\us13/n84 ), .B(\us13/n85 ), .S0(sa13[6]), .Y(
        sa12_sr[6]) );
  INVX1 \us13/U104  ( .A(\us13/n81 ), .Y(\us13/n77 ) );
  AOI21X1 \us13/U103  ( .A0(\us13/n79 ), .A1(\us13/n80 ), .B0(\us13/n27 ), .Y(
        \us13/n78 ) );
  AOI211X1 \us13/U102  ( .A0(\us13/n5 ), .A1(\us13/n76 ), .B0(\us13/n77 ), 
        .C0(\us13/n78 ), .Y(\us13/n51 ) );
  OAI211X1 \us13/U101  ( .A0(\us13/n73 ), .A1(\us13/n27 ), .B0(\us13/n74 ), 
        .C0(\us13/n75 ), .Y(\us13/n72 ) );
  AOI21X1 \us13/U100  ( .A0(\us13/n68 ), .A1(\us13/n69 ), .B0(\us13/n6 ), .Y(
        \us13/n63 ) );
  INVX1 \us13/U99  ( .A(\us13/n67 ), .Y(\us13/n66 ) );
  OAI221XL \us13/U98  ( .A0(\us13/n63 ), .A1(\us13/n64 ), .B0(\us13/n65 ), 
        .B1(\us13/n27 ), .C0(\us13/n66 ), .Y(\us13/n56 ) );
  AOI2BB2X1 \us13/U97  ( .B0(\us13/n61 ), .B1(\us13/n24 ), .A0N(\us13/n62 ), 
        .A1N(\us13/n20 ), .Y(\us13/n60 ) );
  OAI221XL \us13/U96  ( .A0(\us13/n58 ), .A1(\us13/n18 ), .B0(\us13/n59 ), 
        .B1(\us13/n27 ), .C0(\us13/n60 ), .Y(\us13/n57 ) );
  AOI22X1 \us13/U95  ( .A0(\us13/n55 ), .A1(\us13/n56 ), .B0(\us13/n16 ), .B1(
        \us13/n57 ), .Y(\us13/n54 ) );
  OAI221XL \us13/U94  ( .A0(\us13/n51 ), .A1(\us13/n52 ), .B0(\us13/n53 ), 
        .B1(\us13/n10 ), .C0(\us13/n54 ), .Y(\us13/n7 ) );
  INVX1 \us13/U93  ( .A(\us13/n50 ), .Y(\us13/n49 ) );
  OAI221XL \us13/U92  ( .A0(\us13/n47 ), .A1(\us13/n18 ), .B0(\us13/n27 ), 
        .B1(\us13/n48 ), .C0(\us13/n49 ), .Y(\us13/n46 ) );
  NOR2X1 \us13/U91  ( .A(\us13/n41 ), .B(\us13/n42 ), .Y(\us13/n38 ) );
  INVX1 \us13/U90  ( .A(\us13/n40 ), .Y(\us13/n39 ) );
  INVX1 \us13/U89  ( .A(\us13/n32 ), .Y(\us13/n26 ) );
  AOI21X1 \us13/U88  ( .A0(\us13/n5 ), .A1(\us13/n30 ), .B0(\us13/n31 ), .Y(
        \us13/n29 ) );
  OAI221XL \us13/U87  ( .A0(\us13/n26 ), .A1(\us13/n27 ), .B0(\us13/n28 ), 
        .B1(\us13/n20 ), .C0(\us13/n29 ), .Y(\us13/n15 ) );
  OAI221XL \us13/U86  ( .A0(\us13/n18 ), .A1(\us13/n19 ), .B0(\us13/n20 ), 
        .B1(\us13/n21 ), .C0(\us13/n22 ), .Y(\us13/n17 ) );
  AOI22X1 \us13/U85  ( .A0(\us13/n14 ), .A1(\us13/n15 ), .B0(\us13/n16 ), .B1(
        \us13/n17 ), .Y(\us13/n13 ) );
  OAI221XL \us13/U84  ( .A0(\us13/n9 ), .A1(\us13/n10 ), .B0(\us13/n11 ), .B1(
        \us13/n12 ), .C0(\us13/n13 ), .Y(\us13/n8 ) );
  MX2X1 \us13/U83  ( .A(\us13/n7 ), .B(\us13/n8 ), .S0(sa13[6]), .Y(sa12_sr[7]) );
  NOR2X4 \us13/U82  ( .A(\us13/n129 ), .B(sa13[2]), .Y(\us13/n43 ) );
  CLKINVX3 \us13/U81  ( .A(\us13/n14 ), .Y(\us13/n52 ) );
  OAI22XL \us13/U80  ( .A0(\us13/n201 ), .A1(\us13/n52 ), .B0(\us13/n202 ), 
        .B1(\us13/n114 ), .Y(\us13/n193 ) );
  CLKINVX3 \us13/U79  ( .A(sa13[5]), .Y(\us13/n252 ) );
  NOR2X2 \us13/U78  ( .A(\us13/n252 ), .B(\us13/n234 ), .Y(\us13/n55 ) );
  CLKINVX3 \us13/U77  ( .A(sa13[7]), .Y(\us13/n129 ) );
  NOR2X4 \us13/U76  ( .A(\us13/n129 ), .B(\us13/n69 ), .Y(\us13/n24 ) );
  AOI22XL \us13/U75  ( .A0(\us13/n70 ), .A1(\us13/n24 ), .B0(\us13/n96 ), .B1(
        \us13/n129 ), .Y(\us13/n241 ) );
  NOR2X2 \us13/U74  ( .A(\us13/n252 ), .B(sa13[0]), .Y(\us13/n89 ) );
  CLKINVX3 \us13/U73  ( .A(sa13[0]), .Y(\us13/n234 ) );
  NOR2X4 \us13/U72  ( .A(\us13/n69 ), .B(sa13[7]), .Y(\us13/n33 ) );
  INVX12 \us13/U71  ( .A(\us13/n33 ), .Y(\us13/n27 ) );
  CLKINVX3 \us13/U70  ( .A(\us13/n1 ), .Y(\us13/n6 ) );
  CLKINVX3 \us13/U69  ( .A(\us13/n1 ), .Y(\us13/n5 ) );
  INVXL \us13/U68  ( .A(\us13/n24 ), .Y(\us13/n36 ) );
  INVX4 \us13/U67  ( .A(\us13/n3 ), .Y(\us13/n4 ) );
  INVXL \us13/U66  ( .A(\us13/n36 ), .Y(\us13/n3 ) );
  INVX4 \us13/U65  ( .A(sa13[1]), .Y(\us13/n226 ) );
  INVX4 \us13/U64  ( .A(\us13/n43 ), .Y(\us13/n20 ) );
  AOI221X4 \us13/U63  ( .A0(\us13/n24 ), .A1(\us13/n82 ), .B0(\us13/n43 ), 
        .B1(\us13/n295 ), .C0(\us13/n173 ), .Y(\us13/n346 ) );
  AOI221X4 \us13/U62  ( .A0(\us13/n5 ), .A1(\us13/n96 ), .B0(\us13/n43 ), .B1(
        \us13/n239 ), .C0(\us13/n340 ), .Y(\us13/n336 ) );
  AOI222X4 \us13/U61  ( .A0(\us13/n59 ), .A1(\us13/n43 ), .B0(\us13/n6 ), .B1(
        \us13/n221 ), .C0(\us13/n222 ), .C1(\us13/n187 ), .Y(\us13/n218 ) );
  AOI222X4 \us13/U60  ( .A0(\us13/n123 ), .A1(\us13/n43 ), .B0(sa13[2]), .B1(
        \us13/n203 ), .C0(\us13/n6 ), .C1(\us13/n71 ), .Y(\us13/n202 ) );
  AOI221X4 \us13/U59  ( .A0(\us13/n314 ), .A1(\us13/n43 ), .B0(\us13/n160 ), 
        .B1(\us13/n24 ), .C0(\us13/n315 ), .Y(\us13/n307 ) );
  AOI221X4 \us13/U58  ( .A0(\us13/n43 ), .A1(\us13/n208 ), .B0(\us13/n76 ), 
        .B1(\us13/n24 ), .C0(\us13/n209 ), .Y(\us13/n207 ) );
  AOI221X4 \us13/U57  ( .A0(\us13/n43 ), .A1(\us13/n205 ), .B0(\us13/n32 ), 
        .B1(\us13/n6 ), .C0(\us13/n206 ), .Y(\us13/n201 ) );
  AOI221X4 \us13/U56  ( .A0(\us13/n43 ), .A1(\us13/n44 ), .B0(\us13/n45 ), 
        .B1(\us13/n24 ), .C0(\us13/n46 ), .Y(\us13/n9 ) );
  AOI22XL \us13/U55  ( .A0(\us13/n217 ), .A1(\us13/n43 ), .B0(\us13/n33 ), 
        .B1(\us13/n47 ), .Y(\us13/n216 ) );
  AOI22XL \us13/U54  ( .A0(\us13/n98 ), .A1(\us13/n43 ), .B0(\us13/n6 ), .B1(
        \us13/n99 ), .Y(\us13/n97 ) );
  AOI22XL \us13/U53  ( .A0(\us13/n82 ), .A1(\us13/n43 ), .B0(\us13/n83 ), .B1(
        \us13/n24 ), .Y(\us13/n81 ) );
  AOI2BB2XL \us13/U52  ( .B0(\us13/n43 ), .B1(\us13/n94 ), .A0N(\us13/n120 ), 
        .A1N(\us13/n4 ), .Y(\us13/n119 ) );
  AOI222X4 \us13/U51  ( .A0(\us13/n125 ), .A1(\us13/n33 ), .B0(\us13/n145 ), 
        .B1(\us13/n40 ), .C0(\us13/n43 ), .C1(\us13/n184 ), .Y(\us13/n183 ) );
  AOI22XL \us13/U50  ( .A0(\us13/n43 ), .A1(\us13/n303 ), .B0(\us13/n24 ), 
        .B1(\us13/n96 ), .Y(\us13/n358 ) );
  AOI22XL \us13/U49  ( .A0(\us13/n43 ), .A1(\us13/n100 ), .B0(\us13/n24 ), 
        .B1(\us13/n125 ), .Y(\us13/n124 ) );
  AOI21XL \us13/U48  ( .A0(\us13/n159 ), .A1(\us13/n43 ), .B0(\us13/n40 ), .Y(
        \us13/n262 ) );
  AOI22XL \us13/U47  ( .A0(\us13/n40 ), .A1(\us13/n94 ), .B0(\us13/n43 ), .B1(
        \us13/n187 ), .Y(\us13/n244 ) );
  AOI22XL \us13/U46  ( .A0(\us13/n184 ), .A1(\us13/n5 ), .B0(\us13/n198 ), 
        .B1(\us13/n43 ), .Y(\us13/n197 ) );
  NOR2XL \us13/U45  ( .A(\us13/n33 ), .B(\us13/n2 ), .Y(\us13/n302 ) );
  MXI2XL \us13/U44  ( .A(\us13/n2 ), .B(\us13/n6 ), .S0(\us13/n28 ), .Y(
        \us13/n311 ) );
  INVXL \us13/U43  ( .A(\us13/n20 ), .Y(\us13/n2 ) );
  INVX4 \us13/U42  ( .A(\us13/n6 ), .Y(\us13/n18 ) );
  AOI21XL \us13/U41  ( .A0(\us13/n18 ), .A1(\us13/n162 ), .B0(\us13/n25 ), .Y(
        \us13/n161 ) );
  INVX4 \us13/U40  ( .A(sa13[2]), .Y(\us13/n69 ) );
  NOR2X4 \us13/U39  ( .A(\us13/n226 ), .B(\us13/n4 ), .Y(\us13/n40 ) );
  CLKINVX3 \us13/U38  ( .A(sa13[3]), .Y(\us13/n136 ) );
  NOR2X2 \us13/U37  ( .A(\us13/n136 ), .B(sa13[4]), .Y(\us13/n145 ) );
  CLKINVX3 \us13/U36  ( .A(sa13[4]), .Y(\us13/n58 ) );
  NOR2X2 \us13/U35  ( .A(\us13/n58 ), .B(sa13[3]), .Y(\us13/n159 ) );
  NOR2X2 \us13/U34  ( .A(\us13/n136 ), .B(\us13/n58 ), .Y(\us13/n259 ) );
  NOR2X2 \us13/U33  ( .A(sa13[4]), .B(sa13[3]), .Y(\us13/n278 ) );
  NOR2X2 \us13/U32  ( .A(\us13/n259 ), .B(\us13/n278 ), .Y(\us13/n47 ) );
  CLKINVX3 \us13/U31  ( .A(\us13/n259 ), .Y(\us13/n44 ) );
  NOR2X2 \us13/U30  ( .A(\us13/n44 ), .B(sa13[1]), .Y(\us13/n137 ) );
  AOI21XL \us13/U29  ( .A0(\us13/n44 ), .A1(\us13/n111 ), .B0(\us13/n4 ), .Y(
        \us13/n177 ) );
  AOI22XL \us13/U28  ( .A0(\us13/n23 ), .A1(\us13/n24 ), .B0(\us13/n25 ), .B1(
        sa13[2]), .Y(\us13/n22 ) );
  AOI22XL \us13/U27  ( .A0(\us13/n33 ), .A1(sa13[3]), .B0(\us13/n24 ), .B1(
        \us13/n58 ), .Y(\us13/n277 ) );
  NAND2XL \us13/U26  ( .A(\us13/n198 ), .B(\us13/n24 ), .Y(\us13/n132 ) );
  OAI2BB2XL \us13/U25  ( .B0(\us13/n20 ), .B1(\us13/n111 ), .A0N(\us13/n125 ), 
        .A1N(\us13/n24 ), .Y(\us13/n220 ) );
  NAND2XL \us13/U24  ( .A(\us13/n111 ), .B(\us13/n101 ), .Y(\us13/n21 ) );
  NAND2XL \us13/U23  ( .A(\us13/n111 ), .B(\us13/n300 ), .Y(\us13/n187 ) );
  NAND2XL \us13/U22  ( .A(\us13/n111 ), .B(\us13/n121 ), .Y(\us13/n303 ) );
  AOI221XL \us13/U21  ( .A0(\us13/n43 ), .A1(\us13/n151 ), .B0(\us13/n25 ), 
        .B1(\us13/n69 ), .C0(\us13/n275 ), .Y(\us13/n274 ) );
  NOR2BXL \us13/U20  ( .AN(\us13/n101 ), .B(\us13/n25 ), .Y(\us13/n172 ) );
  NAND2X2 \us13/U19  ( .A(\us13/n58 ), .B(\us13/n226 ), .Y(\us13/n34 ) );
  OAI222X1 \us13/U18  ( .A0(\us13/n27 ), .A1(\us13/n34 ), .B0(\us13/n69 ), 
        .B1(\us13/n205 ), .C0(\us13/n20 ), .C1(\us13/n79 ), .Y(\us13/n260 ) );
  OAI222X1 \us13/U17  ( .A0(\us13/n20 ), .A1(\us13/n99 ), .B0(\us13/n27 ), 
        .B1(\us13/n101 ), .C0(\us13/n184 ), .C1(\us13/n4 ), .Y(\us13/n250 ) );
  OAI222X1 \us13/U16  ( .A0(\us13/n4 ), .A1(\us13/n37 ), .B0(\us13/n38 ), .B1(
        \us13/n20 ), .C0(sa13[4]), .C1(\us13/n39 ), .Y(\us13/n35 ) );
  AOI221X1 \us13/U15  ( .A0(\us13/n5 ), .A1(\us13/n19 ), .B0(\us13/n33 ), .B1(
        \us13/n34 ), .C0(\us13/n35 ), .Y(\us13/n11 ) );
  OR2X2 \us13/U14  ( .A(sa13[2]), .B(sa13[7]), .Y(\us13/n1 ) );
  AOI221XL \us13/U13  ( .A0(\us13/n70 ), .A1(\us13/n43 ), .B0(\us13/n24 ), 
        .B1(\us13/n71 ), .C0(\us13/n72 ), .Y(\us13/n53 ) );
  AOI221XL \us13/U12  ( .A0(\us13/n59 ), .A1(\us13/n33 ), .B0(\us13/n43 ), 
        .B1(\us13/n126 ), .C0(\us13/n127 ), .Y(\us13/n113 ) );
  AOI222XL \us13/U11  ( .A0(\us13/n185 ), .A1(\us13/n43 ), .B0(\us13/n186 ), 
        .B1(\us13/n187 ), .C0(\us13/n6 ), .C1(\us13/n188 ), .Y(\us13/n164 ) );
  AOI221X1 \us13/U10  ( .A0(\us13/n313 ), .A1(\us13/n5 ), .B0(\us13/n23 ), 
        .B1(\us13/n2 ), .C0(\us13/n328 ), .Y(\us13/n320 ) );
  AOI221X1 \us13/U9  ( .A0(\us13/n40 ), .A1(\us13/n136 ), .B0(\us13/n33 ), 
        .B1(\us13/n178 ), .C0(\us13/n338 ), .Y(\us13/n337 ) );
  AOI222XL \us13/U8  ( .A0(\us13/n278 ), .A1(\us13/n24 ), .B0(\us13/n42 ), 
        .B1(\us13/n33 ), .C0(\us13/n43 ), .C1(\us13/n136 ), .Y(\us13/n351 ) );
  AOI31X1 \us13/U7  ( .A0(sa13[2]), .A1(\us13/n58 ), .A2(sa13[1]), .B0(
        \us13/n40 ), .Y(\us13/n350 ) );
  AOI31X1 \us13/U6  ( .A0(\us13/n44 ), .A1(\us13/n129 ), .A2(\us13/n130 ), 
        .B0(\us13/n131 ), .Y(\us13/n128 ) );
  AOI221X1 \us13/U5  ( .A0(\us13/n40 ), .A1(\us13/n136 ), .B0(\us13/n33 ), 
        .B1(\us13/n47 ), .C0(\us13/n156 ), .Y(\us13/n141 ) );
  OAI32X1 \us13/U4  ( .A0(\us13/n18 ), .A1(sa13[1]), .A2(\us13/n159 ), .B0(
        sa13[4]), .B1(\us13/n182 ), .Y(\us13/n318 ) );
  OAI32X1 \us13/U3  ( .A0(\us13/n210 ), .A1(\us13/n145 ), .A2(\us13/n18 ), 
        .B0(\us13/n27 ), .B1(\us13/n211 ), .Y(\us13/n209 ) );
  AOI221X1 \us13/U2  ( .A0(\us13/n278 ), .A1(\us13/n40 ), .B0(\us13/n185 ), 
        .B1(\us13/n2 ), .C0(\us13/n279 ), .Y(\us13/n273 ) );
  AOI31XL \us13/U1  ( .A0(\us13/n79 ), .A1(\us13/n44 ), .A2(\us13/n2 ), .B0(
        \us13/n280 ), .Y(\us13/n339 ) );
  NAND2X1 \us20/U366  ( .A(\us20/n47 ), .B(\us20/n226 ), .Y(\us20/n189 ) );
  NOR2X1 \us20/U365  ( .A(\us20/n226 ), .B(sa20[3]), .Y(\us20/n242 ) );
  INVX1 \us20/U364  ( .A(\us20/n242 ), .Y(\us20/n205 ) );
  AND2X1 \us20/U363  ( .A(\us20/n189 ), .B(\us20/n205 ), .Y(\us20/n65 ) );
  NOR2X1 \us20/U362  ( .A(\us20/n226 ), .B(\us20/n47 ), .Y(\us20/n45 ) );
  NOR2X1 \us20/U361  ( .A(\us20/n259 ), .B(\us20/n45 ), .Y(\us20/n73 ) );
  NAND2BX1 \us20/U360  ( .AN(\us20/n73 ), .B(\us20/n6 ), .Y(\us20/n158 ) );
  NOR2X1 \us20/U359  ( .A(\us20/n226 ), .B(\us20/n159 ), .Y(\us20/n95 ) );
  INVX1 \us20/U358  ( .A(\us20/n95 ), .Y(\us20/n111 ) );
  NOR2X1 \us20/U357  ( .A(\us20/n145 ), .B(sa20[1]), .Y(\us20/n42 ) );
  INVX1 \us20/U356  ( .A(\us20/n42 ), .Y(\us20/n121 ) );
  INVX1 \us20/U355  ( .A(\us20/n47 ), .Y(\us20/n96 ) );
  OAI211X1 \us20/U354  ( .A0(\us20/n65 ), .A1(\us20/n27 ), .B0(\us20/n158 ), 
        .C0(\us20/n358 ), .Y(\us20/n355 ) );
  NOR2X1 \us20/U353  ( .A(\us20/n226 ), .B(\us20/n145 ), .Y(\us20/n59 ) );
  NOR2X1 \us20/U352  ( .A(\us20/n96 ), .B(\us20/n59 ), .Y(\us20/n271 ) );
  NOR2X1 \us20/U351  ( .A(\us20/n226 ), .B(\us20/n278 ), .Y(\us20/n217 ) );
  INVX1 \us20/U350  ( .A(\us20/n217 ), .Y(\us20/n150 ) );
  NAND2X1 \us20/U349  ( .A(\us20/n44 ), .B(\us20/n150 ), .Y(\us20/n147 ) );
  NAND2X1 \us20/U348  ( .A(sa20[4]), .B(\us20/n226 ), .Y(\us20/n101 ) );
  INVX1 \us20/U347  ( .A(\us20/n159 ), .Y(\us20/n188 ) );
  NOR2X1 \us20/U346  ( .A(\us20/n188 ), .B(\us20/n226 ), .Y(\us20/n25 ) );
  INVX1 \us20/U345  ( .A(\us20/n172 ), .Y(\us20/n107 ) );
  AOI22X1 \us20/U344  ( .A0(\us20/n33 ), .A1(\us20/n147 ), .B0(\us20/n24 ), 
        .B1(\us20/n107 ), .Y(\us20/n357 ) );
  OAI221XL \us20/U343  ( .A0(\us20/n18 ), .A1(\us20/n121 ), .B0(\us20/n271 ), 
        .B1(\us20/n20 ), .C0(\us20/n357 ), .Y(\us20/n356 ) );
  MXI2X1 \us20/U342  ( .A(\us20/n355 ), .B(\us20/n356 ), .S0(\us20/n252 ), .Y(
        \us20/n331 ) );
  INVX1 \us20/U341  ( .A(\us20/n59 ), .Y(\us20/n79 ) );
  AND2X1 \us20/U340  ( .A(\us20/n101 ), .B(\us20/n79 ), .Y(\us20/n325 ) );
  XNOR2X1 \us20/U339  ( .A(sa20[5]), .B(\us20/n226 ), .Y(\us20/n352 ) );
  NOR2X1 \us20/U338  ( .A(\us20/n226 ), .B(\us20/n136 ), .Y(\us20/n281 ) );
  INVX1 \us20/U337  ( .A(\us20/n281 ), .Y(\us20/n19 ) );
  NAND2X1 \us20/U336  ( .A(\us20/n145 ), .B(\us20/n226 ), .Y(\us20/n223 ) );
  AOI21X1 \us20/U335  ( .A0(\us20/n19 ), .A1(\us20/n223 ), .B0(\us20/n27 ), 
        .Y(\us20/n354 ) );
  AOI31X1 \us20/U334  ( .A0(\us20/n6 ), .A1(\us20/n352 ), .A2(\us20/n259 ), 
        .B0(\us20/n354 ), .Y(\us20/n353 ) );
  OAI221XL \us20/U333  ( .A0(\us20/n20 ), .A1(\us20/n34 ), .B0(\us20/n325 ), 
        .B1(\us20/n4 ), .C0(\us20/n353 ), .Y(\us20/n347 ) );
  INVX1 \us20/U332  ( .A(\us20/n352 ), .Y(\us20/n349 ) );
  NAND2X1 \us20/U331  ( .A(\us20/n278 ), .B(\us20/n6 ), .Y(\us20/n74 ) );
  OAI211X1 \us20/U330  ( .A0(\us20/n349 ), .A1(\us20/n74 ), .B0(\us20/n350 ), 
        .C0(\us20/n351 ), .Y(\us20/n348 ) );
  MXI2X1 \us20/U329  ( .A(\us20/n347 ), .B(\us20/n348 ), .S0(\us20/n252 ), .Y(
        \us20/n332 ) );
  NOR2X1 \us20/U328  ( .A(\us20/n44 ), .B(\us20/n226 ), .Y(\us20/n157 ) );
  INVX1 \us20/U327  ( .A(\us20/n157 ), .Y(\us20/n240 ) );
  NAND2X1 \us20/U326  ( .A(\us20/n240 ), .B(\us20/n189 ), .Y(\us20/n68 ) );
  NOR2X1 \us20/U325  ( .A(\us20/n20 ), .B(\us20/n159 ), .Y(\us20/n225 ) );
  NOR2X1 \us20/U324  ( .A(\us20/n225 ), .B(\us20/n40 ), .Y(\us20/n345 ) );
  INVX1 \us20/U323  ( .A(\us20/n278 ), .Y(\us20/n94 ) );
  NAND2X1 \us20/U322  ( .A(\us20/n94 ), .B(\us20/n226 ), .Y(\us20/n199 ) );
  NAND2X1 \us20/U321  ( .A(\us20/n199 ), .B(\us20/n205 ), .Y(\us20/n82 ) );
  NAND2X1 \us20/U320  ( .A(\us20/n19 ), .B(\us20/n199 ), .Y(\us20/n295 ) );
  NOR2X1 \us20/U319  ( .A(\us20/n226 ), .B(\us20/n259 ), .Y(\us20/n210 ) );
  NOR2X1 \us20/U318  ( .A(\us20/n27 ), .B(\us20/n210 ), .Y(\us20/n173 ) );
  MXI2X1 \us20/U317  ( .A(\us20/n345 ), .B(\us20/n346 ), .S0(\us20/n252 ), .Y(
        \us20/n342 ) );
  NOR2X1 \us20/U316  ( .A(sa20[1]), .B(sa20[3]), .Y(\us20/n163 ) );
  INVX1 \us20/U315  ( .A(\us20/n163 ), .Y(\us20/n37 ) );
  INVX1 \us20/U314  ( .A(\us20/n173 ), .Y(\us20/n344 ) );
  AOI21X1 \us20/U313  ( .A0(\us20/n240 ), .A1(\us20/n37 ), .B0(\us20/n344 ), 
        .Y(\us20/n343 ) );
  AOI211X1 \us20/U312  ( .A0(\us20/n5 ), .A1(\us20/n68 ), .B0(\us20/n342 ), 
        .C0(\us20/n343 ), .Y(\us20/n333 ) );
  NOR2X1 \us20/U311  ( .A(\us20/n18 ), .B(\us20/n226 ), .Y(\us20/n258 ) );
  NAND2X1 \us20/U310  ( .A(\us20/n278 ), .B(sa20[1]), .Y(\us20/n204 ) );
  NOR2X1 \us20/U309  ( .A(\us20/n188 ), .B(sa20[1]), .Y(\us20/n179 ) );
  INVX1 \us20/U308  ( .A(\us20/n179 ), .Y(\us20/n330 ) );
  NAND2X1 \us20/U307  ( .A(\us20/n204 ), .B(\us20/n330 ), .Y(\us20/n239 ) );
  NOR2X1 \us20/U306  ( .A(\us20/n136 ), .B(sa20[1]), .Y(\us20/n299 ) );
  NOR2X1 \us20/U305  ( .A(\us20/n299 ), .B(\us20/n210 ), .Y(\us20/n341 ) );
  OAI32X1 \us20/U304  ( .A0(\us20/n27 ), .A1(\us20/n278 ), .A2(\us20/n95 ), 
        .B0(\us20/n341 ), .B1(\us20/n4 ), .Y(\us20/n340 ) );
  INVX1 \us20/U303  ( .A(\us20/n45 ), .Y(\us20/n126 ) );
  NAND2X1 \us20/U302  ( .A(\us20/n126 ), .B(\us20/n101 ), .Y(\us20/n178 ) );
  NOR2X1 \us20/U301  ( .A(\us20/n18 ), .B(\us20/n136 ), .Y(\us20/n280 ) );
  OAI21XL \us20/U300  ( .A0(\us20/n4 ), .A1(\us20/n121 ), .B0(\us20/n339 ), 
        .Y(\us20/n338 ) );
  MXI2X1 \us20/U299  ( .A(\us20/n336 ), .B(\us20/n337 ), .S0(\us20/n252 ), .Y(
        \us20/n335 ) );
  NOR2X1 \us20/U298  ( .A(\us20/n258 ), .B(\us20/n335 ), .Y(\us20/n334 ) );
  MX4X1 \us20/U297  ( .A(\us20/n331 ), .B(\us20/n332 ), .C(\us20/n333 ), .D(
        \us20/n334 ), .S0(sa20[6]), .S1(\us20/n234 ), .Y(sa22_sr[0]) );
  INVX1 \us20/U296  ( .A(\us20/n299 ), .Y(\us20/n80 ) );
  NOR2X1 \us20/U295  ( .A(\us20/n111 ), .B(\us20/n18 ), .Y(\us20/n269 ) );
  INVX1 \us20/U294  ( .A(\us20/n269 ), .Y(\us20/n75 ) );
  OAI221XL \us20/U293  ( .A0(\us20/n18 ), .A1(\us20/n330 ), .B0(\us20/n20 ), 
        .B1(\us20/n80 ), .C0(\us20/n75 ), .Y(\us20/n329 ) );
  AOI221X1 \us20/U292  ( .A0(\us20/n325 ), .A1(\us20/n33 ), .B0(\us20/n24 ), 
        .B1(\us20/n303 ), .C0(\us20/n329 ), .Y(\us20/n319 ) );
  NOR2X1 \us20/U291  ( .A(\us20/n234 ), .B(sa20[5]), .Y(\us20/n14 ) );
  NOR2X1 \us20/U290  ( .A(\us20/n25 ), .B(\us20/n299 ), .Y(\us20/n313 ) );
  NAND2X1 \us20/U289  ( .A(\us20/n44 ), .B(\us20/n226 ), .Y(\us20/n300 ) );
  AND2X1 \us20/U288  ( .A(\us20/n300 ), .B(\us20/n240 ), .Y(\us20/n23 ) );
  OAI32X1 \us20/U287  ( .A0(\us20/n4 ), .A1(\us20/n145 ), .A2(\us20/n210 ), 
        .B0(\us20/n137 ), .B1(\us20/n27 ), .Y(\us20/n328 ) );
  NOR2X1 \us20/U286  ( .A(sa20[0]), .B(sa20[5]), .Y(\us20/n16 ) );
  INVX1 \us20/U285  ( .A(\us20/n16 ), .Y(\us20/n114 ) );
  INVX1 \us20/U284  ( .A(\us20/n145 ), .Y(\us20/n149 ) );
  NOR2X1 \us20/U283  ( .A(\us20/n47 ), .B(sa20[1]), .Y(\us20/n98 ) );
  INVX1 \us20/U282  ( .A(\us20/n98 ), .Y(\us20/n284 ) );
  OAI21XL \us20/U281  ( .A0(\us20/n69 ), .A1(\us20/n284 ), .B0(\us20/n27 ), 
        .Y(\us20/n327 ) );
  AOI31X1 \us20/U280  ( .A0(\us20/n111 ), .A1(\us20/n149 ), .A2(\us20/n327 ), 
        .B0(\us20/n225 ), .Y(\us20/n326 ) );
  OAI21XL \us20/U279  ( .A0(\us20/n325 ), .A1(\us20/n18 ), .B0(\us20/n326 ), 
        .Y(\us20/n322 ) );
  NAND2X1 \us20/U278  ( .A(\us20/n19 ), .B(\us20/n189 ), .Y(\us20/n71 ) );
  NOR2X1 \us20/U277  ( .A(\us20/n71 ), .B(\us20/n18 ), .Y(\us20/n135 ) );
  AOI21X1 \us20/U276  ( .A0(\us20/n40 ), .A1(sa20[4]), .B0(\us20/n135 ), .Y(
        \us20/n324 ) );
  OAI221XL \us20/U275  ( .A0(\us20/n47 ), .A1(\us20/n27 ), .B0(\us20/n65 ), 
        .B1(\us20/n20 ), .C0(\us20/n324 ), .Y(\us20/n323 ) );
  AOI22X1 \us20/U274  ( .A0(\us20/n55 ), .A1(\us20/n322 ), .B0(\us20/n89 ), 
        .B1(\us20/n323 ), .Y(\us20/n321 ) );
  OAI221XL \us20/U273  ( .A0(\us20/n319 ), .A1(\us20/n52 ), .B0(\us20/n320 ), 
        .B1(\us20/n114 ), .C0(\us20/n321 ), .Y(\us20/n304 ) );
  NOR2X1 \us20/U272  ( .A(\us20/n226 ), .B(\us20/n58 ), .Y(\us20/n290 ) );
  INVX1 \us20/U271  ( .A(\us20/n290 ), .Y(\us20/n200 ) );
  NAND2X1 \us20/U270  ( .A(\us20/n34 ), .B(\us20/n200 ), .Y(\us20/n120 ) );
  INVX1 \us20/U269  ( .A(\us20/n210 ), .Y(\us20/n100 ) );
  OAI221XL \us20/U268  ( .A0(\us20/n20 ), .A1(\us20/n100 ), .B0(sa20[3]), .B1(
        \us20/n4 ), .C0(\us20/n262 ), .Y(\us20/n317 ) );
  INVX1 \us20/U267  ( .A(\us20/n258 ), .Y(\us20/n182 ) );
  AOI211X1 \us20/U266  ( .A0(\us20/n33 ), .A1(\us20/n120 ), .B0(\us20/n317 ), 
        .C0(\us20/n318 ), .Y(\us20/n306 ) );
  NAND2X1 \us20/U265  ( .A(\us20/n100 ), .B(\us20/n199 ), .Y(\us20/n151 ) );
  INVX1 \us20/U264  ( .A(\us20/n151 ), .Y(\us20/n314 ) );
  NOR2X1 \us20/U263  ( .A(\us20/n45 ), .B(\us20/n163 ), .Y(\us20/n160 ) );
  INVX1 \us20/U262  ( .A(\us20/n295 ), .Y(\us20/n92 ) );
  AOI21X1 \us20/U261  ( .A0(sa20[1]), .A1(\us20/n58 ), .B0(\us20/n98 ), .Y(
        \us20/n316 ) );
  OAI22X1 \us20/U260  ( .A0(\us20/n92 ), .A1(\us20/n18 ), .B0(\us20/n316 ), 
        .B1(\us20/n27 ), .Y(\us20/n315 ) );
  NOR2X1 \us20/U259  ( .A(\us20/n149 ), .B(\us20/n226 ), .Y(\us20/n41 ) );
  INVX1 \us20/U258  ( .A(\us20/n41 ), .Y(\us20/n105 ) );
  NAND2X1 \us20/U257  ( .A(\us20/n284 ), .B(\us20/n105 ), .Y(\us20/n227 ) );
  AOI21X1 \us20/U256  ( .A0(\us20/n313 ), .A1(\us20/n33 ), .B0(\us20/n269 ), 
        .Y(\us20/n312 ) );
  OAI221XL \us20/U255  ( .A0(\us20/n149 ), .A1(\us20/n20 ), .B0(\us20/n4 ), 
        .B1(\us20/n227 ), .C0(\us20/n312 ), .Y(\us20/n309 ) );
  AOI21X1 \us20/U254  ( .A0(\us20/n226 ), .A1(\us20/n188 ), .B0(\us20/n242 ), 
        .Y(\us20/n185 ) );
  INVX1 \us20/U253  ( .A(\us20/n185 ), .Y(\us20/n48 ) );
  AND2X1 \us20/U252  ( .A(\us20/n223 ), .B(\us20/n240 ), .Y(\us20/n28 ) );
  OAI221XL \us20/U251  ( .A0(\us20/n27 ), .A1(\us20/n44 ), .B0(\us20/n4 ), 
        .B1(\us20/n48 ), .C0(\us20/n311 ), .Y(\us20/n310 ) );
  AOI22X1 \us20/U250  ( .A0(\us20/n89 ), .A1(\us20/n309 ), .B0(\us20/n55 ), 
        .B1(\us20/n310 ), .Y(\us20/n308 ) );
  OAI221XL \us20/U249  ( .A0(\us20/n306 ), .A1(\us20/n52 ), .B0(\us20/n307 ), 
        .B1(\us20/n114 ), .C0(\us20/n308 ), .Y(\us20/n305 ) );
  MX2X1 \us20/U248  ( .A(\us20/n304 ), .B(\us20/n305 ), .S0(sa20[6]), .Y(
        sa22_sr[1]) );
  INVX1 \us20/U247  ( .A(\us20/n187 ), .Y(\us20/n61 ) );
  MXI2X1 \us20/U246  ( .A(\us20/n303 ), .B(\us20/n61 ), .S0(\us20/n69 ), .Y(
        \us20/n301 ) );
  MXI2X1 \us20/U245  ( .A(\us20/n301 ), .B(\us20/n147 ), .S0(\us20/n302 ), .Y(
        \us20/n285 ) );
  NAND2X1 \us20/U244  ( .A(\us20/n200 ), .B(\us20/n300 ), .Y(\us20/n99 ) );
  INVX1 \us20/U243  ( .A(\us20/n99 ), .Y(\us20/n296 ) );
  NOR2X1 \us20/U242  ( .A(\us20/n299 ), .B(\us20/n242 ), .Y(\us20/n298 ) );
  NAND2X1 \us20/U241  ( .A(sa20[1]), .B(\us20/n47 ), .Y(\us20/n122 ) );
  NOR2X1 \us20/U240  ( .A(\us20/n159 ), .B(\us20/n217 ), .Y(\us20/n198 ) );
  OAI221XL \us20/U239  ( .A0(\us20/n298 ), .A1(\us20/n27 ), .B0(\us20/n20 ), 
        .B1(\us20/n122 ), .C0(\us20/n132 ), .Y(\us20/n297 ) );
  AOI221X1 \us20/U238  ( .A0(\us20/n225 ), .A1(\us20/n226 ), .B0(\us20/n296 ), 
        .B1(\us20/n6 ), .C0(\us20/n297 ), .Y(\us20/n291 ) );
  OAI2BB2X1 \us20/U237  ( .B0(\us20/n27 ), .B1(\us20/n295 ), .A0N(\us20/n34 ), 
        .A1N(\us20/n24 ), .Y(\us20/n293 ) );
  AOI21X1 \us20/U236  ( .A0(\us20/n101 ), .A1(\us20/n150 ), .B0(\us20/n20 ), 
        .Y(\us20/n294 ) );
  AOI211X1 \us20/U235  ( .A0(\us20/n5 ), .A1(\us20/n79 ), .B0(\us20/n293 ), 
        .C0(\us20/n294 ), .Y(\us20/n292 ) );
  INVX1 \us20/U234  ( .A(\us20/n89 ), .Y(\us20/n10 ) );
  OAI22X1 \us20/U233  ( .A0(\us20/n291 ), .A1(\us20/n114 ), .B0(\us20/n292 ), 
        .B1(\us20/n10 ), .Y(\us20/n286 ) );
  INVX1 \us20/U232  ( .A(\us20/n225 ), .Y(\us20/n288 ) );
  NAND2X1 \us20/U231  ( .A(\us20/n200 ), .B(\us20/n284 ), .Y(\us20/n102 ) );
  NOR2X1 \us20/U230  ( .A(\us20/n290 ), .B(\us20/n163 ), .Y(\us20/n184 ) );
  AOI22X1 \us20/U229  ( .A0(\us20/n102 ), .A1(\us20/n69 ), .B0(\us20/n184 ), 
        .B1(\us20/n33 ), .Y(\us20/n289 ) );
  AOI31X1 \us20/U228  ( .A0(\us20/n132 ), .A1(\us20/n288 ), .A2(\us20/n289 ), 
        .B0(\us20/n52 ), .Y(\us20/n287 ) );
  AOI211X1 \us20/U227  ( .A0(\us20/n285 ), .A1(\us20/n55 ), .B0(\us20/n286 ), 
        .C0(\us20/n287 ), .Y(\us20/n263 ) );
  NAND2X1 \us20/U226  ( .A(\us20/n284 ), .B(\us20/n122 ), .Y(\us20/n125 ) );
  NOR2X1 \us20/U225  ( .A(\us20/n199 ), .B(\us20/n4 ), .Y(\us20/n50 ) );
  AOI21X1 \us20/U224  ( .A0(\us20/n200 ), .A1(\us20/n223 ), .B0(\us20/n20 ), 
        .Y(\us20/n283 ) );
  AOI211X1 \us20/U223  ( .A0(\us20/n5 ), .A1(\us20/n125 ), .B0(\us20/n50 ), 
        .C0(\us20/n283 ), .Y(\us20/n282 ) );
  OAI221XL \us20/U222  ( .A0(\us20/n281 ), .A1(\us20/n27 ), .B0(\us20/n4 ), 
        .B1(\us20/n111 ), .C0(\us20/n282 ), .Y(\us20/n265 ) );
  INVX1 \us20/U221  ( .A(\us20/n280 ), .Y(\us20/n247 ) );
  NAND2X1 \us20/U220  ( .A(\us20/n41 ), .B(\us20/n33 ), .Y(\us20/n272 ) );
  OAI221XL \us20/U219  ( .A0(sa20[1]), .A1(\us20/n247 ), .B0(\us20/n4 ), .B1(
        \us20/n189 ), .C0(\us20/n272 ), .Y(\us20/n279 ) );
  NAND2X1 \us20/U218  ( .A(sa20[2]), .B(\us20/n149 ), .Y(\us20/n276 ) );
  XNOR2X1 \us20/U217  ( .A(\us20/n129 ), .B(sa20[1]), .Y(\us20/n155 ) );
  MXI2X1 \us20/U216  ( .A(\us20/n276 ), .B(\us20/n277 ), .S0(\us20/n155 ), .Y(
        \us20/n275 ) );
  OAI22X1 \us20/U215  ( .A0(\us20/n273 ), .A1(\us20/n10 ), .B0(\us20/n274 ), 
        .B1(\us20/n52 ), .Y(\us20/n266 ) );
  NOR2X1 \us20/U214  ( .A(\us20/n20 ), .B(\us20/n226 ), .Y(\us20/n176 ) );
  OAI21XL \us20/U213  ( .A0(\us20/n4 ), .A1(\us20/n271 ), .B0(\us20/n272 ), 
        .Y(\us20/n270 ) );
  OAI31X1 \us20/U212  ( .A0(\us20/n176 ), .A1(\us20/n269 ), .A2(\us20/n270 ), 
        .B0(\us20/n16 ), .Y(\us20/n268 ) );
  INVX1 \us20/U211  ( .A(\us20/n268 ), .Y(\us20/n267 ) );
  AOI211X1 \us20/U210  ( .A0(\us20/n55 ), .A1(\us20/n265 ), .B0(\us20/n266 ), 
        .C0(\us20/n267 ), .Y(\us20/n264 ) );
  MXI2X1 \us20/U209  ( .A(\us20/n263 ), .B(\us20/n264 ), .S0(sa20[6]), .Y(
        sa22_sr[2]) );
  NOR2X1 \us20/U208  ( .A(\us20/n94 ), .B(sa20[1]), .Y(\us20/n211 ) );
  INVX1 \us20/U207  ( .A(\us20/n262 ), .Y(\us20/n261 ) );
  AOI211X1 \us20/U206  ( .A0(\us20/n259 ), .A1(\us20/n24 ), .B0(\us20/n260 ), 
        .C0(\us20/n261 ), .Y(\us20/n255 ) );
  OAI22X1 \us20/U205  ( .A0(\us20/n20 ), .A1(\us20/n68 ), .B0(\us20/n27 ), 
        .B1(\us20/n37 ), .Y(\us20/n257 ) );
  NOR3X1 \us20/U204  ( .A(\us20/n257 ), .B(\us20/n258 ), .C(\us20/n50 ), .Y(
        \us20/n256 ) );
  MXI2X1 \us20/U203  ( .A(\us20/n255 ), .B(\us20/n256 ), .S0(\us20/n252 ), .Y(
        \us20/n254 ) );
  AOI221X1 \us20/U202  ( .A0(\us20/n211 ), .A1(\us20/n5 ), .B0(\us20/n40 ), 
        .B1(sa20[4]), .C0(\us20/n254 ), .Y(\us20/n248 ) );
  INVX1 \us20/U201  ( .A(\us20/n211 ), .Y(\us20/n106 ) );
  NAND2X1 \us20/U200  ( .A(\us20/n200 ), .B(\us20/n106 ), .Y(\us20/n83 ) );
  NAND2X1 \us20/U199  ( .A(\us20/n199 ), .B(\us20/n204 ), .Y(\us20/n169 ) );
  AOI2BB2X1 \us20/U198  ( .B0(\us20/n65 ), .B1(\us20/n24 ), .A0N(\us20/n169 ), 
        .A1N(\us20/n20 ), .Y(\us20/n253 ) );
  OAI221XL \us20/U197  ( .A0(\us20/n172 ), .A1(\us20/n18 ), .B0(\us20/n27 ), 
        .B1(\us20/n83 ), .C0(\us20/n253 ), .Y(\us20/n251 ) );
  MXI2X1 \us20/U196  ( .A(\us20/n250 ), .B(\us20/n251 ), .S0(\us20/n252 ), .Y(
        \us20/n249 ) );
  MXI2X1 \us20/U195  ( .A(\us20/n248 ), .B(\us20/n249 ), .S0(\us20/n234 ), .Y(
        \us20/n228 ) );
  OAI21XL \us20/U194  ( .A0(\us20/n58 ), .A1(\us20/n27 ), .B0(\us20/n247 ), 
        .Y(\us20/n245 ) );
  NOR2X1 \us20/U193  ( .A(sa20[7]), .B(\us20/n145 ), .Y(\us20/n246 ) );
  XNOR2X1 \us20/U192  ( .A(\us20/n69 ), .B(sa20[1]), .Y(\us20/n130 ) );
  MXI2X1 \us20/U191  ( .A(\us20/n245 ), .B(\us20/n246 ), .S0(\us20/n130 ), .Y(
        \us20/n243 ) );
  OAI211X1 \us20/U190  ( .A0(\us20/n4 ), .A1(\us20/n149 ), .B0(\us20/n243 ), 
        .C0(\us20/n244 ), .Y(\us20/n230 ) );
  NOR2X1 \us20/U189  ( .A(\us20/n242 ), .B(\us20/n137 ), .Y(\us20/n70 ) );
  OAI221XL \us20/U188  ( .A0(\us20/n159 ), .A1(\us20/n27 ), .B0(\us20/n20 ), 
        .B1(\us20/n34 ), .C0(\us20/n241 ), .Y(\us20/n231 ) );
  NAND2X1 \us20/U187  ( .A(\us20/n101 ), .B(\us20/n240 ), .Y(\us20/n76 ) );
  AOI21X1 \us20/U186  ( .A0(\us20/n122 ), .A1(\us20/n106 ), .B0(\us20/n129 ), 
        .Y(\us20/n237 ) );
  INVX1 \us20/U185  ( .A(\us20/n239 ), .Y(\us20/n238 ) );
  OAI21XL \us20/U184  ( .A0(\us20/n237 ), .A1(\us20/n43 ), .B0(\us20/n238 ), 
        .Y(\us20/n236 ) );
  OAI221XL \us20/U183  ( .A0(\us20/n18 ), .A1(\us20/n76 ), .B0(\us20/n59 ), 
        .B1(\us20/n27 ), .C0(\us20/n236 ), .Y(\us20/n232 ) );
  AOI2BB2X1 \us20/U182  ( .B0(\us20/n24 ), .B1(\us20/n187 ), .A0N(\us20/n227 ), 
        .A1N(\us20/n20 ), .Y(\us20/n235 ) );
  OAI211X1 \us20/U181  ( .A0(\us20/n27 ), .A1(\us20/n122 ), .B0(\us20/n158 ), 
        .C0(\us20/n235 ), .Y(\us20/n233 ) );
  MX4X1 \us20/U180  ( .A(\us20/n230 ), .B(\us20/n231 ), .C(\us20/n232 ), .D(
        \us20/n233 ), .S0(\us20/n234 ), .S1(sa20[5]), .Y(\us20/n229 ) );
  MX2X1 \us20/U179  ( .A(\us20/n228 ), .B(\us20/n229 ), .S0(sa20[6]), .Y(
        sa22_sr[3]) );
  NOR2BX1 \us20/U178  ( .AN(\us20/n204 ), .B(\us20/n137 ), .Y(\us20/n110 ) );
  INVX1 \us20/U177  ( .A(\us20/n110 ), .Y(\us20/n64 ) );
  AOI22X1 \us20/U176  ( .A0(\us20/n225 ), .A1(\us20/n226 ), .B0(\us20/n6 ), 
        .B1(\us20/n227 ), .Y(\us20/n224 ) );
  OAI221XL \us20/U175  ( .A0(\us20/n27 ), .A1(\us20/n64 ), .B0(\us20/n4 ), 
        .B1(\us20/n83 ), .C0(\us20/n224 ), .Y(\us20/n212 ) );
  NAND2X1 \us20/U174  ( .A(\us20/n34 ), .B(\us20/n204 ), .Y(\us20/n221 ) );
  OAI21XL \us20/U173  ( .A0(\us20/n69 ), .A1(\us20/n223 ), .B0(\us20/n27 ), 
        .Y(\us20/n222 ) );
  NOR2X1 \us20/U172  ( .A(\us20/n217 ), .B(\us20/n42 ), .Y(\us20/n208 ) );
  AOI211X1 \us20/U171  ( .A0(\us20/n208 ), .A1(\us20/n5 ), .B0(\us20/n220 ), 
        .C0(\us20/n173 ), .Y(\us20/n219 ) );
  OAI22X1 \us20/U170  ( .A0(\us20/n218 ), .A1(\us20/n10 ), .B0(\us20/n219 ), 
        .B1(\us20/n114 ), .Y(\us20/n213 ) );
  INVX1 \us20/U169  ( .A(\us20/n135 ), .Y(\us20/n215 ) );
  NOR2X1 \us20/U168  ( .A(\us20/n4 ), .B(\us20/n159 ), .Y(\us20/n31 ) );
  INVX1 \us20/U167  ( .A(\us20/n31 ), .Y(\us20/n196 ) );
  AOI31X1 \us20/U166  ( .A0(\us20/n215 ), .A1(\us20/n196 ), .A2(\us20/n216 ), 
        .B0(\us20/n52 ), .Y(\us20/n214 ) );
  AOI211X1 \us20/U165  ( .A0(\us20/n55 ), .A1(\us20/n212 ), .B0(\us20/n213 ), 
        .C0(\us20/n214 ), .Y(\us20/n190 ) );
  INVX1 \us20/U164  ( .A(\us20/n207 ), .Y(\us20/n192 ) );
  NOR2X1 \us20/U163  ( .A(\us20/n25 ), .B(\us20/n98 ), .Y(\us20/n32 ) );
  OAI22X1 \us20/U162  ( .A0(\us20/n28 ), .A1(\us20/n4 ), .B0(\us20/n188 ), 
        .B1(\us20/n27 ), .Y(\us20/n206 ) );
  NAND2X1 \us20/U161  ( .A(\us20/n204 ), .B(\us20/n80 ), .Y(\us20/n118 ) );
  INVX1 \us20/U160  ( .A(\us20/n118 ), .Y(\us20/n123 ) );
  NAND2X1 \us20/U159  ( .A(\us20/n94 ), .B(\us20/n79 ), .Y(\us20/n203 ) );
  OAI2BB1X1 \us20/U158  ( .A0N(\us20/n199 ), .A1N(\us20/n200 ), .B0(\us20/n33 ), .Y(\us20/n195 ) );
  INVX1 \us20/U157  ( .A(\us20/n55 ), .Y(\us20/n12 ) );
  AOI31X1 \us20/U156  ( .A0(\us20/n195 ), .A1(\us20/n196 ), .A2(\us20/n197 ), 
        .B0(\us20/n12 ), .Y(\us20/n194 ) );
  AOI211X1 \us20/U155  ( .A0(\us20/n89 ), .A1(\us20/n192 ), .B0(\us20/n193 ), 
        .C0(\us20/n194 ), .Y(\us20/n191 ) );
  MXI2X1 \us20/U154  ( .A(\us20/n190 ), .B(\us20/n191 ), .S0(sa20[6]), .Y(
        sa22_sr[4]) );
  OAI21XL \us20/U153  ( .A0(\us20/n69 ), .A1(\us20/n189 ), .B0(\us20/n27 ), 
        .Y(\us20/n186 ) );
  INVX1 \us20/U152  ( .A(\us20/n183 ), .Y(\us20/n180 ) );
  NAND2X1 \us20/U151  ( .A(\us20/n74 ), .B(\us20/n182 ), .Y(\us20/n181 ) );
  AOI211X1 \us20/U150  ( .A0(\us20/n179 ), .A1(\us20/n24 ), .B0(\us20/n180 ), 
        .C0(\us20/n181 ), .Y(\us20/n165 ) );
  INVX1 \us20/U149  ( .A(\us20/n178 ), .Y(\us20/n175 ) );
  AOI211X1 \us20/U148  ( .A0(\us20/n175 ), .A1(\us20/n5 ), .B0(\us20/n176 ), 
        .C0(\us20/n177 ), .Y(\us20/n174 ) );
  OAI221XL \us20/U147  ( .A0(\us20/n159 ), .A1(\us20/n27 ), .B0(\us20/n145 ), 
        .B1(\us20/n20 ), .C0(\us20/n174 ), .Y(\us20/n167 ) );
  MXI2X1 \us20/U146  ( .A(\us20/n40 ), .B(\us20/n173 ), .S0(\us20/n96 ), .Y(
        \us20/n170 ) );
  AOI22X1 \us20/U145  ( .A0(\us20/n137 ), .A1(\us20/n24 ), .B0(\us20/n172 ), 
        .B1(\us20/n6 ), .Y(\us20/n171 ) );
  OAI211X1 \us20/U144  ( .A0(\us20/n20 ), .A1(\us20/n169 ), .B0(\us20/n170 ), 
        .C0(\us20/n171 ), .Y(\us20/n168 ) );
  AOI22X1 \us20/U143  ( .A0(\us20/n89 ), .A1(\us20/n167 ), .B0(\us20/n55 ), 
        .B1(\us20/n168 ), .Y(\us20/n166 ) );
  OAI221XL \us20/U142  ( .A0(\us20/n164 ), .A1(\us20/n114 ), .B0(\us20/n165 ), 
        .B1(\us20/n52 ), .C0(\us20/n166 ), .Y(\us20/n138 ) );
  OAI21XL \us20/U141  ( .A0(\us20/n41 ), .A1(\us20/n163 ), .B0(\us20/n69 ), 
        .Y(\us20/n162 ) );
  AOI221X1 \us20/U140  ( .A0(\us20/n159 ), .A1(\us20/n24 ), .B0(\us20/n160 ), 
        .B1(\us20/n33 ), .C0(\us20/n161 ), .Y(\us20/n140 ) );
  OAI21XL \us20/U139  ( .A0(\us20/n157 ), .A1(\us20/n20 ), .B0(\us20/n158 ), 
        .Y(\us20/n156 ) );
  NOR2X1 \us20/U138  ( .A(\us20/n4 ), .B(\us20/n136 ), .Y(\us20/n153 ) );
  NOR2X1 \us20/U137  ( .A(\us20/n145 ), .B(\us20/n69 ), .Y(\us20/n154 ) );
  MXI2X1 \us20/U136  ( .A(\us20/n153 ), .B(\us20/n154 ), .S0(\us20/n155 ), .Y(
        \us20/n152 ) );
  OAI221XL \us20/U135  ( .A0(\us20/n110 ), .A1(\us20/n18 ), .B0(\us20/n20 ), 
        .B1(\us20/n151 ), .C0(\us20/n152 ), .Y(\us20/n143 ) );
  AOI21X1 \us20/U134  ( .A0(\us20/n149 ), .A1(\us20/n150 ), .B0(\us20/n18 ), 
        .Y(\us20/n148 ) );
  AOI2BB1X1 \us20/U133  ( .A0N(\us20/n147 ), .A1N(\us20/n27 ), .B0(\us20/n148 ), .Y(\us20/n146 ) );
  OAI221XL \us20/U132  ( .A0(\us20/n145 ), .A1(\us20/n20 ), .B0(\us20/n4 ), 
        .B1(\us20/n34 ), .C0(\us20/n146 ), .Y(\us20/n144 ) );
  AOI22X1 \us20/U131  ( .A0(\us20/n89 ), .A1(\us20/n143 ), .B0(\us20/n14 ), 
        .B1(\us20/n144 ), .Y(\us20/n142 ) );
  OAI221XL \us20/U130  ( .A0(\us20/n140 ), .A1(\us20/n12 ), .B0(\us20/n141 ), 
        .B1(\us20/n114 ), .C0(\us20/n142 ), .Y(\us20/n139 ) );
  MX2X1 \us20/U129  ( .A(\us20/n138 ), .B(\us20/n139 ), .S0(sa20[6]), .Y(
        sa22_sr[5]) );
  INVX1 \us20/U128  ( .A(\us20/n70 ), .Y(\us20/n133 ) );
  OAI22X1 \us20/U127  ( .A0(\us20/n4 ), .A1(\us20/n136 ), .B0(\us20/n137 ), 
        .B1(\us20/n27 ), .Y(\us20/n134 ) );
  AOI211X1 \us20/U126  ( .A0(\us20/n133 ), .A1(\us20/n69 ), .B0(\us20/n134 ), 
        .C0(\us20/n135 ), .Y(\us20/n112 ) );
  INVX1 \us20/U125  ( .A(\us20/n132 ), .Y(\us20/n131 ) );
  OAI21XL \us20/U124  ( .A0(\us20/n18 ), .A1(\us20/n37 ), .B0(\us20/n128 ), 
        .Y(\us20/n127 ) );
  OAI221XL \us20/U123  ( .A0(\us20/n18 ), .A1(\us20/n105 ), .B0(\us20/n123 ), 
        .B1(\us20/n27 ), .C0(\us20/n124 ), .Y(\us20/n116 ) );
  NAND2X1 \us20/U122  ( .A(\us20/n121 ), .B(\us20/n122 ), .Y(\us20/n30 ) );
  OAI221XL \us20/U121  ( .A0(\us20/n18 ), .A1(\us20/n118 ), .B0(\us20/n27 ), 
        .B1(\us20/n30 ), .C0(\us20/n119 ), .Y(\us20/n117 ) );
  AOI22X1 \us20/U120  ( .A0(\us20/n89 ), .A1(\us20/n116 ), .B0(\us20/n55 ), 
        .B1(\us20/n117 ), .Y(\us20/n115 ) );
  OAI221XL \us20/U119  ( .A0(\us20/n112 ), .A1(\us20/n52 ), .B0(\us20/n113 ), 
        .B1(\us20/n114 ), .C0(\us20/n115 ), .Y(\us20/n84 ) );
  OAI22X1 \us20/U118  ( .A0(\us20/n110 ), .A1(\us20/n4 ), .B0(\us20/n20 ), 
        .B1(\us20/n21 ), .Y(\us20/n108 ) );
  AOI21X1 \us20/U117  ( .A0(sa20[1]), .A1(\us20/n58 ), .B0(\us20/n27 ), .Y(
        \us20/n109 ) );
  AOI211X1 \us20/U116  ( .A0(\us20/n5 ), .A1(\us20/n107 ), .B0(\us20/n108 ), 
        .C0(\us20/n109 ), .Y(\us20/n86 ) );
  OAI22X1 \us20/U115  ( .A0(\us20/n45 ), .A1(\us20/n4 ), .B0(sa20[4]), .B1(
        \us20/n18 ), .Y(\us20/n103 ) );
  AOI21X1 \us20/U114  ( .A0(\us20/n105 ), .A1(\us20/n106 ), .B0(\us20/n20 ), 
        .Y(\us20/n104 ) );
  AOI211X1 \us20/U113  ( .A0(\us20/n33 ), .A1(\us20/n102 ), .B0(\us20/n103 ), 
        .C0(\us20/n104 ), .Y(\us20/n87 ) );
  NAND2X1 \us20/U112  ( .A(\us20/n100 ), .B(\us20/n101 ), .Y(\us20/n62 ) );
  OAI221XL \us20/U111  ( .A0(\us20/n27 ), .A1(\us20/n62 ), .B0(\us20/n4 ), 
        .B1(\us20/n21 ), .C0(\us20/n97 ), .Y(\us20/n90 ) );
  NOR3X1 \us20/U110  ( .A(\us20/n4 ), .B(\us20/n95 ), .C(\us20/n96 ), .Y(
        \us20/n67 ) );
  AOI31X1 \us20/U109  ( .A0(\us20/n79 ), .A1(\us20/n94 ), .A2(\us20/n6 ), .B0(
        \us20/n67 ), .Y(\us20/n93 ) );
  OAI221XL \us20/U108  ( .A0(\us20/n73 ), .A1(\us20/n27 ), .B0(\us20/n92 ), 
        .B1(\us20/n20 ), .C0(\us20/n93 ), .Y(\us20/n91 ) );
  AOI22X1 \us20/U107  ( .A0(\us20/n89 ), .A1(\us20/n90 ), .B0(\us20/n16 ), 
        .B1(\us20/n91 ), .Y(\us20/n88 ) );
  OAI221XL \us20/U106  ( .A0(\us20/n86 ), .A1(\us20/n52 ), .B0(\us20/n87 ), 
        .B1(\us20/n12 ), .C0(\us20/n88 ), .Y(\us20/n85 ) );
  MX2X1 \us20/U105  ( .A(\us20/n84 ), .B(\us20/n85 ), .S0(sa20[6]), .Y(
        sa22_sr[6]) );
  INVX1 \us20/U104  ( .A(\us20/n81 ), .Y(\us20/n77 ) );
  AOI21X1 \us20/U103  ( .A0(\us20/n79 ), .A1(\us20/n80 ), .B0(\us20/n27 ), .Y(
        \us20/n78 ) );
  AOI211X1 \us20/U102  ( .A0(\us20/n5 ), .A1(\us20/n76 ), .B0(\us20/n77 ), 
        .C0(\us20/n78 ), .Y(\us20/n51 ) );
  OAI211X1 \us20/U101  ( .A0(\us20/n73 ), .A1(\us20/n27 ), .B0(\us20/n74 ), 
        .C0(\us20/n75 ), .Y(\us20/n72 ) );
  AOI21X1 \us20/U100  ( .A0(\us20/n68 ), .A1(\us20/n69 ), .B0(\us20/n6 ), .Y(
        \us20/n63 ) );
  INVX1 \us20/U99  ( .A(\us20/n67 ), .Y(\us20/n66 ) );
  OAI221XL \us20/U98  ( .A0(\us20/n63 ), .A1(\us20/n64 ), .B0(\us20/n65 ), 
        .B1(\us20/n27 ), .C0(\us20/n66 ), .Y(\us20/n56 ) );
  AOI2BB2X1 \us20/U97  ( .B0(\us20/n61 ), .B1(\us20/n24 ), .A0N(\us20/n62 ), 
        .A1N(\us20/n20 ), .Y(\us20/n60 ) );
  OAI221XL \us20/U96  ( .A0(\us20/n58 ), .A1(\us20/n18 ), .B0(\us20/n59 ), 
        .B1(\us20/n27 ), .C0(\us20/n60 ), .Y(\us20/n57 ) );
  AOI22X1 \us20/U95  ( .A0(\us20/n55 ), .A1(\us20/n56 ), .B0(\us20/n16 ), .B1(
        \us20/n57 ), .Y(\us20/n54 ) );
  OAI221XL \us20/U94  ( .A0(\us20/n51 ), .A1(\us20/n52 ), .B0(\us20/n53 ), 
        .B1(\us20/n10 ), .C0(\us20/n54 ), .Y(\us20/n7 ) );
  INVX1 \us20/U93  ( .A(\us20/n50 ), .Y(\us20/n49 ) );
  OAI221XL \us20/U92  ( .A0(\us20/n47 ), .A1(\us20/n18 ), .B0(\us20/n27 ), 
        .B1(\us20/n48 ), .C0(\us20/n49 ), .Y(\us20/n46 ) );
  NOR2X1 \us20/U91  ( .A(\us20/n41 ), .B(\us20/n42 ), .Y(\us20/n38 ) );
  INVX1 \us20/U90  ( .A(\us20/n40 ), .Y(\us20/n39 ) );
  INVX1 \us20/U89  ( .A(\us20/n32 ), .Y(\us20/n26 ) );
  AOI21X1 \us20/U88  ( .A0(\us20/n5 ), .A1(\us20/n30 ), .B0(\us20/n31 ), .Y(
        \us20/n29 ) );
  OAI221XL \us20/U87  ( .A0(\us20/n26 ), .A1(\us20/n27 ), .B0(\us20/n28 ), 
        .B1(\us20/n20 ), .C0(\us20/n29 ), .Y(\us20/n15 ) );
  OAI221XL \us20/U86  ( .A0(\us20/n18 ), .A1(\us20/n19 ), .B0(\us20/n20 ), 
        .B1(\us20/n21 ), .C0(\us20/n22 ), .Y(\us20/n17 ) );
  AOI22X1 \us20/U85  ( .A0(\us20/n14 ), .A1(\us20/n15 ), .B0(\us20/n16 ), .B1(
        \us20/n17 ), .Y(\us20/n13 ) );
  OAI221XL \us20/U84  ( .A0(\us20/n9 ), .A1(\us20/n10 ), .B0(\us20/n11 ), .B1(
        \us20/n12 ), .C0(\us20/n13 ), .Y(\us20/n8 ) );
  MX2X1 \us20/U83  ( .A(\us20/n7 ), .B(\us20/n8 ), .S0(sa20[6]), .Y(sa22_sr[7]) );
  NOR2X4 \us20/U82  ( .A(\us20/n129 ), .B(sa20[2]), .Y(\us20/n43 ) );
  CLKINVX3 \us20/U81  ( .A(\us20/n14 ), .Y(\us20/n52 ) );
  OAI22XL \us20/U80  ( .A0(\us20/n201 ), .A1(\us20/n52 ), .B0(\us20/n202 ), 
        .B1(\us20/n114 ), .Y(\us20/n193 ) );
  CLKINVX3 \us20/U79  ( .A(sa20[5]), .Y(\us20/n252 ) );
  NOR2X2 \us20/U78  ( .A(\us20/n252 ), .B(\us20/n234 ), .Y(\us20/n55 ) );
  CLKINVX3 \us20/U77  ( .A(sa20[7]), .Y(\us20/n129 ) );
  NOR2X4 \us20/U76  ( .A(\us20/n129 ), .B(\us20/n69 ), .Y(\us20/n24 ) );
  AOI22XL \us20/U75  ( .A0(\us20/n70 ), .A1(\us20/n24 ), .B0(\us20/n96 ), .B1(
        \us20/n129 ), .Y(\us20/n241 ) );
  NOR2X2 \us20/U74  ( .A(\us20/n252 ), .B(sa20[0]), .Y(\us20/n89 ) );
  CLKINVX3 \us20/U73  ( .A(sa20[0]), .Y(\us20/n234 ) );
  NOR2X4 \us20/U72  ( .A(\us20/n69 ), .B(sa20[7]), .Y(\us20/n33 ) );
  INVX12 \us20/U71  ( .A(\us20/n33 ), .Y(\us20/n27 ) );
  CLKINVX3 \us20/U70  ( .A(\us20/n1 ), .Y(\us20/n6 ) );
  CLKINVX3 \us20/U69  ( .A(\us20/n1 ), .Y(\us20/n5 ) );
  INVXL \us20/U68  ( .A(\us20/n24 ), .Y(\us20/n36 ) );
  INVX4 \us20/U67  ( .A(\us20/n3 ), .Y(\us20/n4 ) );
  INVXL \us20/U66  ( .A(\us20/n36 ), .Y(\us20/n3 ) );
  INVX4 \us20/U65  ( .A(sa20[1]), .Y(\us20/n226 ) );
  INVX4 \us20/U64  ( .A(\us20/n43 ), .Y(\us20/n20 ) );
  AOI221X4 \us20/U63  ( .A0(\us20/n24 ), .A1(\us20/n82 ), .B0(\us20/n43 ), 
        .B1(\us20/n295 ), .C0(\us20/n173 ), .Y(\us20/n346 ) );
  AOI221X4 \us20/U62  ( .A0(\us20/n5 ), .A1(\us20/n96 ), .B0(\us20/n43 ), .B1(
        \us20/n239 ), .C0(\us20/n340 ), .Y(\us20/n336 ) );
  AOI222X4 \us20/U61  ( .A0(\us20/n59 ), .A1(\us20/n43 ), .B0(\us20/n6 ), .B1(
        \us20/n221 ), .C0(\us20/n222 ), .C1(\us20/n187 ), .Y(\us20/n218 ) );
  AOI222X4 \us20/U60  ( .A0(\us20/n123 ), .A1(\us20/n43 ), .B0(sa20[2]), .B1(
        \us20/n203 ), .C0(\us20/n6 ), .C1(\us20/n71 ), .Y(\us20/n202 ) );
  AOI221X4 \us20/U59  ( .A0(\us20/n314 ), .A1(\us20/n43 ), .B0(\us20/n160 ), 
        .B1(\us20/n24 ), .C0(\us20/n315 ), .Y(\us20/n307 ) );
  AOI221X4 \us20/U58  ( .A0(\us20/n43 ), .A1(\us20/n208 ), .B0(\us20/n76 ), 
        .B1(\us20/n24 ), .C0(\us20/n209 ), .Y(\us20/n207 ) );
  AOI221X4 \us20/U57  ( .A0(\us20/n43 ), .A1(\us20/n205 ), .B0(\us20/n32 ), 
        .B1(\us20/n6 ), .C0(\us20/n206 ), .Y(\us20/n201 ) );
  AOI221X4 \us20/U56  ( .A0(\us20/n43 ), .A1(\us20/n44 ), .B0(\us20/n45 ), 
        .B1(\us20/n24 ), .C0(\us20/n46 ), .Y(\us20/n9 ) );
  AOI22XL \us20/U55  ( .A0(\us20/n217 ), .A1(\us20/n43 ), .B0(\us20/n33 ), 
        .B1(\us20/n47 ), .Y(\us20/n216 ) );
  AOI22XL \us20/U54  ( .A0(\us20/n98 ), .A1(\us20/n43 ), .B0(\us20/n6 ), .B1(
        \us20/n99 ), .Y(\us20/n97 ) );
  AOI22XL \us20/U53  ( .A0(\us20/n82 ), .A1(\us20/n43 ), .B0(\us20/n83 ), .B1(
        \us20/n24 ), .Y(\us20/n81 ) );
  AOI2BB2XL \us20/U52  ( .B0(\us20/n43 ), .B1(\us20/n94 ), .A0N(\us20/n120 ), 
        .A1N(\us20/n4 ), .Y(\us20/n119 ) );
  AOI222X4 \us20/U51  ( .A0(\us20/n125 ), .A1(\us20/n33 ), .B0(\us20/n145 ), 
        .B1(\us20/n40 ), .C0(\us20/n43 ), .C1(\us20/n184 ), .Y(\us20/n183 ) );
  AOI22XL \us20/U50  ( .A0(\us20/n43 ), .A1(\us20/n303 ), .B0(\us20/n24 ), 
        .B1(\us20/n96 ), .Y(\us20/n358 ) );
  AOI22XL \us20/U49  ( .A0(\us20/n43 ), .A1(\us20/n100 ), .B0(\us20/n24 ), 
        .B1(\us20/n125 ), .Y(\us20/n124 ) );
  AOI21XL \us20/U48  ( .A0(\us20/n159 ), .A1(\us20/n43 ), .B0(\us20/n40 ), .Y(
        \us20/n262 ) );
  AOI22XL \us20/U47  ( .A0(\us20/n40 ), .A1(\us20/n94 ), .B0(\us20/n43 ), .B1(
        \us20/n187 ), .Y(\us20/n244 ) );
  AOI22XL \us20/U46  ( .A0(\us20/n184 ), .A1(\us20/n5 ), .B0(\us20/n198 ), 
        .B1(\us20/n43 ), .Y(\us20/n197 ) );
  NOR2XL \us20/U45  ( .A(\us20/n33 ), .B(\us20/n2 ), .Y(\us20/n302 ) );
  MXI2XL \us20/U44  ( .A(\us20/n2 ), .B(\us20/n6 ), .S0(\us20/n28 ), .Y(
        \us20/n311 ) );
  INVXL \us20/U43  ( .A(\us20/n20 ), .Y(\us20/n2 ) );
  INVX4 \us20/U42  ( .A(\us20/n6 ), .Y(\us20/n18 ) );
  AOI21XL \us20/U41  ( .A0(\us20/n18 ), .A1(\us20/n162 ), .B0(\us20/n25 ), .Y(
        \us20/n161 ) );
  INVX4 \us20/U40  ( .A(sa20[2]), .Y(\us20/n69 ) );
  NOR2X4 \us20/U39  ( .A(\us20/n226 ), .B(\us20/n4 ), .Y(\us20/n40 ) );
  CLKINVX3 \us20/U38  ( .A(sa20[3]), .Y(\us20/n136 ) );
  NOR2X2 \us20/U37  ( .A(\us20/n136 ), .B(sa20[4]), .Y(\us20/n145 ) );
  CLKINVX3 \us20/U36  ( .A(sa20[4]), .Y(\us20/n58 ) );
  NOR2X2 \us20/U35  ( .A(\us20/n58 ), .B(sa20[3]), .Y(\us20/n159 ) );
  NOR2X2 \us20/U34  ( .A(\us20/n136 ), .B(\us20/n58 ), .Y(\us20/n259 ) );
  NOR2X2 \us20/U33  ( .A(sa20[4]), .B(sa20[3]), .Y(\us20/n278 ) );
  NOR2X2 \us20/U32  ( .A(\us20/n259 ), .B(\us20/n278 ), .Y(\us20/n47 ) );
  CLKINVX3 \us20/U31  ( .A(\us20/n259 ), .Y(\us20/n44 ) );
  NOR2X2 \us20/U30  ( .A(\us20/n44 ), .B(sa20[1]), .Y(\us20/n137 ) );
  AOI21XL \us20/U29  ( .A0(\us20/n44 ), .A1(\us20/n111 ), .B0(\us20/n4 ), .Y(
        \us20/n177 ) );
  AOI22XL \us20/U28  ( .A0(\us20/n23 ), .A1(\us20/n24 ), .B0(\us20/n25 ), .B1(
        sa20[2]), .Y(\us20/n22 ) );
  AOI22XL \us20/U27  ( .A0(\us20/n33 ), .A1(sa20[3]), .B0(\us20/n24 ), .B1(
        \us20/n58 ), .Y(\us20/n277 ) );
  NAND2XL \us20/U26  ( .A(\us20/n198 ), .B(\us20/n24 ), .Y(\us20/n132 ) );
  OAI2BB2XL \us20/U25  ( .B0(\us20/n20 ), .B1(\us20/n111 ), .A0N(\us20/n125 ), 
        .A1N(\us20/n24 ), .Y(\us20/n220 ) );
  NAND2XL \us20/U24  ( .A(\us20/n111 ), .B(\us20/n101 ), .Y(\us20/n21 ) );
  NAND2XL \us20/U23  ( .A(\us20/n111 ), .B(\us20/n300 ), .Y(\us20/n187 ) );
  NAND2XL \us20/U22  ( .A(\us20/n111 ), .B(\us20/n121 ), .Y(\us20/n303 ) );
  AOI221XL \us20/U21  ( .A0(\us20/n43 ), .A1(\us20/n151 ), .B0(\us20/n25 ), 
        .B1(\us20/n69 ), .C0(\us20/n275 ), .Y(\us20/n274 ) );
  NOR2BXL \us20/U20  ( .AN(\us20/n101 ), .B(\us20/n25 ), .Y(\us20/n172 ) );
  NAND2X2 \us20/U19  ( .A(\us20/n58 ), .B(\us20/n226 ), .Y(\us20/n34 ) );
  OAI222X1 \us20/U18  ( .A0(\us20/n27 ), .A1(\us20/n34 ), .B0(\us20/n69 ), 
        .B1(\us20/n205 ), .C0(\us20/n20 ), .C1(\us20/n79 ), .Y(\us20/n260 ) );
  OAI222X1 \us20/U17  ( .A0(\us20/n20 ), .A1(\us20/n99 ), .B0(\us20/n27 ), 
        .B1(\us20/n101 ), .C0(\us20/n184 ), .C1(\us20/n4 ), .Y(\us20/n250 ) );
  OAI222X1 \us20/U16  ( .A0(\us20/n4 ), .A1(\us20/n37 ), .B0(\us20/n38 ), .B1(
        \us20/n20 ), .C0(sa20[4]), .C1(\us20/n39 ), .Y(\us20/n35 ) );
  AOI221X1 \us20/U15  ( .A0(\us20/n5 ), .A1(\us20/n19 ), .B0(\us20/n33 ), .B1(
        \us20/n34 ), .C0(\us20/n35 ), .Y(\us20/n11 ) );
  OR2X2 \us20/U14  ( .A(sa20[2]), .B(sa20[7]), .Y(\us20/n1 ) );
  AOI221XL \us20/U13  ( .A0(\us20/n59 ), .A1(\us20/n33 ), .B0(\us20/n43 ), 
        .B1(\us20/n126 ), .C0(\us20/n127 ), .Y(\us20/n113 ) );
  AOI221XL \us20/U12  ( .A0(\us20/n70 ), .A1(\us20/n43 ), .B0(\us20/n24 ), 
        .B1(\us20/n71 ), .C0(\us20/n72 ), .Y(\us20/n53 ) );
  AOI221X1 \us20/U11  ( .A0(\us20/n313 ), .A1(\us20/n5 ), .B0(\us20/n23 ), 
        .B1(\us20/n2 ), .C0(\us20/n328 ), .Y(\us20/n320 ) );
  AOI222XL \us20/U10  ( .A0(\us20/n185 ), .A1(\us20/n43 ), .B0(\us20/n186 ), 
        .B1(\us20/n187 ), .C0(\us20/n6 ), .C1(\us20/n188 ), .Y(\us20/n164 ) );
  AOI221X1 \us20/U9  ( .A0(\us20/n40 ), .A1(\us20/n136 ), .B0(\us20/n33 ), 
        .B1(\us20/n178 ), .C0(\us20/n338 ), .Y(\us20/n337 ) );
  AOI222XL \us20/U8  ( .A0(\us20/n278 ), .A1(\us20/n24 ), .B0(\us20/n42 ), 
        .B1(\us20/n33 ), .C0(\us20/n43 ), .C1(\us20/n136 ), .Y(\us20/n351 ) );
  AOI31X1 \us20/U7  ( .A0(sa20[2]), .A1(\us20/n58 ), .A2(sa20[1]), .B0(
        \us20/n40 ), .Y(\us20/n350 ) );
  AOI31X1 \us20/U6  ( .A0(\us20/n44 ), .A1(\us20/n129 ), .A2(\us20/n130 ), 
        .B0(\us20/n131 ), .Y(\us20/n128 ) );
  AOI221X1 \us20/U5  ( .A0(\us20/n278 ), .A1(\us20/n40 ), .B0(\us20/n185 ), 
        .B1(\us20/n2 ), .C0(\us20/n279 ), .Y(\us20/n273 ) );
  OAI32X1 \us20/U4  ( .A0(\us20/n18 ), .A1(sa20[1]), .A2(\us20/n159 ), .B0(
        sa20[4]), .B1(\us20/n182 ), .Y(\us20/n318 ) );
  AOI221X1 \us20/U3  ( .A0(\us20/n40 ), .A1(\us20/n136 ), .B0(\us20/n33 ), 
        .B1(\us20/n47 ), .C0(\us20/n156 ), .Y(\us20/n141 ) );
  OAI32X1 \us20/U2  ( .A0(\us20/n210 ), .A1(\us20/n145 ), .A2(\us20/n18 ), 
        .B0(\us20/n27 ), .B1(\us20/n211 ), .Y(\us20/n209 ) );
  AOI31XL \us20/U1  ( .A0(\us20/n79 ), .A1(\us20/n44 ), .A2(\us20/n2 ), .B0(
        \us20/n280 ), .Y(\us20/n339 ) );
  NAND2X1 \us21/U366  ( .A(\us21/n47 ), .B(\us21/n226 ), .Y(\us21/n189 ) );
  NOR2X1 \us21/U365  ( .A(\us21/n226 ), .B(sa21[3]), .Y(\us21/n242 ) );
  INVX1 \us21/U364  ( .A(\us21/n242 ), .Y(\us21/n205 ) );
  AND2X1 \us21/U363  ( .A(\us21/n189 ), .B(\us21/n205 ), .Y(\us21/n65 ) );
  NOR2X1 \us21/U362  ( .A(\us21/n226 ), .B(\us21/n47 ), .Y(\us21/n45 ) );
  NOR2X1 \us21/U361  ( .A(\us21/n259 ), .B(\us21/n45 ), .Y(\us21/n73 ) );
  NAND2BX1 \us21/U360  ( .AN(\us21/n73 ), .B(\us21/n6 ), .Y(\us21/n158 ) );
  NOR2X1 \us21/U359  ( .A(\us21/n226 ), .B(\us21/n159 ), .Y(\us21/n95 ) );
  INVX1 \us21/U358  ( .A(\us21/n95 ), .Y(\us21/n111 ) );
  NOR2X1 \us21/U357  ( .A(\us21/n145 ), .B(sa21[1]), .Y(\us21/n42 ) );
  INVX1 \us21/U356  ( .A(\us21/n42 ), .Y(\us21/n121 ) );
  INVX1 \us21/U355  ( .A(\us21/n47 ), .Y(\us21/n96 ) );
  OAI211X1 \us21/U354  ( .A0(\us21/n65 ), .A1(\us21/n27 ), .B0(\us21/n158 ), 
        .C0(\us21/n358 ), .Y(\us21/n355 ) );
  NOR2X1 \us21/U353  ( .A(\us21/n226 ), .B(\us21/n145 ), .Y(\us21/n59 ) );
  NOR2X1 \us21/U352  ( .A(\us21/n96 ), .B(\us21/n59 ), .Y(\us21/n271 ) );
  NOR2X1 \us21/U351  ( .A(\us21/n226 ), .B(\us21/n278 ), .Y(\us21/n217 ) );
  INVX1 \us21/U350  ( .A(\us21/n217 ), .Y(\us21/n150 ) );
  NAND2X1 \us21/U349  ( .A(\us21/n44 ), .B(\us21/n150 ), .Y(\us21/n147 ) );
  NAND2X1 \us21/U348  ( .A(sa21[4]), .B(\us21/n226 ), .Y(\us21/n101 ) );
  INVX1 \us21/U347  ( .A(\us21/n159 ), .Y(\us21/n188 ) );
  NOR2X1 \us21/U346  ( .A(\us21/n188 ), .B(\us21/n226 ), .Y(\us21/n25 ) );
  INVX1 \us21/U345  ( .A(\us21/n172 ), .Y(\us21/n107 ) );
  AOI22X1 \us21/U344  ( .A0(\us21/n33 ), .A1(\us21/n147 ), .B0(\us21/n24 ), 
        .B1(\us21/n107 ), .Y(\us21/n357 ) );
  OAI221XL \us21/U343  ( .A0(\us21/n18 ), .A1(\us21/n121 ), .B0(\us21/n271 ), 
        .B1(\us21/n20 ), .C0(\us21/n357 ), .Y(\us21/n356 ) );
  MXI2X1 \us21/U342  ( .A(\us21/n355 ), .B(\us21/n356 ), .S0(\us21/n252 ), .Y(
        \us21/n331 ) );
  INVX1 \us21/U341  ( .A(\us21/n59 ), .Y(\us21/n79 ) );
  AND2X1 \us21/U340  ( .A(\us21/n101 ), .B(\us21/n79 ), .Y(\us21/n325 ) );
  XNOR2X1 \us21/U339  ( .A(sa21[5]), .B(\us21/n226 ), .Y(\us21/n352 ) );
  NOR2X1 \us21/U338  ( .A(\us21/n226 ), .B(\us21/n136 ), .Y(\us21/n281 ) );
  INVX1 \us21/U337  ( .A(\us21/n281 ), .Y(\us21/n19 ) );
  NAND2X1 \us21/U336  ( .A(\us21/n145 ), .B(\us21/n226 ), .Y(\us21/n223 ) );
  AOI21X1 \us21/U335  ( .A0(\us21/n19 ), .A1(\us21/n223 ), .B0(\us21/n27 ), 
        .Y(\us21/n354 ) );
  AOI31X1 \us21/U334  ( .A0(\us21/n6 ), .A1(\us21/n352 ), .A2(\us21/n259 ), 
        .B0(\us21/n354 ), .Y(\us21/n353 ) );
  OAI221XL \us21/U333  ( .A0(\us21/n20 ), .A1(\us21/n34 ), .B0(\us21/n325 ), 
        .B1(\us21/n4 ), .C0(\us21/n353 ), .Y(\us21/n347 ) );
  INVX1 \us21/U332  ( .A(\us21/n352 ), .Y(\us21/n349 ) );
  NAND2X1 \us21/U331  ( .A(\us21/n278 ), .B(\us21/n6 ), .Y(\us21/n74 ) );
  OAI211X1 \us21/U330  ( .A0(\us21/n349 ), .A1(\us21/n74 ), .B0(\us21/n350 ), 
        .C0(\us21/n351 ), .Y(\us21/n348 ) );
  MXI2X1 \us21/U329  ( .A(\us21/n347 ), .B(\us21/n348 ), .S0(\us21/n252 ), .Y(
        \us21/n332 ) );
  NOR2X1 \us21/U328  ( .A(\us21/n44 ), .B(\us21/n226 ), .Y(\us21/n157 ) );
  INVX1 \us21/U327  ( .A(\us21/n157 ), .Y(\us21/n240 ) );
  NAND2X1 \us21/U326  ( .A(\us21/n240 ), .B(\us21/n189 ), .Y(\us21/n68 ) );
  NOR2X1 \us21/U325  ( .A(\us21/n20 ), .B(\us21/n159 ), .Y(\us21/n225 ) );
  NOR2X1 \us21/U324  ( .A(\us21/n225 ), .B(\us21/n40 ), .Y(\us21/n345 ) );
  INVX1 \us21/U323  ( .A(\us21/n278 ), .Y(\us21/n94 ) );
  NAND2X1 \us21/U322  ( .A(\us21/n94 ), .B(\us21/n226 ), .Y(\us21/n199 ) );
  NAND2X1 \us21/U321  ( .A(\us21/n199 ), .B(\us21/n205 ), .Y(\us21/n82 ) );
  NAND2X1 \us21/U320  ( .A(\us21/n19 ), .B(\us21/n199 ), .Y(\us21/n295 ) );
  NOR2X1 \us21/U319  ( .A(\us21/n226 ), .B(\us21/n259 ), .Y(\us21/n210 ) );
  NOR2X1 \us21/U318  ( .A(\us21/n27 ), .B(\us21/n210 ), .Y(\us21/n173 ) );
  MXI2X1 \us21/U317  ( .A(\us21/n345 ), .B(\us21/n346 ), .S0(\us21/n252 ), .Y(
        \us21/n342 ) );
  NOR2X1 \us21/U316  ( .A(sa21[1]), .B(sa21[3]), .Y(\us21/n163 ) );
  INVX1 \us21/U315  ( .A(\us21/n163 ), .Y(\us21/n37 ) );
  INVX1 \us21/U314  ( .A(\us21/n173 ), .Y(\us21/n344 ) );
  AOI21X1 \us21/U313  ( .A0(\us21/n240 ), .A1(\us21/n37 ), .B0(\us21/n344 ), 
        .Y(\us21/n343 ) );
  AOI211X1 \us21/U312  ( .A0(\us21/n5 ), .A1(\us21/n68 ), .B0(\us21/n342 ), 
        .C0(\us21/n343 ), .Y(\us21/n333 ) );
  NOR2X1 \us21/U311  ( .A(\us21/n18 ), .B(\us21/n226 ), .Y(\us21/n258 ) );
  NAND2X1 \us21/U310  ( .A(\us21/n278 ), .B(sa21[1]), .Y(\us21/n204 ) );
  NOR2X1 \us21/U309  ( .A(\us21/n188 ), .B(sa21[1]), .Y(\us21/n179 ) );
  INVX1 \us21/U308  ( .A(\us21/n179 ), .Y(\us21/n330 ) );
  NAND2X1 \us21/U307  ( .A(\us21/n204 ), .B(\us21/n330 ), .Y(\us21/n239 ) );
  NOR2X1 \us21/U306  ( .A(\us21/n136 ), .B(sa21[1]), .Y(\us21/n299 ) );
  NOR2X1 \us21/U305  ( .A(\us21/n299 ), .B(\us21/n210 ), .Y(\us21/n341 ) );
  OAI32X1 \us21/U304  ( .A0(\us21/n27 ), .A1(\us21/n278 ), .A2(\us21/n95 ), 
        .B0(\us21/n341 ), .B1(\us21/n4 ), .Y(\us21/n340 ) );
  INVX1 \us21/U303  ( .A(\us21/n45 ), .Y(\us21/n126 ) );
  NAND2X1 \us21/U302  ( .A(\us21/n126 ), .B(\us21/n101 ), .Y(\us21/n178 ) );
  NOR2X1 \us21/U301  ( .A(\us21/n18 ), .B(\us21/n136 ), .Y(\us21/n280 ) );
  OAI21XL \us21/U300  ( .A0(\us21/n4 ), .A1(\us21/n121 ), .B0(\us21/n339 ), 
        .Y(\us21/n338 ) );
  MXI2X1 \us21/U299  ( .A(\us21/n336 ), .B(\us21/n337 ), .S0(\us21/n252 ), .Y(
        \us21/n335 ) );
  NOR2X1 \us21/U298  ( .A(\us21/n258 ), .B(\us21/n335 ), .Y(\us21/n334 ) );
  MX4X1 \us21/U297  ( .A(\us21/n331 ), .B(\us21/n332 ), .C(\us21/n333 ), .D(
        \us21/n334 ), .S0(sa21[6]), .S1(\us21/n234 ), .Y(sa23_sr[0]) );
  INVX1 \us21/U296  ( .A(\us21/n299 ), .Y(\us21/n80 ) );
  NOR2X1 \us21/U295  ( .A(\us21/n111 ), .B(\us21/n18 ), .Y(\us21/n269 ) );
  INVX1 \us21/U294  ( .A(\us21/n269 ), .Y(\us21/n75 ) );
  OAI221XL \us21/U293  ( .A0(\us21/n18 ), .A1(\us21/n330 ), .B0(\us21/n20 ), 
        .B1(\us21/n80 ), .C0(\us21/n75 ), .Y(\us21/n329 ) );
  AOI221X1 \us21/U292  ( .A0(\us21/n325 ), .A1(\us21/n33 ), .B0(\us21/n24 ), 
        .B1(\us21/n303 ), .C0(\us21/n329 ), .Y(\us21/n319 ) );
  NOR2X1 \us21/U291  ( .A(\us21/n234 ), .B(sa21[5]), .Y(\us21/n14 ) );
  NOR2X1 \us21/U290  ( .A(\us21/n25 ), .B(\us21/n299 ), .Y(\us21/n313 ) );
  NAND2X1 \us21/U289  ( .A(\us21/n44 ), .B(\us21/n226 ), .Y(\us21/n300 ) );
  AND2X1 \us21/U288  ( .A(\us21/n300 ), .B(\us21/n240 ), .Y(\us21/n23 ) );
  OAI32X1 \us21/U287  ( .A0(\us21/n4 ), .A1(\us21/n145 ), .A2(\us21/n210 ), 
        .B0(\us21/n137 ), .B1(\us21/n27 ), .Y(\us21/n328 ) );
  NOR2X1 \us21/U286  ( .A(sa21[0]), .B(sa21[5]), .Y(\us21/n16 ) );
  INVX1 \us21/U285  ( .A(\us21/n16 ), .Y(\us21/n114 ) );
  INVX1 \us21/U284  ( .A(\us21/n145 ), .Y(\us21/n149 ) );
  NOR2X1 \us21/U283  ( .A(\us21/n47 ), .B(sa21[1]), .Y(\us21/n98 ) );
  INVX1 \us21/U282  ( .A(\us21/n98 ), .Y(\us21/n284 ) );
  OAI21XL \us21/U281  ( .A0(\us21/n69 ), .A1(\us21/n284 ), .B0(\us21/n27 ), 
        .Y(\us21/n327 ) );
  AOI31X1 \us21/U280  ( .A0(\us21/n111 ), .A1(\us21/n149 ), .A2(\us21/n327 ), 
        .B0(\us21/n225 ), .Y(\us21/n326 ) );
  OAI21XL \us21/U279  ( .A0(\us21/n325 ), .A1(\us21/n18 ), .B0(\us21/n326 ), 
        .Y(\us21/n322 ) );
  NAND2X1 \us21/U278  ( .A(\us21/n19 ), .B(\us21/n189 ), .Y(\us21/n71 ) );
  NOR2X1 \us21/U277  ( .A(\us21/n71 ), .B(\us21/n18 ), .Y(\us21/n135 ) );
  AOI21X1 \us21/U276  ( .A0(\us21/n40 ), .A1(sa21[4]), .B0(\us21/n135 ), .Y(
        \us21/n324 ) );
  OAI221XL \us21/U275  ( .A0(\us21/n47 ), .A1(\us21/n27 ), .B0(\us21/n65 ), 
        .B1(\us21/n20 ), .C0(\us21/n324 ), .Y(\us21/n323 ) );
  AOI22X1 \us21/U274  ( .A0(\us21/n55 ), .A1(\us21/n322 ), .B0(\us21/n89 ), 
        .B1(\us21/n323 ), .Y(\us21/n321 ) );
  OAI221XL \us21/U273  ( .A0(\us21/n319 ), .A1(\us21/n52 ), .B0(\us21/n320 ), 
        .B1(\us21/n114 ), .C0(\us21/n321 ), .Y(\us21/n304 ) );
  NOR2X1 \us21/U272  ( .A(\us21/n226 ), .B(\us21/n58 ), .Y(\us21/n290 ) );
  INVX1 \us21/U271  ( .A(\us21/n290 ), .Y(\us21/n200 ) );
  NAND2X1 \us21/U270  ( .A(\us21/n34 ), .B(\us21/n200 ), .Y(\us21/n120 ) );
  INVX1 \us21/U269  ( .A(\us21/n210 ), .Y(\us21/n100 ) );
  OAI221XL \us21/U268  ( .A0(\us21/n20 ), .A1(\us21/n100 ), .B0(sa21[3]), .B1(
        \us21/n4 ), .C0(\us21/n262 ), .Y(\us21/n317 ) );
  INVX1 \us21/U267  ( .A(\us21/n258 ), .Y(\us21/n182 ) );
  AOI211X1 \us21/U266  ( .A0(\us21/n33 ), .A1(\us21/n120 ), .B0(\us21/n317 ), 
        .C0(\us21/n318 ), .Y(\us21/n306 ) );
  NAND2X1 \us21/U265  ( .A(\us21/n100 ), .B(\us21/n199 ), .Y(\us21/n151 ) );
  INVX1 \us21/U264  ( .A(\us21/n151 ), .Y(\us21/n314 ) );
  NOR2X1 \us21/U263  ( .A(\us21/n45 ), .B(\us21/n163 ), .Y(\us21/n160 ) );
  INVX1 \us21/U262  ( .A(\us21/n295 ), .Y(\us21/n92 ) );
  AOI21X1 \us21/U261  ( .A0(sa21[1]), .A1(\us21/n58 ), .B0(\us21/n98 ), .Y(
        \us21/n316 ) );
  OAI22X1 \us21/U260  ( .A0(\us21/n92 ), .A1(\us21/n18 ), .B0(\us21/n316 ), 
        .B1(\us21/n27 ), .Y(\us21/n315 ) );
  NOR2X1 \us21/U259  ( .A(\us21/n149 ), .B(\us21/n226 ), .Y(\us21/n41 ) );
  INVX1 \us21/U258  ( .A(\us21/n41 ), .Y(\us21/n105 ) );
  NAND2X1 \us21/U257  ( .A(\us21/n284 ), .B(\us21/n105 ), .Y(\us21/n227 ) );
  AOI21X1 \us21/U256  ( .A0(\us21/n313 ), .A1(\us21/n33 ), .B0(\us21/n269 ), 
        .Y(\us21/n312 ) );
  OAI221XL \us21/U255  ( .A0(\us21/n149 ), .A1(\us21/n20 ), .B0(\us21/n4 ), 
        .B1(\us21/n227 ), .C0(\us21/n312 ), .Y(\us21/n309 ) );
  AOI21X1 \us21/U254  ( .A0(\us21/n226 ), .A1(\us21/n188 ), .B0(\us21/n242 ), 
        .Y(\us21/n185 ) );
  INVX1 \us21/U253  ( .A(\us21/n185 ), .Y(\us21/n48 ) );
  AND2X1 \us21/U252  ( .A(\us21/n223 ), .B(\us21/n240 ), .Y(\us21/n28 ) );
  OAI221XL \us21/U251  ( .A0(\us21/n27 ), .A1(\us21/n44 ), .B0(\us21/n4 ), 
        .B1(\us21/n48 ), .C0(\us21/n311 ), .Y(\us21/n310 ) );
  AOI22X1 \us21/U250  ( .A0(\us21/n89 ), .A1(\us21/n309 ), .B0(\us21/n55 ), 
        .B1(\us21/n310 ), .Y(\us21/n308 ) );
  OAI221XL \us21/U249  ( .A0(\us21/n306 ), .A1(\us21/n52 ), .B0(\us21/n307 ), 
        .B1(\us21/n114 ), .C0(\us21/n308 ), .Y(\us21/n305 ) );
  MX2X1 \us21/U248  ( .A(\us21/n304 ), .B(\us21/n305 ), .S0(sa21[6]), .Y(
        sa23_sr[1]) );
  INVX1 \us21/U247  ( .A(\us21/n187 ), .Y(\us21/n61 ) );
  MXI2X1 \us21/U246  ( .A(\us21/n303 ), .B(\us21/n61 ), .S0(\us21/n69 ), .Y(
        \us21/n301 ) );
  MXI2X1 \us21/U245  ( .A(\us21/n301 ), .B(\us21/n147 ), .S0(\us21/n302 ), .Y(
        \us21/n285 ) );
  NAND2X1 \us21/U244  ( .A(\us21/n200 ), .B(\us21/n300 ), .Y(\us21/n99 ) );
  INVX1 \us21/U243  ( .A(\us21/n99 ), .Y(\us21/n296 ) );
  NOR2X1 \us21/U242  ( .A(\us21/n299 ), .B(\us21/n242 ), .Y(\us21/n298 ) );
  NAND2X1 \us21/U241  ( .A(sa21[1]), .B(\us21/n47 ), .Y(\us21/n122 ) );
  NOR2X1 \us21/U240  ( .A(\us21/n159 ), .B(\us21/n217 ), .Y(\us21/n198 ) );
  OAI221XL \us21/U239  ( .A0(\us21/n298 ), .A1(\us21/n27 ), .B0(\us21/n20 ), 
        .B1(\us21/n122 ), .C0(\us21/n132 ), .Y(\us21/n297 ) );
  AOI221X1 \us21/U238  ( .A0(\us21/n225 ), .A1(\us21/n226 ), .B0(\us21/n296 ), 
        .B1(\us21/n6 ), .C0(\us21/n297 ), .Y(\us21/n291 ) );
  OAI2BB2X1 \us21/U237  ( .B0(\us21/n27 ), .B1(\us21/n295 ), .A0N(\us21/n34 ), 
        .A1N(\us21/n24 ), .Y(\us21/n293 ) );
  AOI21X1 \us21/U236  ( .A0(\us21/n101 ), .A1(\us21/n150 ), .B0(\us21/n20 ), 
        .Y(\us21/n294 ) );
  AOI211X1 \us21/U235  ( .A0(\us21/n5 ), .A1(\us21/n79 ), .B0(\us21/n293 ), 
        .C0(\us21/n294 ), .Y(\us21/n292 ) );
  INVX1 \us21/U234  ( .A(\us21/n89 ), .Y(\us21/n10 ) );
  OAI22X1 \us21/U233  ( .A0(\us21/n291 ), .A1(\us21/n114 ), .B0(\us21/n292 ), 
        .B1(\us21/n10 ), .Y(\us21/n286 ) );
  INVX1 \us21/U232  ( .A(\us21/n225 ), .Y(\us21/n288 ) );
  NAND2X1 \us21/U231  ( .A(\us21/n200 ), .B(\us21/n284 ), .Y(\us21/n102 ) );
  NOR2X1 \us21/U230  ( .A(\us21/n290 ), .B(\us21/n163 ), .Y(\us21/n184 ) );
  AOI22X1 \us21/U229  ( .A0(\us21/n102 ), .A1(\us21/n69 ), .B0(\us21/n184 ), 
        .B1(\us21/n33 ), .Y(\us21/n289 ) );
  AOI31X1 \us21/U228  ( .A0(\us21/n132 ), .A1(\us21/n288 ), .A2(\us21/n289 ), 
        .B0(\us21/n52 ), .Y(\us21/n287 ) );
  AOI211X1 \us21/U227  ( .A0(\us21/n285 ), .A1(\us21/n55 ), .B0(\us21/n286 ), 
        .C0(\us21/n287 ), .Y(\us21/n263 ) );
  NAND2X1 \us21/U226  ( .A(\us21/n284 ), .B(\us21/n122 ), .Y(\us21/n125 ) );
  NOR2X1 \us21/U225  ( .A(\us21/n199 ), .B(\us21/n4 ), .Y(\us21/n50 ) );
  AOI21X1 \us21/U224  ( .A0(\us21/n200 ), .A1(\us21/n223 ), .B0(\us21/n20 ), 
        .Y(\us21/n283 ) );
  AOI211X1 \us21/U223  ( .A0(\us21/n5 ), .A1(\us21/n125 ), .B0(\us21/n50 ), 
        .C0(\us21/n283 ), .Y(\us21/n282 ) );
  OAI221XL \us21/U222  ( .A0(\us21/n281 ), .A1(\us21/n27 ), .B0(\us21/n4 ), 
        .B1(\us21/n111 ), .C0(\us21/n282 ), .Y(\us21/n265 ) );
  INVX1 \us21/U221  ( .A(\us21/n280 ), .Y(\us21/n247 ) );
  NAND2X1 \us21/U220  ( .A(\us21/n41 ), .B(\us21/n33 ), .Y(\us21/n272 ) );
  OAI221XL \us21/U219  ( .A0(sa21[1]), .A1(\us21/n247 ), .B0(\us21/n4 ), .B1(
        \us21/n189 ), .C0(\us21/n272 ), .Y(\us21/n279 ) );
  NAND2X1 \us21/U218  ( .A(sa21[2]), .B(\us21/n149 ), .Y(\us21/n276 ) );
  XNOR2X1 \us21/U217  ( .A(\us21/n129 ), .B(sa21[1]), .Y(\us21/n155 ) );
  MXI2X1 \us21/U216  ( .A(\us21/n276 ), .B(\us21/n277 ), .S0(\us21/n155 ), .Y(
        \us21/n275 ) );
  OAI22X1 \us21/U215  ( .A0(\us21/n273 ), .A1(\us21/n10 ), .B0(\us21/n274 ), 
        .B1(\us21/n52 ), .Y(\us21/n266 ) );
  NOR2X1 \us21/U214  ( .A(\us21/n20 ), .B(\us21/n226 ), .Y(\us21/n176 ) );
  OAI21XL \us21/U213  ( .A0(\us21/n4 ), .A1(\us21/n271 ), .B0(\us21/n272 ), 
        .Y(\us21/n270 ) );
  OAI31X1 \us21/U212  ( .A0(\us21/n176 ), .A1(\us21/n269 ), .A2(\us21/n270 ), 
        .B0(\us21/n16 ), .Y(\us21/n268 ) );
  INVX1 \us21/U211  ( .A(\us21/n268 ), .Y(\us21/n267 ) );
  AOI211X1 \us21/U210  ( .A0(\us21/n55 ), .A1(\us21/n265 ), .B0(\us21/n266 ), 
        .C0(\us21/n267 ), .Y(\us21/n264 ) );
  MXI2X1 \us21/U209  ( .A(\us21/n263 ), .B(\us21/n264 ), .S0(sa21[6]), .Y(
        sa23_sr[2]) );
  NOR2X1 \us21/U208  ( .A(\us21/n94 ), .B(sa21[1]), .Y(\us21/n211 ) );
  INVX1 \us21/U207  ( .A(\us21/n262 ), .Y(\us21/n261 ) );
  AOI211X1 \us21/U206  ( .A0(\us21/n259 ), .A1(\us21/n24 ), .B0(\us21/n260 ), 
        .C0(\us21/n261 ), .Y(\us21/n255 ) );
  OAI22X1 \us21/U205  ( .A0(\us21/n20 ), .A1(\us21/n68 ), .B0(\us21/n27 ), 
        .B1(\us21/n37 ), .Y(\us21/n257 ) );
  NOR3X1 \us21/U204  ( .A(\us21/n257 ), .B(\us21/n258 ), .C(\us21/n50 ), .Y(
        \us21/n256 ) );
  MXI2X1 \us21/U203  ( .A(\us21/n255 ), .B(\us21/n256 ), .S0(\us21/n252 ), .Y(
        \us21/n254 ) );
  AOI221X1 \us21/U202  ( .A0(\us21/n211 ), .A1(\us21/n5 ), .B0(\us21/n40 ), 
        .B1(sa21[4]), .C0(\us21/n254 ), .Y(\us21/n248 ) );
  INVX1 \us21/U201  ( .A(\us21/n211 ), .Y(\us21/n106 ) );
  NAND2X1 \us21/U200  ( .A(\us21/n200 ), .B(\us21/n106 ), .Y(\us21/n83 ) );
  NAND2X1 \us21/U199  ( .A(\us21/n199 ), .B(\us21/n204 ), .Y(\us21/n169 ) );
  AOI2BB2X1 \us21/U198  ( .B0(\us21/n65 ), .B1(\us21/n24 ), .A0N(\us21/n169 ), 
        .A1N(\us21/n20 ), .Y(\us21/n253 ) );
  OAI221XL \us21/U197  ( .A0(\us21/n172 ), .A1(\us21/n18 ), .B0(\us21/n27 ), 
        .B1(\us21/n83 ), .C0(\us21/n253 ), .Y(\us21/n251 ) );
  MXI2X1 \us21/U196  ( .A(\us21/n250 ), .B(\us21/n251 ), .S0(\us21/n252 ), .Y(
        \us21/n249 ) );
  MXI2X1 \us21/U195  ( .A(\us21/n248 ), .B(\us21/n249 ), .S0(\us21/n234 ), .Y(
        \us21/n228 ) );
  OAI21XL \us21/U194  ( .A0(\us21/n58 ), .A1(\us21/n27 ), .B0(\us21/n247 ), 
        .Y(\us21/n245 ) );
  NOR2X1 \us21/U193  ( .A(sa21[7]), .B(\us21/n145 ), .Y(\us21/n246 ) );
  XNOR2X1 \us21/U192  ( .A(\us21/n69 ), .B(sa21[1]), .Y(\us21/n130 ) );
  MXI2X1 \us21/U191  ( .A(\us21/n245 ), .B(\us21/n246 ), .S0(\us21/n130 ), .Y(
        \us21/n243 ) );
  OAI211X1 \us21/U190  ( .A0(\us21/n4 ), .A1(\us21/n149 ), .B0(\us21/n243 ), 
        .C0(\us21/n244 ), .Y(\us21/n230 ) );
  NOR2X1 \us21/U189  ( .A(\us21/n242 ), .B(\us21/n137 ), .Y(\us21/n70 ) );
  OAI221XL \us21/U188  ( .A0(\us21/n159 ), .A1(\us21/n27 ), .B0(\us21/n20 ), 
        .B1(\us21/n34 ), .C0(\us21/n241 ), .Y(\us21/n231 ) );
  NAND2X1 \us21/U187  ( .A(\us21/n101 ), .B(\us21/n240 ), .Y(\us21/n76 ) );
  AOI21X1 \us21/U186  ( .A0(\us21/n122 ), .A1(\us21/n106 ), .B0(\us21/n129 ), 
        .Y(\us21/n237 ) );
  INVX1 \us21/U185  ( .A(\us21/n239 ), .Y(\us21/n238 ) );
  OAI21XL \us21/U184  ( .A0(\us21/n237 ), .A1(\us21/n43 ), .B0(\us21/n238 ), 
        .Y(\us21/n236 ) );
  OAI221XL \us21/U183  ( .A0(\us21/n18 ), .A1(\us21/n76 ), .B0(\us21/n59 ), 
        .B1(\us21/n27 ), .C0(\us21/n236 ), .Y(\us21/n232 ) );
  AOI2BB2X1 \us21/U182  ( .B0(\us21/n24 ), .B1(\us21/n187 ), .A0N(\us21/n227 ), 
        .A1N(\us21/n20 ), .Y(\us21/n235 ) );
  OAI211X1 \us21/U181  ( .A0(\us21/n27 ), .A1(\us21/n122 ), .B0(\us21/n158 ), 
        .C0(\us21/n235 ), .Y(\us21/n233 ) );
  MX4X1 \us21/U180  ( .A(\us21/n230 ), .B(\us21/n231 ), .C(\us21/n232 ), .D(
        \us21/n233 ), .S0(\us21/n234 ), .S1(sa21[5]), .Y(\us21/n229 ) );
  MX2X1 \us21/U179  ( .A(\us21/n228 ), .B(\us21/n229 ), .S0(sa21[6]), .Y(
        sa23_sr[3]) );
  NOR2BX1 \us21/U178  ( .AN(\us21/n204 ), .B(\us21/n137 ), .Y(\us21/n110 ) );
  INVX1 \us21/U177  ( .A(\us21/n110 ), .Y(\us21/n64 ) );
  AOI22X1 \us21/U176  ( .A0(\us21/n225 ), .A1(\us21/n226 ), .B0(\us21/n6 ), 
        .B1(\us21/n227 ), .Y(\us21/n224 ) );
  OAI221XL \us21/U175  ( .A0(\us21/n27 ), .A1(\us21/n64 ), .B0(\us21/n4 ), 
        .B1(\us21/n83 ), .C0(\us21/n224 ), .Y(\us21/n212 ) );
  NAND2X1 \us21/U174  ( .A(\us21/n34 ), .B(\us21/n204 ), .Y(\us21/n221 ) );
  OAI21XL \us21/U173  ( .A0(\us21/n69 ), .A1(\us21/n223 ), .B0(\us21/n27 ), 
        .Y(\us21/n222 ) );
  NOR2X1 \us21/U172  ( .A(\us21/n217 ), .B(\us21/n42 ), .Y(\us21/n208 ) );
  AOI211X1 \us21/U171  ( .A0(\us21/n208 ), .A1(\us21/n5 ), .B0(\us21/n220 ), 
        .C0(\us21/n173 ), .Y(\us21/n219 ) );
  OAI22X1 \us21/U170  ( .A0(\us21/n218 ), .A1(\us21/n10 ), .B0(\us21/n219 ), 
        .B1(\us21/n114 ), .Y(\us21/n213 ) );
  INVX1 \us21/U169  ( .A(\us21/n135 ), .Y(\us21/n215 ) );
  NOR2X1 \us21/U168  ( .A(\us21/n4 ), .B(\us21/n159 ), .Y(\us21/n31 ) );
  INVX1 \us21/U167  ( .A(\us21/n31 ), .Y(\us21/n196 ) );
  AOI31X1 \us21/U166  ( .A0(\us21/n215 ), .A1(\us21/n196 ), .A2(\us21/n216 ), 
        .B0(\us21/n52 ), .Y(\us21/n214 ) );
  AOI211X1 \us21/U165  ( .A0(\us21/n55 ), .A1(\us21/n212 ), .B0(\us21/n213 ), 
        .C0(\us21/n214 ), .Y(\us21/n190 ) );
  INVX1 \us21/U164  ( .A(\us21/n207 ), .Y(\us21/n192 ) );
  NOR2X1 \us21/U163  ( .A(\us21/n25 ), .B(\us21/n98 ), .Y(\us21/n32 ) );
  OAI22X1 \us21/U162  ( .A0(\us21/n28 ), .A1(\us21/n4 ), .B0(\us21/n188 ), 
        .B1(\us21/n27 ), .Y(\us21/n206 ) );
  NAND2X1 \us21/U161  ( .A(\us21/n204 ), .B(\us21/n80 ), .Y(\us21/n118 ) );
  INVX1 \us21/U160  ( .A(\us21/n118 ), .Y(\us21/n123 ) );
  NAND2X1 \us21/U159  ( .A(\us21/n94 ), .B(\us21/n79 ), .Y(\us21/n203 ) );
  OAI2BB1X1 \us21/U158  ( .A0N(\us21/n199 ), .A1N(\us21/n200 ), .B0(\us21/n33 ), .Y(\us21/n195 ) );
  INVX1 \us21/U157  ( .A(\us21/n55 ), .Y(\us21/n12 ) );
  AOI31X1 \us21/U156  ( .A0(\us21/n195 ), .A1(\us21/n196 ), .A2(\us21/n197 ), 
        .B0(\us21/n12 ), .Y(\us21/n194 ) );
  AOI211X1 \us21/U155  ( .A0(\us21/n89 ), .A1(\us21/n192 ), .B0(\us21/n193 ), 
        .C0(\us21/n194 ), .Y(\us21/n191 ) );
  MXI2X1 \us21/U154  ( .A(\us21/n190 ), .B(\us21/n191 ), .S0(sa21[6]), .Y(
        sa23_sr[4]) );
  OAI21XL \us21/U153  ( .A0(\us21/n69 ), .A1(\us21/n189 ), .B0(\us21/n27 ), 
        .Y(\us21/n186 ) );
  INVX1 \us21/U152  ( .A(\us21/n183 ), .Y(\us21/n180 ) );
  NAND2X1 \us21/U151  ( .A(\us21/n74 ), .B(\us21/n182 ), .Y(\us21/n181 ) );
  AOI211X1 \us21/U150  ( .A0(\us21/n179 ), .A1(\us21/n24 ), .B0(\us21/n180 ), 
        .C0(\us21/n181 ), .Y(\us21/n165 ) );
  INVX1 \us21/U149  ( .A(\us21/n178 ), .Y(\us21/n175 ) );
  AOI211X1 \us21/U148  ( .A0(\us21/n175 ), .A1(\us21/n5 ), .B0(\us21/n176 ), 
        .C0(\us21/n177 ), .Y(\us21/n174 ) );
  OAI221XL \us21/U147  ( .A0(\us21/n159 ), .A1(\us21/n27 ), .B0(\us21/n145 ), 
        .B1(\us21/n20 ), .C0(\us21/n174 ), .Y(\us21/n167 ) );
  MXI2X1 \us21/U146  ( .A(\us21/n40 ), .B(\us21/n173 ), .S0(\us21/n96 ), .Y(
        \us21/n170 ) );
  AOI22X1 \us21/U145  ( .A0(\us21/n137 ), .A1(\us21/n24 ), .B0(\us21/n172 ), 
        .B1(\us21/n6 ), .Y(\us21/n171 ) );
  OAI211X1 \us21/U144  ( .A0(\us21/n20 ), .A1(\us21/n169 ), .B0(\us21/n170 ), 
        .C0(\us21/n171 ), .Y(\us21/n168 ) );
  AOI22X1 \us21/U143  ( .A0(\us21/n89 ), .A1(\us21/n167 ), .B0(\us21/n55 ), 
        .B1(\us21/n168 ), .Y(\us21/n166 ) );
  OAI221XL \us21/U142  ( .A0(\us21/n164 ), .A1(\us21/n114 ), .B0(\us21/n165 ), 
        .B1(\us21/n52 ), .C0(\us21/n166 ), .Y(\us21/n138 ) );
  OAI21XL \us21/U141  ( .A0(\us21/n41 ), .A1(\us21/n163 ), .B0(\us21/n69 ), 
        .Y(\us21/n162 ) );
  AOI221X1 \us21/U140  ( .A0(\us21/n159 ), .A1(\us21/n24 ), .B0(\us21/n160 ), 
        .B1(\us21/n33 ), .C0(\us21/n161 ), .Y(\us21/n140 ) );
  OAI21XL \us21/U139  ( .A0(\us21/n157 ), .A1(\us21/n20 ), .B0(\us21/n158 ), 
        .Y(\us21/n156 ) );
  NOR2X1 \us21/U138  ( .A(\us21/n4 ), .B(\us21/n136 ), .Y(\us21/n153 ) );
  NOR2X1 \us21/U137  ( .A(\us21/n145 ), .B(\us21/n69 ), .Y(\us21/n154 ) );
  MXI2X1 \us21/U136  ( .A(\us21/n153 ), .B(\us21/n154 ), .S0(\us21/n155 ), .Y(
        \us21/n152 ) );
  OAI221XL \us21/U135  ( .A0(\us21/n110 ), .A1(\us21/n18 ), .B0(\us21/n20 ), 
        .B1(\us21/n151 ), .C0(\us21/n152 ), .Y(\us21/n143 ) );
  AOI21X1 \us21/U134  ( .A0(\us21/n149 ), .A1(\us21/n150 ), .B0(\us21/n18 ), 
        .Y(\us21/n148 ) );
  AOI2BB1X1 \us21/U133  ( .A0N(\us21/n147 ), .A1N(\us21/n27 ), .B0(\us21/n148 ), .Y(\us21/n146 ) );
  OAI221XL \us21/U132  ( .A0(\us21/n145 ), .A1(\us21/n20 ), .B0(\us21/n4 ), 
        .B1(\us21/n34 ), .C0(\us21/n146 ), .Y(\us21/n144 ) );
  AOI22X1 \us21/U131  ( .A0(\us21/n89 ), .A1(\us21/n143 ), .B0(\us21/n14 ), 
        .B1(\us21/n144 ), .Y(\us21/n142 ) );
  OAI221XL \us21/U130  ( .A0(\us21/n140 ), .A1(\us21/n12 ), .B0(\us21/n141 ), 
        .B1(\us21/n114 ), .C0(\us21/n142 ), .Y(\us21/n139 ) );
  MX2X1 \us21/U129  ( .A(\us21/n138 ), .B(\us21/n139 ), .S0(sa21[6]), .Y(
        sa23_sr[5]) );
  INVX1 \us21/U128  ( .A(\us21/n70 ), .Y(\us21/n133 ) );
  OAI22X1 \us21/U127  ( .A0(\us21/n4 ), .A1(\us21/n136 ), .B0(\us21/n137 ), 
        .B1(\us21/n27 ), .Y(\us21/n134 ) );
  AOI211X1 \us21/U126  ( .A0(\us21/n133 ), .A1(\us21/n69 ), .B0(\us21/n134 ), 
        .C0(\us21/n135 ), .Y(\us21/n112 ) );
  INVX1 \us21/U125  ( .A(\us21/n132 ), .Y(\us21/n131 ) );
  OAI21XL \us21/U124  ( .A0(\us21/n18 ), .A1(\us21/n37 ), .B0(\us21/n128 ), 
        .Y(\us21/n127 ) );
  OAI221XL \us21/U123  ( .A0(\us21/n18 ), .A1(\us21/n105 ), .B0(\us21/n123 ), 
        .B1(\us21/n27 ), .C0(\us21/n124 ), .Y(\us21/n116 ) );
  NAND2X1 \us21/U122  ( .A(\us21/n121 ), .B(\us21/n122 ), .Y(\us21/n30 ) );
  OAI221XL \us21/U121  ( .A0(\us21/n18 ), .A1(\us21/n118 ), .B0(\us21/n27 ), 
        .B1(\us21/n30 ), .C0(\us21/n119 ), .Y(\us21/n117 ) );
  AOI22X1 \us21/U120  ( .A0(\us21/n89 ), .A1(\us21/n116 ), .B0(\us21/n55 ), 
        .B1(\us21/n117 ), .Y(\us21/n115 ) );
  OAI221XL \us21/U119  ( .A0(\us21/n112 ), .A1(\us21/n52 ), .B0(\us21/n113 ), 
        .B1(\us21/n114 ), .C0(\us21/n115 ), .Y(\us21/n84 ) );
  OAI22X1 \us21/U118  ( .A0(\us21/n110 ), .A1(\us21/n4 ), .B0(\us21/n20 ), 
        .B1(\us21/n21 ), .Y(\us21/n108 ) );
  AOI21X1 \us21/U117  ( .A0(sa21[1]), .A1(\us21/n58 ), .B0(\us21/n27 ), .Y(
        \us21/n109 ) );
  AOI211X1 \us21/U116  ( .A0(\us21/n5 ), .A1(\us21/n107 ), .B0(\us21/n108 ), 
        .C0(\us21/n109 ), .Y(\us21/n86 ) );
  OAI22X1 \us21/U115  ( .A0(\us21/n45 ), .A1(\us21/n4 ), .B0(sa21[4]), .B1(
        \us21/n18 ), .Y(\us21/n103 ) );
  AOI21X1 \us21/U114  ( .A0(\us21/n105 ), .A1(\us21/n106 ), .B0(\us21/n20 ), 
        .Y(\us21/n104 ) );
  AOI211X1 \us21/U113  ( .A0(\us21/n33 ), .A1(\us21/n102 ), .B0(\us21/n103 ), 
        .C0(\us21/n104 ), .Y(\us21/n87 ) );
  NAND2X1 \us21/U112  ( .A(\us21/n100 ), .B(\us21/n101 ), .Y(\us21/n62 ) );
  OAI221XL \us21/U111  ( .A0(\us21/n27 ), .A1(\us21/n62 ), .B0(\us21/n4 ), 
        .B1(\us21/n21 ), .C0(\us21/n97 ), .Y(\us21/n90 ) );
  NOR3X1 \us21/U110  ( .A(\us21/n4 ), .B(\us21/n95 ), .C(\us21/n96 ), .Y(
        \us21/n67 ) );
  AOI31X1 \us21/U109  ( .A0(\us21/n79 ), .A1(\us21/n94 ), .A2(\us21/n6 ), .B0(
        \us21/n67 ), .Y(\us21/n93 ) );
  OAI221XL \us21/U108  ( .A0(\us21/n73 ), .A1(\us21/n27 ), .B0(\us21/n92 ), 
        .B1(\us21/n20 ), .C0(\us21/n93 ), .Y(\us21/n91 ) );
  AOI22X1 \us21/U107  ( .A0(\us21/n89 ), .A1(\us21/n90 ), .B0(\us21/n16 ), 
        .B1(\us21/n91 ), .Y(\us21/n88 ) );
  OAI221XL \us21/U106  ( .A0(\us21/n86 ), .A1(\us21/n52 ), .B0(\us21/n87 ), 
        .B1(\us21/n12 ), .C0(\us21/n88 ), .Y(\us21/n85 ) );
  MX2X1 \us21/U105  ( .A(\us21/n84 ), .B(\us21/n85 ), .S0(sa21[6]), .Y(
        sa23_sr[6]) );
  INVX1 \us21/U104  ( .A(\us21/n81 ), .Y(\us21/n77 ) );
  AOI21X1 \us21/U103  ( .A0(\us21/n79 ), .A1(\us21/n80 ), .B0(\us21/n27 ), .Y(
        \us21/n78 ) );
  AOI211X1 \us21/U102  ( .A0(\us21/n5 ), .A1(\us21/n76 ), .B0(\us21/n77 ), 
        .C0(\us21/n78 ), .Y(\us21/n51 ) );
  OAI211X1 \us21/U101  ( .A0(\us21/n73 ), .A1(\us21/n27 ), .B0(\us21/n74 ), 
        .C0(\us21/n75 ), .Y(\us21/n72 ) );
  AOI21X1 \us21/U100  ( .A0(\us21/n68 ), .A1(\us21/n69 ), .B0(\us21/n6 ), .Y(
        \us21/n63 ) );
  INVX1 \us21/U99  ( .A(\us21/n67 ), .Y(\us21/n66 ) );
  OAI221XL \us21/U98  ( .A0(\us21/n63 ), .A1(\us21/n64 ), .B0(\us21/n65 ), 
        .B1(\us21/n27 ), .C0(\us21/n66 ), .Y(\us21/n56 ) );
  AOI2BB2X1 \us21/U97  ( .B0(\us21/n61 ), .B1(\us21/n24 ), .A0N(\us21/n62 ), 
        .A1N(\us21/n20 ), .Y(\us21/n60 ) );
  OAI221XL \us21/U96  ( .A0(\us21/n58 ), .A1(\us21/n18 ), .B0(\us21/n59 ), 
        .B1(\us21/n27 ), .C0(\us21/n60 ), .Y(\us21/n57 ) );
  AOI22X1 \us21/U95  ( .A0(\us21/n55 ), .A1(\us21/n56 ), .B0(\us21/n16 ), .B1(
        \us21/n57 ), .Y(\us21/n54 ) );
  OAI221XL \us21/U94  ( .A0(\us21/n51 ), .A1(\us21/n52 ), .B0(\us21/n53 ), 
        .B1(\us21/n10 ), .C0(\us21/n54 ), .Y(\us21/n7 ) );
  INVX1 \us21/U93  ( .A(\us21/n50 ), .Y(\us21/n49 ) );
  OAI221XL \us21/U92  ( .A0(\us21/n47 ), .A1(\us21/n18 ), .B0(\us21/n27 ), 
        .B1(\us21/n48 ), .C0(\us21/n49 ), .Y(\us21/n46 ) );
  NOR2X1 \us21/U91  ( .A(\us21/n41 ), .B(\us21/n42 ), .Y(\us21/n38 ) );
  INVX1 \us21/U90  ( .A(\us21/n40 ), .Y(\us21/n39 ) );
  INVX1 \us21/U89  ( .A(\us21/n32 ), .Y(\us21/n26 ) );
  AOI21X1 \us21/U88  ( .A0(\us21/n5 ), .A1(\us21/n30 ), .B0(\us21/n31 ), .Y(
        \us21/n29 ) );
  OAI221XL \us21/U87  ( .A0(\us21/n26 ), .A1(\us21/n27 ), .B0(\us21/n28 ), 
        .B1(\us21/n20 ), .C0(\us21/n29 ), .Y(\us21/n15 ) );
  OAI221XL \us21/U86  ( .A0(\us21/n18 ), .A1(\us21/n19 ), .B0(\us21/n20 ), 
        .B1(\us21/n21 ), .C0(\us21/n22 ), .Y(\us21/n17 ) );
  AOI22X1 \us21/U85  ( .A0(\us21/n14 ), .A1(\us21/n15 ), .B0(\us21/n16 ), .B1(
        \us21/n17 ), .Y(\us21/n13 ) );
  OAI221XL \us21/U84  ( .A0(\us21/n9 ), .A1(\us21/n10 ), .B0(\us21/n11 ), .B1(
        \us21/n12 ), .C0(\us21/n13 ), .Y(\us21/n8 ) );
  MX2X1 \us21/U83  ( .A(\us21/n7 ), .B(\us21/n8 ), .S0(sa21[6]), .Y(sa23_sr[7]) );
  NOR2X4 \us21/U82  ( .A(\us21/n129 ), .B(sa21[2]), .Y(\us21/n43 ) );
  CLKINVX3 \us21/U81  ( .A(\us21/n14 ), .Y(\us21/n52 ) );
  OAI22XL \us21/U80  ( .A0(\us21/n201 ), .A1(\us21/n52 ), .B0(\us21/n202 ), 
        .B1(\us21/n114 ), .Y(\us21/n193 ) );
  CLKINVX3 \us21/U79  ( .A(sa21[5]), .Y(\us21/n252 ) );
  NOR2X2 \us21/U78  ( .A(\us21/n252 ), .B(\us21/n234 ), .Y(\us21/n55 ) );
  CLKINVX3 \us21/U77  ( .A(sa21[7]), .Y(\us21/n129 ) );
  NOR2X4 \us21/U76  ( .A(\us21/n129 ), .B(\us21/n69 ), .Y(\us21/n24 ) );
  AOI22XL \us21/U75  ( .A0(\us21/n70 ), .A1(\us21/n24 ), .B0(\us21/n96 ), .B1(
        \us21/n129 ), .Y(\us21/n241 ) );
  NOR2X2 \us21/U74  ( .A(\us21/n252 ), .B(sa21[0]), .Y(\us21/n89 ) );
  CLKINVX3 \us21/U73  ( .A(sa21[0]), .Y(\us21/n234 ) );
  NOR2X4 \us21/U72  ( .A(\us21/n69 ), .B(sa21[7]), .Y(\us21/n33 ) );
  INVX12 \us21/U71  ( .A(\us21/n33 ), .Y(\us21/n27 ) );
  CLKINVX3 \us21/U70  ( .A(\us21/n1 ), .Y(\us21/n6 ) );
  CLKINVX3 \us21/U69  ( .A(\us21/n1 ), .Y(\us21/n5 ) );
  INVXL \us21/U68  ( .A(\us21/n24 ), .Y(\us21/n36 ) );
  INVX4 \us21/U67  ( .A(\us21/n3 ), .Y(\us21/n4 ) );
  INVXL \us21/U66  ( .A(\us21/n36 ), .Y(\us21/n3 ) );
  INVX4 \us21/U65  ( .A(sa21[1]), .Y(\us21/n226 ) );
  INVX4 \us21/U64  ( .A(\us21/n43 ), .Y(\us21/n20 ) );
  AOI221X4 \us21/U63  ( .A0(\us21/n24 ), .A1(\us21/n82 ), .B0(\us21/n43 ), 
        .B1(\us21/n295 ), .C0(\us21/n173 ), .Y(\us21/n346 ) );
  AOI221X4 \us21/U62  ( .A0(\us21/n5 ), .A1(\us21/n96 ), .B0(\us21/n43 ), .B1(
        \us21/n239 ), .C0(\us21/n340 ), .Y(\us21/n336 ) );
  AOI222X4 \us21/U61  ( .A0(\us21/n59 ), .A1(\us21/n43 ), .B0(\us21/n6 ), .B1(
        \us21/n221 ), .C0(\us21/n222 ), .C1(\us21/n187 ), .Y(\us21/n218 ) );
  AOI222X4 \us21/U60  ( .A0(\us21/n123 ), .A1(\us21/n43 ), .B0(sa21[2]), .B1(
        \us21/n203 ), .C0(\us21/n6 ), .C1(\us21/n71 ), .Y(\us21/n202 ) );
  AOI221X4 \us21/U59  ( .A0(\us21/n314 ), .A1(\us21/n43 ), .B0(\us21/n160 ), 
        .B1(\us21/n24 ), .C0(\us21/n315 ), .Y(\us21/n307 ) );
  AOI221X4 \us21/U58  ( .A0(\us21/n43 ), .A1(\us21/n208 ), .B0(\us21/n76 ), 
        .B1(\us21/n24 ), .C0(\us21/n209 ), .Y(\us21/n207 ) );
  AOI221X4 \us21/U57  ( .A0(\us21/n43 ), .A1(\us21/n205 ), .B0(\us21/n32 ), 
        .B1(\us21/n6 ), .C0(\us21/n206 ), .Y(\us21/n201 ) );
  AOI221X4 \us21/U56  ( .A0(\us21/n43 ), .A1(\us21/n44 ), .B0(\us21/n45 ), 
        .B1(\us21/n24 ), .C0(\us21/n46 ), .Y(\us21/n9 ) );
  AOI22XL \us21/U55  ( .A0(\us21/n217 ), .A1(\us21/n43 ), .B0(\us21/n33 ), 
        .B1(\us21/n47 ), .Y(\us21/n216 ) );
  AOI22XL \us21/U54  ( .A0(\us21/n98 ), .A1(\us21/n43 ), .B0(\us21/n6 ), .B1(
        \us21/n99 ), .Y(\us21/n97 ) );
  AOI22XL \us21/U53  ( .A0(\us21/n82 ), .A1(\us21/n43 ), .B0(\us21/n83 ), .B1(
        \us21/n24 ), .Y(\us21/n81 ) );
  AOI2BB2XL \us21/U52  ( .B0(\us21/n43 ), .B1(\us21/n94 ), .A0N(\us21/n120 ), 
        .A1N(\us21/n4 ), .Y(\us21/n119 ) );
  AOI222X4 \us21/U51  ( .A0(\us21/n125 ), .A1(\us21/n33 ), .B0(\us21/n145 ), 
        .B1(\us21/n40 ), .C0(\us21/n43 ), .C1(\us21/n184 ), .Y(\us21/n183 ) );
  AOI22XL \us21/U50  ( .A0(\us21/n43 ), .A1(\us21/n303 ), .B0(\us21/n24 ), 
        .B1(\us21/n96 ), .Y(\us21/n358 ) );
  AOI22XL \us21/U49  ( .A0(\us21/n43 ), .A1(\us21/n100 ), .B0(\us21/n24 ), 
        .B1(\us21/n125 ), .Y(\us21/n124 ) );
  AOI21XL \us21/U48  ( .A0(\us21/n159 ), .A1(\us21/n43 ), .B0(\us21/n40 ), .Y(
        \us21/n262 ) );
  AOI22XL \us21/U47  ( .A0(\us21/n40 ), .A1(\us21/n94 ), .B0(\us21/n43 ), .B1(
        \us21/n187 ), .Y(\us21/n244 ) );
  AOI22XL \us21/U46  ( .A0(\us21/n184 ), .A1(\us21/n5 ), .B0(\us21/n198 ), 
        .B1(\us21/n43 ), .Y(\us21/n197 ) );
  NOR2XL \us21/U45  ( .A(\us21/n33 ), .B(\us21/n2 ), .Y(\us21/n302 ) );
  MXI2XL \us21/U44  ( .A(\us21/n2 ), .B(\us21/n6 ), .S0(\us21/n28 ), .Y(
        \us21/n311 ) );
  INVXL \us21/U43  ( .A(\us21/n20 ), .Y(\us21/n2 ) );
  INVX4 \us21/U42  ( .A(\us21/n6 ), .Y(\us21/n18 ) );
  AOI21XL \us21/U41  ( .A0(\us21/n18 ), .A1(\us21/n162 ), .B0(\us21/n25 ), .Y(
        \us21/n161 ) );
  INVX4 \us21/U40  ( .A(sa21[2]), .Y(\us21/n69 ) );
  NOR2X4 \us21/U39  ( .A(\us21/n226 ), .B(\us21/n4 ), .Y(\us21/n40 ) );
  CLKINVX3 \us21/U38  ( .A(sa21[3]), .Y(\us21/n136 ) );
  NOR2X2 \us21/U37  ( .A(\us21/n136 ), .B(sa21[4]), .Y(\us21/n145 ) );
  CLKINVX3 \us21/U36  ( .A(sa21[4]), .Y(\us21/n58 ) );
  NOR2X2 \us21/U35  ( .A(\us21/n58 ), .B(sa21[3]), .Y(\us21/n159 ) );
  NOR2X2 \us21/U34  ( .A(\us21/n136 ), .B(\us21/n58 ), .Y(\us21/n259 ) );
  NOR2X2 \us21/U33  ( .A(sa21[4]), .B(sa21[3]), .Y(\us21/n278 ) );
  NOR2X2 \us21/U32  ( .A(\us21/n259 ), .B(\us21/n278 ), .Y(\us21/n47 ) );
  CLKINVX3 \us21/U31  ( .A(\us21/n259 ), .Y(\us21/n44 ) );
  NOR2X2 \us21/U30  ( .A(\us21/n44 ), .B(sa21[1]), .Y(\us21/n137 ) );
  AOI21XL \us21/U29  ( .A0(\us21/n44 ), .A1(\us21/n111 ), .B0(\us21/n4 ), .Y(
        \us21/n177 ) );
  AOI22XL \us21/U28  ( .A0(\us21/n23 ), .A1(\us21/n24 ), .B0(\us21/n25 ), .B1(
        sa21[2]), .Y(\us21/n22 ) );
  AOI22XL \us21/U27  ( .A0(\us21/n33 ), .A1(sa21[3]), .B0(\us21/n24 ), .B1(
        \us21/n58 ), .Y(\us21/n277 ) );
  NAND2XL \us21/U26  ( .A(\us21/n198 ), .B(\us21/n24 ), .Y(\us21/n132 ) );
  OAI2BB2XL \us21/U25  ( .B0(\us21/n20 ), .B1(\us21/n111 ), .A0N(\us21/n125 ), 
        .A1N(\us21/n24 ), .Y(\us21/n220 ) );
  NAND2XL \us21/U24  ( .A(\us21/n111 ), .B(\us21/n101 ), .Y(\us21/n21 ) );
  NAND2XL \us21/U23  ( .A(\us21/n111 ), .B(\us21/n300 ), .Y(\us21/n187 ) );
  NAND2XL \us21/U22  ( .A(\us21/n111 ), .B(\us21/n121 ), .Y(\us21/n303 ) );
  AOI221XL \us21/U21  ( .A0(\us21/n43 ), .A1(\us21/n151 ), .B0(\us21/n25 ), 
        .B1(\us21/n69 ), .C0(\us21/n275 ), .Y(\us21/n274 ) );
  NOR2BXL \us21/U20  ( .AN(\us21/n101 ), .B(\us21/n25 ), .Y(\us21/n172 ) );
  NAND2X2 \us21/U19  ( .A(\us21/n58 ), .B(\us21/n226 ), .Y(\us21/n34 ) );
  OAI222X1 \us21/U18  ( .A0(\us21/n27 ), .A1(\us21/n34 ), .B0(\us21/n69 ), 
        .B1(\us21/n205 ), .C0(\us21/n20 ), .C1(\us21/n79 ), .Y(\us21/n260 ) );
  OAI222X1 \us21/U17  ( .A0(\us21/n20 ), .A1(\us21/n99 ), .B0(\us21/n27 ), 
        .B1(\us21/n101 ), .C0(\us21/n184 ), .C1(\us21/n4 ), .Y(\us21/n250 ) );
  OAI222X1 \us21/U16  ( .A0(\us21/n4 ), .A1(\us21/n37 ), .B0(\us21/n38 ), .B1(
        \us21/n20 ), .C0(sa21[4]), .C1(\us21/n39 ), .Y(\us21/n35 ) );
  AOI221X1 \us21/U15  ( .A0(\us21/n5 ), .A1(\us21/n19 ), .B0(\us21/n33 ), .B1(
        \us21/n34 ), .C0(\us21/n35 ), .Y(\us21/n11 ) );
  OR2X2 \us21/U14  ( .A(sa21[2]), .B(sa21[7]), .Y(\us21/n1 ) );
  AOI221XL \us21/U13  ( .A0(\us21/n59 ), .A1(\us21/n33 ), .B0(\us21/n43 ), 
        .B1(\us21/n126 ), .C0(\us21/n127 ), .Y(\us21/n113 ) );
  AOI221XL \us21/U12  ( .A0(\us21/n70 ), .A1(\us21/n43 ), .B0(\us21/n24 ), 
        .B1(\us21/n71 ), .C0(\us21/n72 ), .Y(\us21/n53 ) );
  AOI221X1 \us21/U11  ( .A0(\us21/n313 ), .A1(\us21/n5 ), .B0(\us21/n23 ), 
        .B1(\us21/n2 ), .C0(\us21/n328 ), .Y(\us21/n320 ) );
  AOI222XL \us21/U10  ( .A0(\us21/n185 ), .A1(\us21/n43 ), .B0(\us21/n186 ), 
        .B1(\us21/n187 ), .C0(\us21/n6 ), .C1(\us21/n188 ), .Y(\us21/n164 ) );
  AOI221X1 \us21/U9  ( .A0(\us21/n40 ), .A1(\us21/n136 ), .B0(\us21/n33 ), 
        .B1(\us21/n178 ), .C0(\us21/n338 ), .Y(\us21/n337 ) );
  AOI222XL \us21/U8  ( .A0(\us21/n278 ), .A1(\us21/n24 ), .B0(\us21/n42 ), 
        .B1(\us21/n33 ), .C0(\us21/n43 ), .C1(\us21/n136 ), .Y(\us21/n351 ) );
  AOI31X1 \us21/U7  ( .A0(sa21[2]), .A1(\us21/n58 ), .A2(sa21[1]), .B0(
        \us21/n40 ), .Y(\us21/n350 ) );
  AOI31X1 \us21/U6  ( .A0(\us21/n44 ), .A1(\us21/n129 ), .A2(\us21/n130 ), 
        .B0(\us21/n131 ), .Y(\us21/n128 ) );
  AOI221X1 \us21/U5  ( .A0(\us21/n278 ), .A1(\us21/n40 ), .B0(\us21/n185 ), 
        .B1(\us21/n2 ), .C0(\us21/n279 ), .Y(\us21/n273 ) );
  OAI32X1 \us21/U4  ( .A0(\us21/n18 ), .A1(sa21[1]), .A2(\us21/n159 ), .B0(
        sa21[4]), .B1(\us21/n182 ), .Y(\us21/n318 ) );
  AOI221X1 \us21/U3  ( .A0(\us21/n40 ), .A1(\us21/n136 ), .B0(\us21/n33 ), 
        .B1(\us21/n47 ), .C0(\us21/n156 ), .Y(\us21/n141 ) );
  OAI32X1 \us21/U2  ( .A0(\us21/n210 ), .A1(\us21/n145 ), .A2(\us21/n18 ), 
        .B0(\us21/n27 ), .B1(\us21/n211 ), .Y(\us21/n209 ) );
  AOI31XL \us21/U1  ( .A0(\us21/n79 ), .A1(\us21/n44 ), .A2(\us21/n2 ), .B0(
        \us21/n280 ), .Y(\us21/n339 ) );
  NAND2X1 \us22/U366  ( .A(\us22/n47 ), .B(\us22/n226 ), .Y(\us22/n189 ) );
  NOR2X1 \us22/U365  ( .A(\us22/n226 ), .B(sa22[3]), .Y(\us22/n242 ) );
  INVX1 \us22/U364  ( .A(\us22/n242 ), .Y(\us22/n205 ) );
  AND2X1 \us22/U363  ( .A(\us22/n189 ), .B(\us22/n205 ), .Y(\us22/n65 ) );
  NOR2X1 \us22/U362  ( .A(\us22/n226 ), .B(\us22/n47 ), .Y(\us22/n45 ) );
  NOR2X1 \us22/U361  ( .A(\us22/n259 ), .B(\us22/n45 ), .Y(\us22/n73 ) );
  NAND2BX1 \us22/U360  ( .AN(\us22/n73 ), .B(\us22/n6 ), .Y(\us22/n158 ) );
  NOR2X1 \us22/U359  ( .A(\us22/n226 ), .B(\us22/n159 ), .Y(\us22/n95 ) );
  INVX1 \us22/U358  ( .A(\us22/n95 ), .Y(\us22/n111 ) );
  NOR2X1 \us22/U357  ( .A(\us22/n145 ), .B(sa22[1]), .Y(\us22/n42 ) );
  INVX1 \us22/U356  ( .A(\us22/n42 ), .Y(\us22/n121 ) );
  INVX1 \us22/U355  ( .A(\us22/n47 ), .Y(\us22/n96 ) );
  OAI211X1 \us22/U354  ( .A0(\us22/n65 ), .A1(\us22/n27 ), .B0(\us22/n158 ), 
        .C0(\us22/n358 ), .Y(\us22/n355 ) );
  NOR2X1 \us22/U353  ( .A(\us22/n226 ), .B(\us22/n145 ), .Y(\us22/n59 ) );
  NOR2X1 \us22/U352  ( .A(\us22/n96 ), .B(\us22/n59 ), .Y(\us22/n271 ) );
  NOR2X1 \us22/U351  ( .A(\us22/n226 ), .B(\us22/n278 ), .Y(\us22/n217 ) );
  INVX1 \us22/U350  ( .A(\us22/n217 ), .Y(\us22/n150 ) );
  NAND2X1 \us22/U349  ( .A(\us22/n44 ), .B(\us22/n150 ), .Y(\us22/n147 ) );
  NAND2X1 \us22/U348  ( .A(sa22[4]), .B(\us22/n226 ), .Y(\us22/n101 ) );
  INVX1 \us22/U347  ( .A(\us22/n159 ), .Y(\us22/n188 ) );
  NOR2X1 \us22/U346  ( .A(\us22/n188 ), .B(\us22/n226 ), .Y(\us22/n25 ) );
  INVX1 \us22/U345  ( .A(\us22/n172 ), .Y(\us22/n107 ) );
  AOI22X1 \us22/U344  ( .A0(\us22/n33 ), .A1(\us22/n147 ), .B0(\us22/n24 ), 
        .B1(\us22/n107 ), .Y(\us22/n357 ) );
  OAI221XL \us22/U343  ( .A0(\us22/n18 ), .A1(\us22/n121 ), .B0(\us22/n271 ), 
        .B1(\us22/n20 ), .C0(\us22/n357 ), .Y(\us22/n356 ) );
  MXI2X1 \us22/U342  ( .A(\us22/n355 ), .B(\us22/n356 ), .S0(\us22/n252 ), .Y(
        \us22/n331 ) );
  INVX1 \us22/U341  ( .A(\us22/n59 ), .Y(\us22/n79 ) );
  AND2X1 \us22/U340  ( .A(\us22/n101 ), .B(\us22/n79 ), .Y(\us22/n325 ) );
  XNOR2X1 \us22/U339  ( .A(sa22[5]), .B(\us22/n226 ), .Y(\us22/n352 ) );
  NOR2X1 \us22/U338  ( .A(\us22/n226 ), .B(\us22/n136 ), .Y(\us22/n281 ) );
  INVX1 \us22/U337  ( .A(\us22/n281 ), .Y(\us22/n19 ) );
  NAND2X1 \us22/U336  ( .A(\us22/n145 ), .B(\us22/n226 ), .Y(\us22/n223 ) );
  AOI21X1 \us22/U335  ( .A0(\us22/n19 ), .A1(\us22/n223 ), .B0(\us22/n27 ), 
        .Y(\us22/n354 ) );
  AOI31X1 \us22/U334  ( .A0(\us22/n6 ), .A1(\us22/n352 ), .A2(\us22/n259 ), 
        .B0(\us22/n354 ), .Y(\us22/n353 ) );
  OAI221XL \us22/U333  ( .A0(\us22/n20 ), .A1(\us22/n34 ), .B0(\us22/n325 ), 
        .B1(\us22/n4 ), .C0(\us22/n353 ), .Y(\us22/n347 ) );
  INVX1 \us22/U332  ( .A(\us22/n352 ), .Y(\us22/n349 ) );
  NAND2X1 \us22/U331  ( .A(\us22/n278 ), .B(\us22/n6 ), .Y(\us22/n74 ) );
  OAI211X1 \us22/U330  ( .A0(\us22/n349 ), .A1(\us22/n74 ), .B0(\us22/n350 ), 
        .C0(\us22/n351 ), .Y(\us22/n348 ) );
  MXI2X1 \us22/U329  ( .A(\us22/n347 ), .B(\us22/n348 ), .S0(\us22/n252 ), .Y(
        \us22/n332 ) );
  NOR2X1 \us22/U328  ( .A(\us22/n44 ), .B(\us22/n226 ), .Y(\us22/n157 ) );
  INVX1 \us22/U327  ( .A(\us22/n157 ), .Y(\us22/n240 ) );
  NAND2X1 \us22/U326  ( .A(\us22/n240 ), .B(\us22/n189 ), .Y(\us22/n68 ) );
  NOR2X1 \us22/U325  ( .A(\us22/n20 ), .B(\us22/n159 ), .Y(\us22/n225 ) );
  NOR2X1 \us22/U324  ( .A(\us22/n225 ), .B(\us22/n40 ), .Y(\us22/n345 ) );
  INVX1 \us22/U323  ( .A(\us22/n278 ), .Y(\us22/n94 ) );
  NAND2X1 \us22/U322  ( .A(\us22/n94 ), .B(\us22/n226 ), .Y(\us22/n199 ) );
  NAND2X1 \us22/U321  ( .A(\us22/n199 ), .B(\us22/n205 ), .Y(\us22/n82 ) );
  NAND2X1 \us22/U320  ( .A(\us22/n19 ), .B(\us22/n199 ), .Y(\us22/n295 ) );
  NOR2X1 \us22/U319  ( .A(\us22/n226 ), .B(\us22/n259 ), .Y(\us22/n210 ) );
  NOR2X1 \us22/U318  ( .A(\us22/n27 ), .B(\us22/n210 ), .Y(\us22/n173 ) );
  MXI2X1 \us22/U317  ( .A(\us22/n345 ), .B(\us22/n346 ), .S0(\us22/n252 ), .Y(
        \us22/n342 ) );
  NOR2X1 \us22/U316  ( .A(sa22[1]), .B(sa22[3]), .Y(\us22/n163 ) );
  INVX1 \us22/U315  ( .A(\us22/n163 ), .Y(\us22/n37 ) );
  INVX1 \us22/U314  ( .A(\us22/n173 ), .Y(\us22/n344 ) );
  AOI21X1 \us22/U313  ( .A0(\us22/n240 ), .A1(\us22/n37 ), .B0(\us22/n344 ), 
        .Y(\us22/n343 ) );
  AOI211X1 \us22/U312  ( .A0(\us22/n5 ), .A1(\us22/n68 ), .B0(\us22/n342 ), 
        .C0(\us22/n343 ), .Y(\us22/n333 ) );
  NOR2X1 \us22/U311  ( .A(\us22/n18 ), .B(\us22/n226 ), .Y(\us22/n258 ) );
  NAND2X1 \us22/U310  ( .A(\us22/n278 ), .B(sa22[1]), .Y(\us22/n204 ) );
  NOR2X1 \us22/U309  ( .A(\us22/n188 ), .B(sa22[1]), .Y(\us22/n179 ) );
  INVX1 \us22/U308  ( .A(\us22/n179 ), .Y(\us22/n330 ) );
  NAND2X1 \us22/U307  ( .A(\us22/n204 ), .B(\us22/n330 ), .Y(\us22/n239 ) );
  NOR2X1 \us22/U306  ( .A(\us22/n136 ), .B(sa22[1]), .Y(\us22/n299 ) );
  NOR2X1 \us22/U305  ( .A(\us22/n299 ), .B(\us22/n210 ), .Y(\us22/n341 ) );
  OAI32X1 \us22/U304  ( .A0(\us22/n27 ), .A1(\us22/n278 ), .A2(\us22/n95 ), 
        .B0(\us22/n341 ), .B1(\us22/n4 ), .Y(\us22/n340 ) );
  INVX1 \us22/U303  ( .A(\us22/n45 ), .Y(\us22/n126 ) );
  NAND2X1 \us22/U302  ( .A(\us22/n126 ), .B(\us22/n101 ), .Y(\us22/n178 ) );
  NOR2X1 \us22/U301  ( .A(\us22/n18 ), .B(\us22/n136 ), .Y(\us22/n280 ) );
  OAI21XL \us22/U300  ( .A0(\us22/n4 ), .A1(\us22/n121 ), .B0(\us22/n339 ), 
        .Y(\us22/n338 ) );
  MXI2X1 \us22/U299  ( .A(\us22/n336 ), .B(\us22/n337 ), .S0(\us22/n252 ), .Y(
        \us22/n335 ) );
  NOR2X1 \us22/U298  ( .A(\us22/n258 ), .B(\us22/n335 ), .Y(\us22/n334 ) );
  MX4X1 \us22/U297  ( .A(\us22/n331 ), .B(\us22/n332 ), .C(\us22/n333 ), .D(
        \us22/n334 ), .S0(sa22[6]), .S1(\us22/n234 ), .Y(sa20_sr[0]) );
  INVX1 \us22/U296  ( .A(\us22/n299 ), .Y(\us22/n80 ) );
  NOR2X1 \us22/U295  ( .A(\us22/n111 ), .B(\us22/n18 ), .Y(\us22/n269 ) );
  INVX1 \us22/U294  ( .A(\us22/n269 ), .Y(\us22/n75 ) );
  OAI221XL \us22/U293  ( .A0(\us22/n18 ), .A1(\us22/n330 ), .B0(\us22/n20 ), 
        .B1(\us22/n80 ), .C0(\us22/n75 ), .Y(\us22/n329 ) );
  AOI221X1 \us22/U292  ( .A0(\us22/n325 ), .A1(\us22/n33 ), .B0(\us22/n24 ), 
        .B1(\us22/n303 ), .C0(\us22/n329 ), .Y(\us22/n319 ) );
  NOR2X1 \us22/U291  ( .A(\us22/n234 ), .B(sa22[5]), .Y(\us22/n14 ) );
  NOR2X1 \us22/U290  ( .A(\us22/n25 ), .B(\us22/n299 ), .Y(\us22/n313 ) );
  NAND2X1 \us22/U289  ( .A(\us22/n44 ), .B(\us22/n226 ), .Y(\us22/n300 ) );
  AND2X1 \us22/U288  ( .A(\us22/n300 ), .B(\us22/n240 ), .Y(\us22/n23 ) );
  OAI32X1 \us22/U287  ( .A0(\us22/n4 ), .A1(\us22/n145 ), .A2(\us22/n210 ), 
        .B0(\us22/n137 ), .B1(\us22/n27 ), .Y(\us22/n328 ) );
  NOR2X1 \us22/U286  ( .A(sa22[0]), .B(sa22[5]), .Y(\us22/n16 ) );
  INVX1 \us22/U285  ( .A(\us22/n16 ), .Y(\us22/n114 ) );
  INVX1 \us22/U284  ( .A(\us22/n145 ), .Y(\us22/n149 ) );
  NOR2X1 \us22/U283  ( .A(\us22/n47 ), .B(sa22[1]), .Y(\us22/n98 ) );
  INVX1 \us22/U282  ( .A(\us22/n98 ), .Y(\us22/n284 ) );
  OAI21XL \us22/U281  ( .A0(\us22/n69 ), .A1(\us22/n284 ), .B0(\us22/n27 ), 
        .Y(\us22/n327 ) );
  AOI31X1 \us22/U280  ( .A0(\us22/n111 ), .A1(\us22/n149 ), .A2(\us22/n327 ), 
        .B0(\us22/n225 ), .Y(\us22/n326 ) );
  OAI21XL \us22/U279  ( .A0(\us22/n325 ), .A1(\us22/n18 ), .B0(\us22/n326 ), 
        .Y(\us22/n322 ) );
  NAND2X1 \us22/U278  ( .A(\us22/n19 ), .B(\us22/n189 ), .Y(\us22/n71 ) );
  NOR2X1 \us22/U277  ( .A(\us22/n71 ), .B(\us22/n18 ), .Y(\us22/n135 ) );
  AOI21X1 \us22/U276  ( .A0(\us22/n40 ), .A1(sa22[4]), .B0(\us22/n135 ), .Y(
        \us22/n324 ) );
  OAI221XL \us22/U275  ( .A0(\us22/n47 ), .A1(\us22/n27 ), .B0(\us22/n65 ), 
        .B1(\us22/n20 ), .C0(\us22/n324 ), .Y(\us22/n323 ) );
  AOI22X1 \us22/U274  ( .A0(\us22/n55 ), .A1(\us22/n322 ), .B0(\us22/n89 ), 
        .B1(\us22/n323 ), .Y(\us22/n321 ) );
  OAI221XL \us22/U273  ( .A0(\us22/n319 ), .A1(\us22/n52 ), .B0(\us22/n320 ), 
        .B1(\us22/n114 ), .C0(\us22/n321 ), .Y(\us22/n304 ) );
  NOR2X1 \us22/U272  ( .A(\us22/n226 ), .B(\us22/n58 ), .Y(\us22/n290 ) );
  INVX1 \us22/U271  ( .A(\us22/n290 ), .Y(\us22/n200 ) );
  NAND2X1 \us22/U270  ( .A(\us22/n34 ), .B(\us22/n200 ), .Y(\us22/n120 ) );
  INVX1 \us22/U269  ( .A(\us22/n210 ), .Y(\us22/n100 ) );
  OAI221XL \us22/U268  ( .A0(\us22/n20 ), .A1(\us22/n100 ), .B0(sa22[3]), .B1(
        \us22/n4 ), .C0(\us22/n262 ), .Y(\us22/n317 ) );
  INVX1 \us22/U267  ( .A(\us22/n258 ), .Y(\us22/n182 ) );
  AOI211X1 \us22/U266  ( .A0(\us22/n33 ), .A1(\us22/n120 ), .B0(\us22/n317 ), 
        .C0(\us22/n318 ), .Y(\us22/n306 ) );
  NAND2X1 \us22/U265  ( .A(\us22/n100 ), .B(\us22/n199 ), .Y(\us22/n151 ) );
  INVX1 \us22/U264  ( .A(\us22/n151 ), .Y(\us22/n314 ) );
  NOR2X1 \us22/U263  ( .A(\us22/n45 ), .B(\us22/n163 ), .Y(\us22/n160 ) );
  INVX1 \us22/U262  ( .A(\us22/n295 ), .Y(\us22/n92 ) );
  AOI21X1 \us22/U261  ( .A0(sa22[1]), .A1(\us22/n58 ), .B0(\us22/n98 ), .Y(
        \us22/n316 ) );
  OAI22X1 \us22/U260  ( .A0(\us22/n92 ), .A1(\us22/n18 ), .B0(\us22/n316 ), 
        .B1(\us22/n27 ), .Y(\us22/n315 ) );
  NOR2X1 \us22/U259  ( .A(\us22/n149 ), .B(\us22/n226 ), .Y(\us22/n41 ) );
  INVX1 \us22/U258  ( .A(\us22/n41 ), .Y(\us22/n105 ) );
  NAND2X1 \us22/U257  ( .A(\us22/n284 ), .B(\us22/n105 ), .Y(\us22/n227 ) );
  AOI21X1 \us22/U256  ( .A0(\us22/n313 ), .A1(\us22/n33 ), .B0(\us22/n269 ), 
        .Y(\us22/n312 ) );
  OAI221XL \us22/U255  ( .A0(\us22/n149 ), .A1(\us22/n20 ), .B0(\us22/n4 ), 
        .B1(\us22/n227 ), .C0(\us22/n312 ), .Y(\us22/n309 ) );
  AOI21X1 \us22/U254  ( .A0(\us22/n226 ), .A1(\us22/n188 ), .B0(\us22/n242 ), 
        .Y(\us22/n185 ) );
  INVX1 \us22/U253  ( .A(\us22/n185 ), .Y(\us22/n48 ) );
  AND2X1 \us22/U252  ( .A(\us22/n223 ), .B(\us22/n240 ), .Y(\us22/n28 ) );
  OAI221XL \us22/U251  ( .A0(\us22/n27 ), .A1(\us22/n44 ), .B0(\us22/n4 ), 
        .B1(\us22/n48 ), .C0(\us22/n311 ), .Y(\us22/n310 ) );
  AOI22X1 \us22/U250  ( .A0(\us22/n89 ), .A1(\us22/n309 ), .B0(\us22/n55 ), 
        .B1(\us22/n310 ), .Y(\us22/n308 ) );
  OAI221XL \us22/U249  ( .A0(\us22/n306 ), .A1(\us22/n52 ), .B0(\us22/n307 ), 
        .B1(\us22/n114 ), .C0(\us22/n308 ), .Y(\us22/n305 ) );
  MX2X1 \us22/U248  ( .A(\us22/n304 ), .B(\us22/n305 ), .S0(sa22[6]), .Y(
        sa20_sr[1]) );
  INVX1 \us22/U247  ( .A(\us22/n187 ), .Y(\us22/n61 ) );
  MXI2X1 \us22/U246  ( .A(\us22/n303 ), .B(\us22/n61 ), .S0(\us22/n69 ), .Y(
        \us22/n301 ) );
  MXI2X1 \us22/U245  ( .A(\us22/n301 ), .B(\us22/n147 ), .S0(\us22/n302 ), .Y(
        \us22/n285 ) );
  NAND2X1 \us22/U244  ( .A(\us22/n200 ), .B(\us22/n300 ), .Y(\us22/n99 ) );
  INVX1 \us22/U243  ( .A(\us22/n99 ), .Y(\us22/n296 ) );
  NOR2X1 \us22/U242  ( .A(\us22/n299 ), .B(\us22/n242 ), .Y(\us22/n298 ) );
  NAND2X1 \us22/U241  ( .A(sa22[1]), .B(\us22/n47 ), .Y(\us22/n122 ) );
  NOR2X1 \us22/U240  ( .A(\us22/n159 ), .B(\us22/n217 ), .Y(\us22/n198 ) );
  OAI221XL \us22/U239  ( .A0(\us22/n298 ), .A1(\us22/n27 ), .B0(\us22/n20 ), 
        .B1(\us22/n122 ), .C0(\us22/n132 ), .Y(\us22/n297 ) );
  AOI221X1 \us22/U238  ( .A0(\us22/n225 ), .A1(\us22/n226 ), .B0(\us22/n296 ), 
        .B1(\us22/n6 ), .C0(\us22/n297 ), .Y(\us22/n291 ) );
  OAI2BB2X1 \us22/U237  ( .B0(\us22/n27 ), .B1(\us22/n295 ), .A0N(\us22/n34 ), 
        .A1N(\us22/n24 ), .Y(\us22/n293 ) );
  AOI21X1 \us22/U236  ( .A0(\us22/n101 ), .A1(\us22/n150 ), .B0(\us22/n20 ), 
        .Y(\us22/n294 ) );
  AOI211X1 \us22/U235  ( .A0(\us22/n5 ), .A1(\us22/n79 ), .B0(\us22/n293 ), 
        .C0(\us22/n294 ), .Y(\us22/n292 ) );
  INVX1 \us22/U234  ( .A(\us22/n89 ), .Y(\us22/n10 ) );
  OAI22X1 \us22/U233  ( .A0(\us22/n291 ), .A1(\us22/n114 ), .B0(\us22/n292 ), 
        .B1(\us22/n10 ), .Y(\us22/n286 ) );
  INVX1 \us22/U232  ( .A(\us22/n225 ), .Y(\us22/n288 ) );
  NAND2X1 \us22/U231  ( .A(\us22/n200 ), .B(\us22/n284 ), .Y(\us22/n102 ) );
  NOR2X1 \us22/U230  ( .A(\us22/n290 ), .B(\us22/n163 ), .Y(\us22/n184 ) );
  AOI22X1 \us22/U229  ( .A0(\us22/n102 ), .A1(\us22/n69 ), .B0(\us22/n184 ), 
        .B1(\us22/n33 ), .Y(\us22/n289 ) );
  AOI31X1 \us22/U228  ( .A0(\us22/n132 ), .A1(\us22/n288 ), .A2(\us22/n289 ), 
        .B0(\us22/n52 ), .Y(\us22/n287 ) );
  AOI211X1 \us22/U227  ( .A0(\us22/n285 ), .A1(\us22/n55 ), .B0(\us22/n286 ), 
        .C0(\us22/n287 ), .Y(\us22/n263 ) );
  NAND2X1 \us22/U226  ( .A(\us22/n284 ), .B(\us22/n122 ), .Y(\us22/n125 ) );
  NOR2X1 \us22/U225  ( .A(\us22/n199 ), .B(\us22/n4 ), .Y(\us22/n50 ) );
  AOI21X1 \us22/U224  ( .A0(\us22/n200 ), .A1(\us22/n223 ), .B0(\us22/n20 ), 
        .Y(\us22/n283 ) );
  AOI211X1 \us22/U223  ( .A0(\us22/n5 ), .A1(\us22/n125 ), .B0(\us22/n50 ), 
        .C0(\us22/n283 ), .Y(\us22/n282 ) );
  OAI221XL \us22/U222  ( .A0(\us22/n281 ), .A1(\us22/n27 ), .B0(\us22/n4 ), 
        .B1(\us22/n111 ), .C0(\us22/n282 ), .Y(\us22/n265 ) );
  INVX1 \us22/U221  ( .A(\us22/n280 ), .Y(\us22/n247 ) );
  NAND2X1 \us22/U220  ( .A(\us22/n41 ), .B(\us22/n33 ), .Y(\us22/n272 ) );
  OAI221XL \us22/U219  ( .A0(sa22[1]), .A1(\us22/n247 ), .B0(\us22/n4 ), .B1(
        \us22/n189 ), .C0(\us22/n272 ), .Y(\us22/n279 ) );
  NAND2X1 \us22/U218  ( .A(sa22[2]), .B(\us22/n149 ), .Y(\us22/n276 ) );
  XNOR2X1 \us22/U217  ( .A(\us22/n129 ), .B(sa22[1]), .Y(\us22/n155 ) );
  MXI2X1 \us22/U216  ( .A(\us22/n276 ), .B(\us22/n277 ), .S0(\us22/n155 ), .Y(
        \us22/n275 ) );
  OAI22X1 \us22/U215  ( .A0(\us22/n273 ), .A1(\us22/n10 ), .B0(\us22/n274 ), 
        .B1(\us22/n52 ), .Y(\us22/n266 ) );
  NOR2X1 \us22/U214  ( .A(\us22/n20 ), .B(\us22/n226 ), .Y(\us22/n176 ) );
  OAI21XL \us22/U213  ( .A0(\us22/n4 ), .A1(\us22/n271 ), .B0(\us22/n272 ), 
        .Y(\us22/n270 ) );
  OAI31X1 \us22/U212  ( .A0(\us22/n176 ), .A1(\us22/n269 ), .A2(\us22/n270 ), 
        .B0(\us22/n16 ), .Y(\us22/n268 ) );
  INVX1 \us22/U211  ( .A(\us22/n268 ), .Y(\us22/n267 ) );
  AOI211X1 \us22/U210  ( .A0(\us22/n55 ), .A1(\us22/n265 ), .B0(\us22/n266 ), 
        .C0(\us22/n267 ), .Y(\us22/n264 ) );
  MXI2X1 \us22/U209  ( .A(\us22/n263 ), .B(\us22/n264 ), .S0(sa22[6]), .Y(
        sa20_sr[2]) );
  NOR2X1 \us22/U208  ( .A(\us22/n94 ), .B(sa22[1]), .Y(\us22/n211 ) );
  INVX1 \us22/U207  ( .A(\us22/n262 ), .Y(\us22/n261 ) );
  AOI211X1 \us22/U206  ( .A0(\us22/n259 ), .A1(\us22/n24 ), .B0(\us22/n260 ), 
        .C0(\us22/n261 ), .Y(\us22/n255 ) );
  OAI22X1 \us22/U205  ( .A0(\us22/n20 ), .A1(\us22/n68 ), .B0(\us22/n27 ), 
        .B1(\us22/n37 ), .Y(\us22/n257 ) );
  NOR3X1 \us22/U204  ( .A(\us22/n257 ), .B(\us22/n258 ), .C(\us22/n50 ), .Y(
        \us22/n256 ) );
  MXI2X1 \us22/U203  ( .A(\us22/n255 ), .B(\us22/n256 ), .S0(\us22/n252 ), .Y(
        \us22/n254 ) );
  AOI221X1 \us22/U202  ( .A0(\us22/n211 ), .A1(\us22/n5 ), .B0(\us22/n40 ), 
        .B1(sa22[4]), .C0(\us22/n254 ), .Y(\us22/n248 ) );
  INVX1 \us22/U201  ( .A(\us22/n211 ), .Y(\us22/n106 ) );
  NAND2X1 \us22/U200  ( .A(\us22/n200 ), .B(\us22/n106 ), .Y(\us22/n83 ) );
  NAND2X1 \us22/U199  ( .A(\us22/n199 ), .B(\us22/n204 ), .Y(\us22/n169 ) );
  AOI2BB2X1 \us22/U198  ( .B0(\us22/n65 ), .B1(\us22/n24 ), .A0N(\us22/n169 ), 
        .A1N(\us22/n20 ), .Y(\us22/n253 ) );
  OAI221XL \us22/U197  ( .A0(\us22/n172 ), .A1(\us22/n18 ), .B0(\us22/n27 ), 
        .B1(\us22/n83 ), .C0(\us22/n253 ), .Y(\us22/n251 ) );
  MXI2X1 \us22/U196  ( .A(\us22/n250 ), .B(\us22/n251 ), .S0(\us22/n252 ), .Y(
        \us22/n249 ) );
  MXI2X1 \us22/U195  ( .A(\us22/n248 ), .B(\us22/n249 ), .S0(\us22/n234 ), .Y(
        \us22/n228 ) );
  OAI21XL \us22/U194  ( .A0(\us22/n58 ), .A1(\us22/n27 ), .B0(\us22/n247 ), 
        .Y(\us22/n245 ) );
  NOR2X1 \us22/U193  ( .A(sa22[7]), .B(\us22/n145 ), .Y(\us22/n246 ) );
  XNOR2X1 \us22/U192  ( .A(\us22/n69 ), .B(sa22[1]), .Y(\us22/n130 ) );
  MXI2X1 \us22/U191  ( .A(\us22/n245 ), .B(\us22/n246 ), .S0(\us22/n130 ), .Y(
        \us22/n243 ) );
  OAI211X1 \us22/U190  ( .A0(\us22/n4 ), .A1(\us22/n149 ), .B0(\us22/n243 ), 
        .C0(\us22/n244 ), .Y(\us22/n230 ) );
  NOR2X1 \us22/U189  ( .A(\us22/n242 ), .B(\us22/n137 ), .Y(\us22/n70 ) );
  OAI221XL \us22/U188  ( .A0(\us22/n159 ), .A1(\us22/n27 ), .B0(\us22/n20 ), 
        .B1(\us22/n34 ), .C0(\us22/n241 ), .Y(\us22/n231 ) );
  NAND2X1 \us22/U187  ( .A(\us22/n101 ), .B(\us22/n240 ), .Y(\us22/n76 ) );
  AOI21X1 \us22/U186  ( .A0(\us22/n122 ), .A1(\us22/n106 ), .B0(\us22/n129 ), 
        .Y(\us22/n237 ) );
  INVX1 \us22/U185  ( .A(\us22/n239 ), .Y(\us22/n238 ) );
  OAI21XL \us22/U184  ( .A0(\us22/n237 ), .A1(\us22/n43 ), .B0(\us22/n238 ), 
        .Y(\us22/n236 ) );
  OAI221XL \us22/U183  ( .A0(\us22/n18 ), .A1(\us22/n76 ), .B0(\us22/n59 ), 
        .B1(\us22/n27 ), .C0(\us22/n236 ), .Y(\us22/n232 ) );
  AOI2BB2X1 \us22/U182  ( .B0(\us22/n24 ), .B1(\us22/n187 ), .A0N(\us22/n227 ), 
        .A1N(\us22/n20 ), .Y(\us22/n235 ) );
  OAI211X1 \us22/U181  ( .A0(\us22/n27 ), .A1(\us22/n122 ), .B0(\us22/n158 ), 
        .C0(\us22/n235 ), .Y(\us22/n233 ) );
  MX4X1 \us22/U180  ( .A(\us22/n230 ), .B(\us22/n231 ), .C(\us22/n232 ), .D(
        \us22/n233 ), .S0(\us22/n234 ), .S1(sa22[5]), .Y(\us22/n229 ) );
  MX2X1 \us22/U179  ( .A(\us22/n228 ), .B(\us22/n229 ), .S0(sa22[6]), .Y(
        sa20_sr[3]) );
  NOR2BX1 \us22/U178  ( .AN(\us22/n204 ), .B(\us22/n137 ), .Y(\us22/n110 ) );
  INVX1 \us22/U177  ( .A(\us22/n110 ), .Y(\us22/n64 ) );
  AOI22X1 \us22/U176  ( .A0(\us22/n225 ), .A1(\us22/n226 ), .B0(\us22/n6 ), 
        .B1(\us22/n227 ), .Y(\us22/n224 ) );
  OAI221XL \us22/U175  ( .A0(\us22/n27 ), .A1(\us22/n64 ), .B0(\us22/n4 ), 
        .B1(\us22/n83 ), .C0(\us22/n224 ), .Y(\us22/n212 ) );
  NAND2X1 \us22/U174  ( .A(\us22/n34 ), .B(\us22/n204 ), .Y(\us22/n221 ) );
  OAI21XL \us22/U173  ( .A0(\us22/n69 ), .A1(\us22/n223 ), .B0(\us22/n27 ), 
        .Y(\us22/n222 ) );
  NOR2X1 \us22/U172  ( .A(\us22/n217 ), .B(\us22/n42 ), .Y(\us22/n208 ) );
  AOI211X1 \us22/U171  ( .A0(\us22/n208 ), .A1(\us22/n5 ), .B0(\us22/n220 ), 
        .C0(\us22/n173 ), .Y(\us22/n219 ) );
  OAI22X1 \us22/U170  ( .A0(\us22/n218 ), .A1(\us22/n10 ), .B0(\us22/n219 ), 
        .B1(\us22/n114 ), .Y(\us22/n213 ) );
  INVX1 \us22/U169  ( .A(\us22/n135 ), .Y(\us22/n215 ) );
  NOR2X1 \us22/U168  ( .A(\us22/n4 ), .B(\us22/n159 ), .Y(\us22/n31 ) );
  INVX1 \us22/U167  ( .A(\us22/n31 ), .Y(\us22/n196 ) );
  AOI31X1 \us22/U166  ( .A0(\us22/n215 ), .A1(\us22/n196 ), .A2(\us22/n216 ), 
        .B0(\us22/n52 ), .Y(\us22/n214 ) );
  AOI211X1 \us22/U165  ( .A0(\us22/n55 ), .A1(\us22/n212 ), .B0(\us22/n213 ), 
        .C0(\us22/n214 ), .Y(\us22/n190 ) );
  INVX1 \us22/U164  ( .A(\us22/n207 ), .Y(\us22/n192 ) );
  NOR2X1 \us22/U163  ( .A(\us22/n25 ), .B(\us22/n98 ), .Y(\us22/n32 ) );
  OAI22X1 \us22/U162  ( .A0(\us22/n28 ), .A1(\us22/n4 ), .B0(\us22/n188 ), 
        .B1(\us22/n27 ), .Y(\us22/n206 ) );
  NAND2X1 \us22/U161  ( .A(\us22/n204 ), .B(\us22/n80 ), .Y(\us22/n118 ) );
  INVX1 \us22/U160  ( .A(\us22/n118 ), .Y(\us22/n123 ) );
  NAND2X1 \us22/U159  ( .A(\us22/n94 ), .B(\us22/n79 ), .Y(\us22/n203 ) );
  OAI2BB1X1 \us22/U158  ( .A0N(\us22/n199 ), .A1N(\us22/n200 ), .B0(\us22/n33 ), .Y(\us22/n195 ) );
  INVX1 \us22/U157  ( .A(\us22/n55 ), .Y(\us22/n12 ) );
  AOI31X1 \us22/U156  ( .A0(\us22/n195 ), .A1(\us22/n196 ), .A2(\us22/n197 ), 
        .B0(\us22/n12 ), .Y(\us22/n194 ) );
  AOI211X1 \us22/U155  ( .A0(\us22/n89 ), .A1(\us22/n192 ), .B0(\us22/n193 ), 
        .C0(\us22/n194 ), .Y(\us22/n191 ) );
  MXI2X1 \us22/U154  ( .A(\us22/n190 ), .B(\us22/n191 ), .S0(sa22[6]), .Y(
        sa20_sr[4]) );
  OAI21XL \us22/U153  ( .A0(\us22/n69 ), .A1(\us22/n189 ), .B0(\us22/n27 ), 
        .Y(\us22/n186 ) );
  INVX1 \us22/U152  ( .A(\us22/n183 ), .Y(\us22/n180 ) );
  NAND2X1 \us22/U151  ( .A(\us22/n74 ), .B(\us22/n182 ), .Y(\us22/n181 ) );
  AOI211X1 \us22/U150  ( .A0(\us22/n179 ), .A1(\us22/n24 ), .B0(\us22/n180 ), 
        .C0(\us22/n181 ), .Y(\us22/n165 ) );
  INVX1 \us22/U149  ( .A(\us22/n178 ), .Y(\us22/n175 ) );
  AOI211X1 \us22/U148  ( .A0(\us22/n175 ), .A1(\us22/n5 ), .B0(\us22/n176 ), 
        .C0(\us22/n177 ), .Y(\us22/n174 ) );
  OAI221XL \us22/U147  ( .A0(\us22/n159 ), .A1(\us22/n27 ), .B0(\us22/n145 ), 
        .B1(\us22/n20 ), .C0(\us22/n174 ), .Y(\us22/n167 ) );
  MXI2X1 \us22/U146  ( .A(\us22/n40 ), .B(\us22/n173 ), .S0(\us22/n96 ), .Y(
        \us22/n170 ) );
  AOI22X1 \us22/U145  ( .A0(\us22/n137 ), .A1(\us22/n24 ), .B0(\us22/n172 ), 
        .B1(\us22/n6 ), .Y(\us22/n171 ) );
  OAI211X1 \us22/U144  ( .A0(\us22/n20 ), .A1(\us22/n169 ), .B0(\us22/n170 ), 
        .C0(\us22/n171 ), .Y(\us22/n168 ) );
  AOI22X1 \us22/U143  ( .A0(\us22/n89 ), .A1(\us22/n167 ), .B0(\us22/n55 ), 
        .B1(\us22/n168 ), .Y(\us22/n166 ) );
  OAI221XL \us22/U142  ( .A0(\us22/n164 ), .A1(\us22/n114 ), .B0(\us22/n165 ), 
        .B1(\us22/n52 ), .C0(\us22/n166 ), .Y(\us22/n138 ) );
  OAI21XL \us22/U141  ( .A0(\us22/n41 ), .A1(\us22/n163 ), .B0(\us22/n69 ), 
        .Y(\us22/n162 ) );
  AOI221X1 \us22/U140  ( .A0(\us22/n159 ), .A1(\us22/n24 ), .B0(\us22/n160 ), 
        .B1(\us22/n33 ), .C0(\us22/n161 ), .Y(\us22/n140 ) );
  OAI21XL \us22/U139  ( .A0(\us22/n157 ), .A1(\us22/n20 ), .B0(\us22/n158 ), 
        .Y(\us22/n156 ) );
  NOR2X1 \us22/U138  ( .A(\us22/n4 ), .B(\us22/n136 ), .Y(\us22/n153 ) );
  NOR2X1 \us22/U137  ( .A(\us22/n145 ), .B(\us22/n69 ), .Y(\us22/n154 ) );
  MXI2X1 \us22/U136  ( .A(\us22/n153 ), .B(\us22/n154 ), .S0(\us22/n155 ), .Y(
        \us22/n152 ) );
  OAI221XL \us22/U135  ( .A0(\us22/n110 ), .A1(\us22/n18 ), .B0(\us22/n20 ), 
        .B1(\us22/n151 ), .C0(\us22/n152 ), .Y(\us22/n143 ) );
  AOI21X1 \us22/U134  ( .A0(\us22/n149 ), .A1(\us22/n150 ), .B0(\us22/n18 ), 
        .Y(\us22/n148 ) );
  AOI2BB1X1 \us22/U133  ( .A0N(\us22/n147 ), .A1N(\us22/n27 ), .B0(\us22/n148 ), .Y(\us22/n146 ) );
  OAI221XL \us22/U132  ( .A0(\us22/n145 ), .A1(\us22/n20 ), .B0(\us22/n4 ), 
        .B1(\us22/n34 ), .C0(\us22/n146 ), .Y(\us22/n144 ) );
  AOI22X1 \us22/U131  ( .A0(\us22/n89 ), .A1(\us22/n143 ), .B0(\us22/n14 ), 
        .B1(\us22/n144 ), .Y(\us22/n142 ) );
  OAI221XL \us22/U130  ( .A0(\us22/n140 ), .A1(\us22/n12 ), .B0(\us22/n141 ), 
        .B1(\us22/n114 ), .C0(\us22/n142 ), .Y(\us22/n139 ) );
  MX2X1 \us22/U129  ( .A(\us22/n138 ), .B(\us22/n139 ), .S0(sa22[6]), .Y(
        sa20_sr[5]) );
  INVX1 \us22/U128  ( .A(\us22/n70 ), .Y(\us22/n133 ) );
  OAI22X1 \us22/U127  ( .A0(\us22/n4 ), .A1(\us22/n136 ), .B0(\us22/n137 ), 
        .B1(\us22/n27 ), .Y(\us22/n134 ) );
  AOI211X1 \us22/U126  ( .A0(\us22/n133 ), .A1(\us22/n69 ), .B0(\us22/n134 ), 
        .C0(\us22/n135 ), .Y(\us22/n112 ) );
  INVX1 \us22/U125  ( .A(\us22/n132 ), .Y(\us22/n131 ) );
  OAI21XL \us22/U124  ( .A0(\us22/n18 ), .A1(\us22/n37 ), .B0(\us22/n128 ), 
        .Y(\us22/n127 ) );
  OAI221XL \us22/U123  ( .A0(\us22/n18 ), .A1(\us22/n105 ), .B0(\us22/n123 ), 
        .B1(\us22/n27 ), .C0(\us22/n124 ), .Y(\us22/n116 ) );
  NAND2X1 \us22/U122  ( .A(\us22/n121 ), .B(\us22/n122 ), .Y(\us22/n30 ) );
  OAI221XL \us22/U121  ( .A0(\us22/n18 ), .A1(\us22/n118 ), .B0(\us22/n27 ), 
        .B1(\us22/n30 ), .C0(\us22/n119 ), .Y(\us22/n117 ) );
  AOI22X1 \us22/U120  ( .A0(\us22/n89 ), .A1(\us22/n116 ), .B0(\us22/n55 ), 
        .B1(\us22/n117 ), .Y(\us22/n115 ) );
  OAI221XL \us22/U119  ( .A0(\us22/n112 ), .A1(\us22/n52 ), .B0(\us22/n113 ), 
        .B1(\us22/n114 ), .C0(\us22/n115 ), .Y(\us22/n84 ) );
  OAI22X1 \us22/U118  ( .A0(\us22/n110 ), .A1(\us22/n4 ), .B0(\us22/n20 ), 
        .B1(\us22/n21 ), .Y(\us22/n108 ) );
  AOI21X1 \us22/U117  ( .A0(sa22[1]), .A1(\us22/n58 ), .B0(\us22/n27 ), .Y(
        \us22/n109 ) );
  AOI211X1 \us22/U116  ( .A0(\us22/n5 ), .A1(\us22/n107 ), .B0(\us22/n108 ), 
        .C0(\us22/n109 ), .Y(\us22/n86 ) );
  OAI22X1 \us22/U115  ( .A0(\us22/n45 ), .A1(\us22/n4 ), .B0(sa22[4]), .B1(
        \us22/n18 ), .Y(\us22/n103 ) );
  AOI21X1 \us22/U114  ( .A0(\us22/n105 ), .A1(\us22/n106 ), .B0(\us22/n20 ), 
        .Y(\us22/n104 ) );
  AOI211X1 \us22/U113  ( .A0(\us22/n33 ), .A1(\us22/n102 ), .B0(\us22/n103 ), 
        .C0(\us22/n104 ), .Y(\us22/n87 ) );
  NAND2X1 \us22/U112  ( .A(\us22/n100 ), .B(\us22/n101 ), .Y(\us22/n62 ) );
  OAI221XL \us22/U111  ( .A0(\us22/n27 ), .A1(\us22/n62 ), .B0(\us22/n4 ), 
        .B1(\us22/n21 ), .C0(\us22/n97 ), .Y(\us22/n90 ) );
  NOR3X1 \us22/U110  ( .A(\us22/n4 ), .B(\us22/n95 ), .C(\us22/n96 ), .Y(
        \us22/n67 ) );
  AOI31X1 \us22/U109  ( .A0(\us22/n79 ), .A1(\us22/n94 ), .A2(\us22/n6 ), .B0(
        \us22/n67 ), .Y(\us22/n93 ) );
  OAI221XL \us22/U108  ( .A0(\us22/n73 ), .A1(\us22/n27 ), .B0(\us22/n92 ), 
        .B1(\us22/n20 ), .C0(\us22/n93 ), .Y(\us22/n91 ) );
  AOI22X1 \us22/U107  ( .A0(\us22/n89 ), .A1(\us22/n90 ), .B0(\us22/n16 ), 
        .B1(\us22/n91 ), .Y(\us22/n88 ) );
  OAI221XL \us22/U106  ( .A0(\us22/n86 ), .A1(\us22/n52 ), .B0(\us22/n87 ), 
        .B1(\us22/n12 ), .C0(\us22/n88 ), .Y(\us22/n85 ) );
  MX2X1 \us22/U105  ( .A(\us22/n84 ), .B(\us22/n85 ), .S0(sa22[6]), .Y(
        sa20_sr[6]) );
  INVX1 \us22/U104  ( .A(\us22/n81 ), .Y(\us22/n77 ) );
  AOI21X1 \us22/U103  ( .A0(\us22/n79 ), .A1(\us22/n80 ), .B0(\us22/n27 ), .Y(
        \us22/n78 ) );
  AOI211X1 \us22/U102  ( .A0(\us22/n5 ), .A1(\us22/n76 ), .B0(\us22/n77 ), 
        .C0(\us22/n78 ), .Y(\us22/n51 ) );
  OAI211X1 \us22/U101  ( .A0(\us22/n73 ), .A1(\us22/n27 ), .B0(\us22/n74 ), 
        .C0(\us22/n75 ), .Y(\us22/n72 ) );
  AOI21X1 \us22/U100  ( .A0(\us22/n68 ), .A1(\us22/n69 ), .B0(\us22/n6 ), .Y(
        \us22/n63 ) );
  INVX1 \us22/U99  ( .A(\us22/n67 ), .Y(\us22/n66 ) );
  OAI221XL \us22/U98  ( .A0(\us22/n63 ), .A1(\us22/n64 ), .B0(\us22/n65 ), 
        .B1(\us22/n27 ), .C0(\us22/n66 ), .Y(\us22/n56 ) );
  AOI2BB2X1 \us22/U97  ( .B0(\us22/n61 ), .B1(\us22/n24 ), .A0N(\us22/n62 ), 
        .A1N(\us22/n20 ), .Y(\us22/n60 ) );
  OAI221XL \us22/U96  ( .A0(\us22/n58 ), .A1(\us22/n18 ), .B0(\us22/n59 ), 
        .B1(\us22/n27 ), .C0(\us22/n60 ), .Y(\us22/n57 ) );
  AOI22X1 \us22/U95  ( .A0(\us22/n55 ), .A1(\us22/n56 ), .B0(\us22/n16 ), .B1(
        \us22/n57 ), .Y(\us22/n54 ) );
  OAI221XL \us22/U94  ( .A0(\us22/n51 ), .A1(\us22/n52 ), .B0(\us22/n53 ), 
        .B1(\us22/n10 ), .C0(\us22/n54 ), .Y(\us22/n7 ) );
  INVX1 \us22/U93  ( .A(\us22/n50 ), .Y(\us22/n49 ) );
  OAI221XL \us22/U92  ( .A0(\us22/n47 ), .A1(\us22/n18 ), .B0(\us22/n27 ), 
        .B1(\us22/n48 ), .C0(\us22/n49 ), .Y(\us22/n46 ) );
  NOR2X1 \us22/U91  ( .A(\us22/n41 ), .B(\us22/n42 ), .Y(\us22/n38 ) );
  INVX1 \us22/U90  ( .A(\us22/n40 ), .Y(\us22/n39 ) );
  INVX1 \us22/U89  ( .A(\us22/n32 ), .Y(\us22/n26 ) );
  AOI21X1 \us22/U88  ( .A0(\us22/n5 ), .A1(\us22/n30 ), .B0(\us22/n31 ), .Y(
        \us22/n29 ) );
  OAI221XL \us22/U87  ( .A0(\us22/n26 ), .A1(\us22/n27 ), .B0(\us22/n28 ), 
        .B1(\us22/n20 ), .C0(\us22/n29 ), .Y(\us22/n15 ) );
  OAI221XL \us22/U86  ( .A0(\us22/n18 ), .A1(\us22/n19 ), .B0(\us22/n20 ), 
        .B1(\us22/n21 ), .C0(\us22/n22 ), .Y(\us22/n17 ) );
  AOI22X1 \us22/U85  ( .A0(\us22/n14 ), .A1(\us22/n15 ), .B0(\us22/n16 ), .B1(
        \us22/n17 ), .Y(\us22/n13 ) );
  OAI221XL \us22/U84  ( .A0(\us22/n9 ), .A1(\us22/n10 ), .B0(\us22/n11 ), .B1(
        \us22/n12 ), .C0(\us22/n13 ), .Y(\us22/n8 ) );
  MX2X1 \us22/U83  ( .A(\us22/n7 ), .B(\us22/n8 ), .S0(sa22[6]), .Y(sa20_sr[7]) );
  NOR2X4 \us22/U82  ( .A(\us22/n129 ), .B(sa22[2]), .Y(\us22/n43 ) );
  CLKINVX3 \us22/U81  ( .A(\us22/n14 ), .Y(\us22/n52 ) );
  OAI22XL \us22/U80  ( .A0(\us22/n201 ), .A1(\us22/n52 ), .B0(\us22/n202 ), 
        .B1(\us22/n114 ), .Y(\us22/n193 ) );
  CLKINVX3 \us22/U79  ( .A(sa22[5]), .Y(\us22/n252 ) );
  NOR2X2 \us22/U78  ( .A(\us22/n252 ), .B(\us22/n234 ), .Y(\us22/n55 ) );
  CLKINVX3 \us22/U77  ( .A(sa22[7]), .Y(\us22/n129 ) );
  NOR2X4 \us22/U76  ( .A(\us22/n129 ), .B(\us22/n69 ), .Y(\us22/n24 ) );
  AOI22XL \us22/U75  ( .A0(\us22/n70 ), .A1(\us22/n24 ), .B0(\us22/n96 ), .B1(
        \us22/n129 ), .Y(\us22/n241 ) );
  NOR2X2 \us22/U74  ( .A(\us22/n252 ), .B(sa22[0]), .Y(\us22/n89 ) );
  CLKINVX3 \us22/U73  ( .A(sa22[0]), .Y(\us22/n234 ) );
  NOR2X4 \us22/U72  ( .A(\us22/n69 ), .B(sa22[7]), .Y(\us22/n33 ) );
  INVX12 \us22/U71  ( .A(\us22/n33 ), .Y(\us22/n27 ) );
  CLKINVX3 \us22/U70  ( .A(\us22/n1 ), .Y(\us22/n6 ) );
  CLKINVX3 \us22/U69  ( .A(\us22/n1 ), .Y(\us22/n5 ) );
  INVXL \us22/U68  ( .A(\us22/n24 ), .Y(\us22/n36 ) );
  INVX4 \us22/U67  ( .A(\us22/n3 ), .Y(\us22/n4 ) );
  INVXL \us22/U66  ( .A(\us22/n36 ), .Y(\us22/n3 ) );
  INVX4 \us22/U65  ( .A(sa22[1]), .Y(\us22/n226 ) );
  INVX4 \us22/U64  ( .A(\us22/n43 ), .Y(\us22/n20 ) );
  AOI221X4 \us22/U63  ( .A0(\us22/n24 ), .A1(\us22/n82 ), .B0(\us22/n43 ), 
        .B1(\us22/n295 ), .C0(\us22/n173 ), .Y(\us22/n346 ) );
  AOI221X4 \us22/U62  ( .A0(\us22/n5 ), .A1(\us22/n96 ), .B0(\us22/n43 ), .B1(
        \us22/n239 ), .C0(\us22/n340 ), .Y(\us22/n336 ) );
  AOI222X4 \us22/U61  ( .A0(\us22/n59 ), .A1(\us22/n43 ), .B0(\us22/n6 ), .B1(
        \us22/n221 ), .C0(\us22/n222 ), .C1(\us22/n187 ), .Y(\us22/n218 ) );
  AOI222X4 \us22/U60  ( .A0(\us22/n123 ), .A1(\us22/n43 ), .B0(sa22[2]), .B1(
        \us22/n203 ), .C0(\us22/n6 ), .C1(\us22/n71 ), .Y(\us22/n202 ) );
  AOI221X4 \us22/U59  ( .A0(\us22/n314 ), .A1(\us22/n43 ), .B0(\us22/n160 ), 
        .B1(\us22/n24 ), .C0(\us22/n315 ), .Y(\us22/n307 ) );
  AOI221X4 \us22/U58  ( .A0(\us22/n43 ), .A1(\us22/n208 ), .B0(\us22/n76 ), 
        .B1(\us22/n24 ), .C0(\us22/n209 ), .Y(\us22/n207 ) );
  AOI221X4 \us22/U57  ( .A0(\us22/n43 ), .A1(\us22/n205 ), .B0(\us22/n32 ), 
        .B1(\us22/n6 ), .C0(\us22/n206 ), .Y(\us22/n201 ) );
  AOI221X4 \us22/U56  ( .A0(\us22/n43 ), .A1(\us22/n44 ), .B0(\us22/n45 ), 
        .B1(\us22/n24 ), .C0(\us22/n46 ), .Y(\us22/n9 ) );
  AOI22XL \us22/U55  ( .A0(\us22/n217 ), .A1(\us22/n43 ), .B0(\us22/n33 ), 
        .B1(\us22/n47 ), .Y(\us22/n216 ) );
  AOI22XL \us22/U54  ( .A0(\us22/n98 ), .A1(\us22/n43 ), .B0(\us22/n6 ), .B1(
        \us22/n99 ), .Y(\us22/n97 ) );
  AOI22XL \us22/U53  ( .A0(\us22/n82 ), .A1(\us22/n43 ), .B0(\us22/n83 ), .B1(
        \us22/n24 ), .Y(\us22/n81 ) );
  AOI2BB2XL \us22/U52  ( .B0(\us22/n43 ), .B1(\us22/n94 ), .A0N(\us22/n120 ), 
        .A1N(\us22/n4 ), .Y(\us22/n119 ) );
  AOI222X4 \us22/U51  ( .A0(\us22/n125 ), .A1(\us22/n33 ), .B0(\us22/n145 ), 
        .B1(\us22/n40 ), .C0(\us22/n43 ), .C1(\us22/n184 ), .Y(\us22/n183 ) );
  AOI22XL \us22/U50  ( .A0(\us22/n43 ), .A1(\us22/n303 ), .B0(\us22/n24 ), 
        .B1(\us22/n96 ), .Y(\us22/n358 ) );
  AOI22XL \us22/U49  ( .A0(\us22/n43 ), .A1(\us22/n100 ), .B0(\us22/n24 ), 
        .B1(\us22/n125 ), .Y(\us22/n124 ) );
  AOI21XL \us22/U48  ( .A0(\us22/n159 ), .A1(\us22/n43 ), .B0(\us22/n40 ), .Y(
        \us22/n262 ) );
  AOI22XL \us22/U47  ( .A0(\us22/n40 ), .A1(\us22/n94 ), .B0(\us22/n43 ), .B1(
        \us22/n187 ), .Y(\us22/n244 ) );
  AOI22XL \us22/U46  ( .A0(\us22/n184 ), .A1(\us22/n5 ), .B0(\us22/n198 ), 
        .B1(\us22/n43 ), .Y(\us22/n197 ) );
  NOR2XL \us22/U45  ( .A(\us22/n33 ), .B(\us22/n2 ), .Y(\us22/n302 ) );
  MXI2XL \us22/U44  ( .A(\us22/n2 ), .B(\us22/n6 ), .S0(\us22/n28 ), .Y(
        \us22/n311 ) );
  INVXL \us22/U43  ( .A(\us22/n20 ), .Y(\us22/n2 ) );
  INVX4 \us22/U42  ( .A(\us22/n6 ), .Y(\us22/n18 ) );
  AOI21XL \us22/U41  ( .A0(\us22/n18 ), .A1(\us22/n162 ), .B0(\us22/n25 ), .Y(
        \us22/n161 ) );
  INVX4 \us22/U40  ( .A(sa22[2]), .Y(\us22/n69 ) );
  NOR2X4 \us22/U39  ( .A(\us22/n226 ), .B(\us22/n4 ), .Y(\us22/n40 ) );
  CLKINVX3 \us22/U38  ( .A(sa22[3]), .Y(\us22/n136 ) );
  NOR2X2 \us22/U37  ( .A(\us22/n136 ), .B(sa22[4]), .Y(\us22/n145 ) );
  CLKINVX3 \us22/U36  ( .A(sa22[4]), .Y(\us22/n58 ) );
  NOR2X2 \us22/U35  ( .A(\us22/n58 ), .B(sa22[3]), .Y(\us22/n159 ) );
  NOR2X2 \us22/U34  ( .A(\us22/n136 ), .B(\us22/n58 ), .Y(\us22/n259 ) );
  NOR2X2 \us22/U33  ( .A(sa22[4]), .B(sa22[3]), .Y(\us22/n278 ) );
  NOR2X2 \us22/U32  ( .A(\us22/n259 ), .B(\us22/n278 ), .Y(\us22/n47 ) );
  CLKINVX3 \us22/U31  ( .A(\us22/n259 ), .Y(\us22/n44 ) );
  NOR2X2 \us22/U30  ( .A(\us22/n44 ), .B(sa22[1]), .Y(\us22/n137 ) );
  AOI21XL \us22/U29  ( .A0(\us22/n44 ), .A1(\us22/n111 ), .B0(\us22/n4 ), .Y(
        \us22/n177 ) );
  AOI22XL \us22/U28  ( .A0(\us22/n23 ), .A1(\us22/n24 ), .B0(\us22/n25 ), .B1(
        sa22[2]), .Y(\us22/n22 ) );
  AOI22XL \us22/U27  ( .A0(\us22/n33 ), .A1(sa22[3]), .B0(\us22/n24 ), .B1(
        \us22/n58 ), .Y(\us22/n277 ) );
  NAND2XL \us22/U26  ( .A(\us22/n198 ), .B(\us22/n24 ), .Y(\us22/n132 ) );
  OAI2BB2XL \us22/U25  ( .B0(\us22/n20 ), .B1(\us22/n111 ), .A0N(\us22/n125 ), 
        .A1N(\us22/n24 ), .Y(\us22/n220 ) );
  NAND2XL \us22/U24  ( .A(\us22/n111 ), .B(\us22/n101 ), .Y(\us22/n21 ) );
  NAND2XL \us22/U23  ( .A(\us22/n111 ), .B(\us22/n300 ), .Y(\us22/n187 ) );
  NAND2XL \us22/U22  ( .A(\us22/n111 ), .B(\us22/n121 ), .Y(\us22/n303 ) );
  AOI221XL \us22/U21  ( .A0(\us22/n43 ), .A1(\us22/n151 ), .B0(\us22/n25 ), 
        .B1(\us22/n69 ), .C0(\us22/n275 ), .Y(\us22/n274 ) );
  NOR2BXL \us22/U20  ( .AN(\us22/n101 ), .B(\us22/n25 ), .Y(\us22/n172 ) );
  NAND2X2 \us22/U19  ( .A(\us22/n58 ), .B(\us22/n226 ), .Y(\us22/n34 ) );
  OAI222X1 \us22/U18  ( .A0(\us22/n27 ), .A1(\us22/n34 ), .B0(\us22/n69 ), 
        .B1(\us22/n205 ), .C0(\us22/n20 ), .C1(\us22/n79 ), .Y(\us22/n260 ) );
  OAI222X1 \us22/U17  ( .A0(\us22/n20 ), .A1(\us22/n99 ), .B0(\us22/n27 ), 
        .B1(\us22/n101 ), .C0(\us22/n184 ), .C1(\us22/n4 ), .Y(\us22/n250 ) );
  OAI222X1 \us22/U16  ( .A0(\us22/n4 ), .A1(\us22/n37 ), .B0(\us22/n38 ), .B1(
        \us22/n20 ), .C0(sa22[4]), .C1(\us22/n39 ), .Y(\us22/n35 ) );
  AOI221X1 \us22/U15  ( .A0(\us22/n5 ), .A1(\us22/n19 ), .B0(\us22/n33 ), .B1(
        \us22/n34 ), .C0(\us22/n35 ), .Y(\us22/n11 ) );
  OR2X2 \us22/U14  ( .A(sa22[2]), .B(sa22[7]), .Y(\us22/n1 ) );
  AOI221XL \us22/U13  ( .A0(\us22/n59 ), .A1(\us22/n33 ), .B0(\us22/n43 ), 
        .B1(\us22/n126 ), .C0(\us22/n127 ), .Y(\us22/n113 ) );
  AOI221XL \us22/U12  ( .A0(\us22/n70 ), .A1(\us22/n43 ), .B0(\us22/n24 ), 
        .B1(\us22/n71 ), .C0(\us22/n72 ), .Y(\us22/n53 ) );
  AOI221X1 \us22/U11  ( .A0(\us22/n313 ), .A1(\us22/n5 ), .B0(\us22/n23 ), 
        .B1(\us22/n2 ), .C0(\us22/n328 ), .Y(\us22/n320 ) );
  AOI222XL \us22/U10  ( .A0(\us22/n185 ), .A1(\us22/n43 ), .B0(\us22/n186 ), 
        .B1(\us22/n187 ), .C0(\us22/n6 ), .C1(\us22/n188 ), .Y(\us22/n164 ) );
  AOI221X1 \us22/U9  ( .A0(\us22/n40 ), .A1(\us22/n136 ), .B0(\us22/n33 ), 
        .B1(\us22/n178 ), .C0(\us22/n338 ), .Y(\us22/n337 ) );
  AOI222XL \us22/U8  ( .A0(\us22/n278 ), .A1(\us22/n24 ), .B0(\us22/n42 ), 
        .B1(\us22/n33 ), .C0(\us22/n43 ), .C1(\us22/n136 ), .Y(\us22/n351 ) );
  AOI31X1 \us22/U7  ( .A0(sa22[2]), .A1(\us22/n58 ), .A2(sa22[1]), .B0(
        \us22/n40 ), .Y(\us22/n350 ) );
  AOI31X1 \us22/U6  ( .A0(\us22/n44 ), .A1(\us22/n129 ), .A2(\us22/n130 ), 
        .B0(\us22/n131 ), .Y(\us22/n128 ) );
  OAI32X1 \us22/U5  ( .A0(\us22/n18 ), .A1(sa22[1]), .A2(\us22/n159 ), .B0(
        sa22[4]), .B1(\us22/n182 ), .Y(\us22/n318 ) );
  AOI221X1 \us22/U4  ( .A0(\us22/n278 ), .A1(\us22/n40 ), .B0(\us22/n185 ), 
        .B1(\us22/n2 ), .C0(\us22/n279 ), .Y(\us22/n273 ) );
  AOI221X1 \us22/U3  ( .A0(\us22/n40 ), .A1(\us22/n136 ), .B0(\us22/n33 ), 
        .B1(\us22/n47 ), .C0(\us22/n156 ), .Y(\us22/n141 ) );
  OAI32X1 \us22/U2  ( .A0(\us22/n210 ), .A1(\us22/n145 ), .A2(\us22/n18 ), 
        .B0(\us22/n27 ), .B1(\us22/n211 ), .Y(\us22/n209 ) );
  AOI31XL \us22/U1  ( .A0(\us22/n79 ), .A1(\us22/n44 ), .A2(\us22/n2 ), .B0(
        \us22/n280 ), .Y(\us22/n339 ) );
  NAND2X1 \us23/U366  ( .A(\us23/n47 ), .B(\us23/n226 ), .Y(\us23/n189 ) );
  NOR2X1 \us23/U365  ( .A(\us23/n226 ), .B(sa23[3]), .Y(\us23/n242 ) );
  INVX1 \us23/U364  ( .A(\us23/n242 ), .Y(\us23/n205 ) );
  AND2X1 \us23/U363  ( .A(\us23/n189 ), .B(\us23/n205 ), .Y(\us23/n65 ) );
  NOR2X1 \us23/U362  ( .A(\us23/n226 ), .B(\us23/n47 ), .Y(\us23/n45 ) );
  NOR2X1 \us23/U361  ( .A(\us23/n259 ), .B(\us23/n45 ), .Y(\us23/n73 ) );
  NAND2BX1 \us23/U360  ( .AN(\us23/n73 ), .B(\us23/n6 ), .Y(\us23/n158 ) );
  NOR2X1 \us23/U359  ( .A(\us23/n226 ), .B(\us23/n159 ), .Y(\us23/n95 ) );
  INVX1 \us23/U358  ( .A(\us23/n95 ), .Y(\us23/n111 ) );
  NOR2X1 \us23/U357  ( .A(\us23/n145 ), .B(sa23[1]), .Y(\us23/n42 ) );
  INVX1 \us23/U356  ( .A(\us23/n42 ), .Y(\us23/n121 ) );
  INVX1 \us23/U355  ( .A(\us23/n47 ), .Y(\us23/n96 ) );
  OAI211X1 \us23/U354  ( .A0(\us23/n65 ), .A1(\us23/n27 ), .B0(\us23/n158 ), 
        .C0(\us23/n358 ), .Y(\us23/n355 ) );
  NOR2X1 \us23/U353  ( .A(\us23/n226 ), .B(\us23/n145 ), .Y(\us23/n59 ) );
  NOR2X1 \us23/U352  ( .A(\us23/n96 ), .B(\us23/n59 ), .Y(\us23/n271 ) );
  NOR2X1 \us23/U351  ( .A(\us23/n226 ), .B(\us23/n278 ), .Y(\us23/n217 ) );
  INVX1 \us23/U350  ( .A(\us23/n217 ), .Y(\us23/n150 ) );
  NAND2X1 \us23/U349  ( .A(\us23/n44 ), .B(\us23/n150 ), .Y(\us23/n147 ) );
  NAND2X1 \us23/U348  ( .A(sa23[4]), .B(\us23/n226 ), .Y(\us23/n101 ) );
  INVX1 \us23/U347  ( .A(\us23/n159 ), .Y(\us23/n188 ) );
  NOR2X1 \us23/U346  ( .A(\us23/n188 ), .B(\us23/n226 ), .Y(\us23/n25 ) );
  INVX1 \us23/U345  ( .A(\us23/n172 ), .Y(\us23/n107 ) );
  AOI22X1 \us23/U344  ( .A0(\us23/n33 ), .A1(\us23/n147 ), .B0(\us23/n24 ), 
        .B1(\us23/n107 ), .Y(\us23/n357 ) );
  OAI221XL \us23/U343  ( .A0(\us23/n18 ), .A1(\us23/n121 ), .B0(\us23/n271 ), 
        .B1(\us23/n20 ), .C0(\us23/n357 ), .Y(\us23/n356 ) );
  MXI2X1 \us23/U342  ( .A(\us23/n355 ), .B(\us23/n356 ), .S0(\us23/n252 ), .Y(
        \us23/n331 ) );
  INVX1 \us23/U341  ( .A(\us23/n59 ), .Y(\us23/n79 ) );
  AND2X1 \us23/U340  ( .A(\us23/n101 ), .B(\us23/n79 ), .Y(\us23/n325 ) );
  XNOR2X1 \us23/U339  ( .A(sa23[5]), .B(\us23/n226 ), .Y(\us23/n352 ) );
  NOR2X1 \us23/U338  ( .A(\us23/n226 ), .B(\us23/n136 ), .Y(\us23/n281 ) );
  INVX1 \us23/U337  ( .A(\us23/n281 ), .Y(\us23/n19 ) );
  NAND2X1 \us23/U336  ( .A(\us23/n145 ), .B(\us23/n226 ), .Y(\us23/n223 ) );
  AOI21X1 \us23/U335  ( .A0(\us23/n19 ), .A1(\us23/n223 ), .B0(\us23/n27 ), 
        .Y(\us23/n354 ) );
  AOI31X1 \us23/U334  ( .A0(\us23/n6 ), .A1(\us23/n352 ), .A2(\us23/n259 ), 
        .B0(\us23/n354 ), .Y(\us23/n353 ) );
  OAI221XL \us23/U333  ( .A0(\us23/n20 ), .A1(\us23/n34 ), .B0(\us23/n325 ), 
        .B1(\us23/n4 ), .C0(\us23/n353 ), .Y(\us23/n347 ) );
  INVX1 \us23/U332  ( .A(\us23/n352 ), .Y(\us23/n349 ) );
  NAND2X1 \us23/U331  ( .A(\us23/n278 ), .B(\us23/n6 ), .Y(\us23/n74 ) );
  OAI211X1 \us23/U330  ( .A0(\us23/n349 ), .A1(\us23/n74 ), .B0(\us23/n350 ), 
        .C0(\us23/n351 ), .Y(\us23/n348 ) );
  MXI2X1 \us23/U329  ( .A(\us23/n347 ), .B(\us23/n348 ), .S0(\us23/n252 ), .Y(
        \us23/n332 ) );
  NOR2X1 \us23/U328  ( .A(\us23/n44 ), .B(\us23/n226 ), .Y(\us23/n157 ) );
  INVX1 \us23/U327  ( .A(\us23/n157 ), .Y(\us23/n240 ) );
  NAND2X1 \us23/U326  ( .A(\us23/n240 ), .B(\us23/n189 ), .Y(\us23/n68 ) );
  NOR2X1 \us23/U325  ( .A(\us23/n20 ), .B(\us23/n159 ), .Y(\us23/n225 ) );
  NOR2X1 \us23/U324  ( .A(\us23/n225 ), .B(\us23/n40 ), .Y(\us23/n345 ) );
  INVX1 \us23/U323  ( .A(\us23/n278 ), .Y(\us23/n94 ) );
  NAND2X1 \us23/U322  ( .A(\us23/n94 ), .B(\us23/n226 ), .Y(\us23/n199 ) );
  NAND2X1 \us23/U321  ( .A(\us23/n199 ), .B(\us23/n205 ), .Y(\us23/n82 ) );
  NAND2X1 \us23/U320  ( .A(\us23/n19 ), .B(\us23/n199 ), .Y(\us23/n295 ) );
  NOR2X1 \us23/U319  ( .A(\us23/n226 ), .B(\us23/n259 ), .Y(\us23/n210 ) );
  NOR2X1 \us23/U318  ( .A(\us23/n27 ), .B(\us23/n210 ), .Y(\us23/n173 ) );
  MXI2X1 \us23/U317  ( .A(\us23/n345 ), .B(\us23/n346 ), .S0(\us23/n252 ), .Y(
        \us23/n342 ) );
  NOR2X1 \us23/U316  ( .A(sa23[1]), .B(sa23[3]), .Y(\us23/n163 ) );
  INVX1 \us23/U315  ( .A(\us23/n163 ), .Y(\us23/n37 ) );
  INVX1 \us23/U314  ( .A(\us23/n173 ), .Y(\us23/n344 ) );
  AOI21X1 \us23/U313  ( .A0(\us23/n240 ), .A1(\us23/n37 ), .B0(\us23/n344 ), 
        .Y(\us23/n343 ) );
  AOI211X1 \us23/U312  ( .A0(\us23/n5 ), .A1(\us23/n68 ), .B0(\us23/n342 ), 
        .C0(\us23/n343 ), .Y(\us23/n333 ) );
  NOR2X1 \us23/U311  ( .A(\us23/n18 ), .B(\us23/n226 ), .Y(\us23/n258 ) );
  NAND2X1 \us23/U310  ( .A(\us23/n278 ), .B(sa23[1]), .Y(\us23/n204 ) );
  NOR2X1 \us23/U309  ( .A(\us23/n188 ), .B(sa23[1]), .Y(\us23/n179 ) );
  INVX1 \us23/U308  ( .A(\us23/n179 ), .Y(\us23/n330 ) );
  NAND2X1 \us23/U307  ( .A(\us23/n204 ), .B(\us23/n330 ), .Y(\us23/n239 ) );
  NOR2X1 \us23/U306  ( .A(\us23/n136 ), .B(sa23[1]), .Y(\us23/n299 ) );
  NOR2X1 \us23/U305  ( .A(\us23/n299 ), .B(\us23/n210 ), .Y(\us23/n341 ) );
  OAI32X1 \us23/U304  ( .A0(\us23/n27 ), .A1(\us23/n278 ), .A2(\us23/n95 ), 
        .B0(\us23/n341 ), .B1(\us23/n4 ), .Y(\us23/n340 ) );
  INVX1 \us23/U303  ( .A(\us23/n45 ), .Y(\us23/n126 ) );
  NAND2X1 \us23/U302  ( .A(\us23/n126 ), .B(\us23/n101 ), .Y(\us23/n178 ) );
  NOR2X1 \us23/U301  ( .A(\us23/n18 ), .B(\us23/n136 ), .Y(\us23/n280 ) );
  OAI21XL \us23/U300  ( .A0(\us23/n4 ), .A1(\us23/n121 ), .B0(\us23/n339 ), 
        .Y(\us23/n338 ) );
  MXI2X1 \us23/U299  ( .A(\us23/n336 ), .B(\us23/n337 ), .S0(\us23/n252 ), .Y(
        \us23/n335 ) );
  NOR2X1 \us23/U298  ( .A(\us23/n258 ), .B(\us23/n335 ), .Y(\us23/n334 ) );
  MX4X1 \us23/U297  ( .A(\us23/n331 ), .B(\us23/n332 ), .C(\us23/n333 ), .D(
        \us23/n334 ), .S0(sa23[6]), .S1(\us23/n234 ), .Y(sa21_sr[0]) );
  INVX1 \us23/U296  ( .A(\us23/n299 ), .Y(\us23/n80 ) );
  NOR2X1 \us23/U295  ( .A(\us23/n111 ), .B(\us23/n18 ), .Y(\us23/n269 ) );
  INVX1 \us23/U294  ( .A(\us23/n269 ), .Y(\us23/n75 ) );
  OAI221XL \us23/U293  ( .A0(\us23/n18 ), .A1(\us23/n330 ), .B0(\us23/n20 ), 
        .B1(\us23/n80 ), .C0(\us23/n75 ), .Y(\us23/n329 ) );
  AOI221X1 \us23/U292  ( .A0(\us23/n325 ), .A1(\us23/n33 ), .B0(\us23/n24 ), 
        .B1(\us23/n303 ), .C0(\us23/n329 ), .Y(\us23/n319 ) );
  NOR2X1 \us23/U291  ( .A(\us23/n234 ), .B(sa23[5]), .Y(\us23/n14 ) );
  NOR2X1 \us23/U290  ( .A(\us23/n25 ), .B(\us23/n299 ), .Y(\us23/n313 ) );
  NAND2X1 \us23/U289  ( .A(\us23/n44 ), .B(\us23/n226 ), .Y(\us23/n300 ) );
  AND2X1 \us23/U288  ( .A(\us23/n300 ), .B(\us23/n240 ), .Y(\us23/n23 ) );
  OAI32X1 \us23/U287  ( .A0(\us23/n4 ), .A1(\us23/n145 ), .A2(\us23/n210 ), 
        .B0(\us23/n137 ), .B1(\us23/n27 ), .Y(\us23/n328 ) );
  NOR2X1 \us23/U286  ( .A(sa23[0]), .B(sa23[5]), .Y(\us23/n16 ) );
  INVX1 \us23/U285  ( .A(\us23/n16 ), .Y(\us23/n114 ) );
  INVX1 \us23/U284  ( .A(\us23/n145 ), .Y(\us23/n149 ) );
  NOR2X1 \us23/U283  ( .A(\us23/n47 ), .B(sa23[1]), .Y(\us23/n98 ) );
  INVX1 \us23/U282  ( .A(\us23/n98 ), .Y(\us23/n284 ) );
  OAI21XL \us23/U281  ( .A0(\us23/n69 ), .A1(\us23/n284 ), .B0(\us23/n27 ), 
        .Y(\us23/n327 ) );
  AOI31X1 \us23/U280  ( .A0(\us23/n111 ), .A1(\us23/n149 ), .A2(\us23/n327 ), 
        .B0(\us23/n225 ), .Y(\us23/n326 ) );
  OAI21XL \us23/U279  ( .A0(\us23/n325 ), .A1(\us23/n18 ), .B0(\us23/n326 ), 
        .Y(\us23/n322 ) );
  NAND2X1 \us23/U278  ( .A(\us23/n19 ), .B(\us23/n189 ), .Y(\us23/n71 ) );
  NOR2X1 \us23/U277  ( .A(\us23/n71 ), .B(\us23/n18 ), .Y(\us23/n135 ) );
  AOI21X1 \us23/U276  ( .A0(\us23/n40 ), .A1(sa23[4]), .B0(\us23/n135 ), .Y(
        \us23/n324 ) );
  OAI221XL \us23/U275  ( .A0(\us23/n47 ), .A1(\us23/n27 ), .B0(\us23/n65 ), 
        .B1(\us23/n20 ), .C0(\us23/n324 ), .Y(\us23/n323 ) );
  AOI22X1 \us23/U274  ( .A0(\us23/n55 ), .A1(\us23/n322 ), .B0(\us23/n89 ), 
        .B1(\us23/n323 ), .Y(\us23/n321 ) );
  OAI221XL \us23/U273  ( .A0(\us23/n319 ), .A1(\us23/n52 ), .B0(\us23/n320 ), 
        .B1(\us23/n114 ), .C0(\us23/n321 ), .Y(\us23/n304 ) );
  NOR2X1 \us23/U272  ( .A(\us23/n226 ), .B(\us23/n58 ), .Y(\us23/n290 ) );
  INVX1 \us23/U271  ( .A(\us23/n290 ), .Y(\us23/n200 ) );
  NAND2X1 \us23/U270  ( .A(\us23/n34 ), .B(\us23/n200 ), .Y(\us23/n120 ) );
  INVX1 \us23/U269  ( .A(\us23/n210 ), .Y(\us23/n100 ) );
  OAI221XL \us23/U268  ( .A0(\us23/n20 ), .A1(\us23/n100 ), .B0(sa23[3]), .B1(
        \us23/n4 ), .C0(\us23/n262 ), .Y(\us23/n317 ) );
  INVX1 \us23/U267  ( .A(\us23/n258 ), .Y(\us23/n182 ) );
  AOI211X1 \us23/U266  ( .A0(\us23/n33 ), .A1(\us23/n120 ), .B0(\us23/n317 ), 
        .C0(\us23/n318 ), .Y(\us23/n306 ) );
  NAND2X1 \us23/U265  ( .A(\us23/n100 ), .B(\us23/n199 ), .Y(\us23/n151 ) );
  INVX1 \us23/U264  ( .A(\us23/n151 ), .Y(\us23/n314 ) );
  NOR2X1 \us23/U263  ( .A(\us23/n45 ), .B(\us23/n163 ), .Y(\us23/n160 ) );
  INVX1 \us23/U262  ( .A(\us23/n295 ), .Y(\us23/n92 ) );
  AOI21X1 \us23/U261  ( .A0(sa23[1]), .A1(\us23/n58 ), .B0(\us23/n98 ), .Y(
        \us23/n316 ) );
  OAI22X1 \us23/U260  ( .A0(\us23/n92 ), .A1(\us23/n18 ), .B0(\us23/n316 ), 
        .B1(\us23/n27 ), .Y(\us23/n315 ) );
  NOR2X1 \us23/U259  ( .A(\us23/n149 ), .B(\us23/n226 ), .Y(\us23/n41 ) );
  INVX1 \us23/U258  ( .A(\us23/n41 ), .Y(\us23/n105 ) );
  NAND2X1 \us23/U257  ( .A(\us23/n284 ), .B(\us23/n105 ), .Y(\us23/n227 ) );
  AOI21X1 \us23/U256  ( .A0(\us23/n313 ), .A1(\us23/n33 ), .B0(\us23/n269 ), 
        .Y(\us23/n312 ) );
  OAI221XL \us23/U255  ( .A0(\us23/n149 ), .A1(\us23/n20 ), .B0(\us23/n4 ), 
        .B1(\us23/n227 ), .C0(\us23/n312 ), .Y(\us23/n309 ) );
  AOI21X1 \us23/U254  ( .A0(\us23/n226 ), .A1(\us23/n188 ), .B0(\us23/n242 ), 
        .Y(\us23/n185 ) );
  INVX1 \us23/U253  ( .A(\us23/n185 ), .Y(\us23/n48 ) );
  AND2X1 \us23/U252  ( .A(\us23/n223 ), .B(\us23/n240 ), .Y(\us23/n28 ) );
  OAI221XL \us23/U251  ( .A0(\us23/n27 ), .A1(\us23/n44 ), .B0(\us23/n4 ), 
        .B1(\us23/n48 ), .C0(\us23/n311 ), .Y(\us23/n310 ) );
  AOI22X1 \us23/U250  ( .A0(\us23/n89 ), .A1(\us23/n309 ), .B0(\us23/n55 ), 
        .B1(\us23/n310 ), .Y(\us23/n308 ) );
  OAI221XL \us23/U249  ( .A0(\us23/n306 ), .A1(\us23/n52 ), .B0(\us23/n307 ), 
        .B1(\us23/n114 ), .C0(\us23/n308 ), .Y(\us23/n305 ) );
  MX2X1 \us23/U248  ( .A(\us23/n304 ), .B(\us23/n305 ), .S0(sa23[6]), .Y(
        sa21_sr[1]) );
  INVX1 \us23/U247  ( .A(\us23/n187 ), .Y(\us23/n61 ) );
  MXI2X1 \us23/U246  ( .A(\us23/n303 ), .B(\us23/n61 ), .S0(\us23/n69 ), .Y(
        \us23/n301 ) );
  MXI2X1 \us23/U245  ( .A(\us23/n301 ), .B(\us23/n147 ), .S0(\us23/n302 ), .Y(
        \us23/n285 ) );
  NAND2X1 \us23/U244  ( .A(\us23/n200 ), .B(\us23/n300 ), .Y(\us23/n99 ) );
  INVX1 \us23/U243  ( .A(\us23/n99 ), .Y(\us23/n296 ) );
  NOR2X1 \us23/U242  ( .A(\us23/n299 ), .B(\us23/n242 ), .Y(\us23/n298 ) );
  NAND2X1 \us23/U241  ( .A(sa23[1]), .B(\us23/n47 ), .Y(\us23/n122 ) );
  NOR2X1 \us23/U240  ( .A(\us23/n159 ), .B(\us23/n217 ), .Y(\us23/n198 ) );
  OAI221XL \us23/U239  ( .A0(\us23/n298 ), .A1(\us23/n27 ), .B0(\us23/n20 ), 
        .B1(\us23/n122 ), .C0(\us23/n132 ), .Y(\us23/n297 ) );
  AOI221X1 \us23/U238  ( .A0(\us23/n225 ), .A1(\us23/n226 ), .B0(\us23/n296 ), 
        .B1(\us23/n6 ), .C0(\us23/n297 ), .Y(\us23/n291 ) );
  OAI2BB2X1 \us23/U237  ( .B0(\us23/n27 ), .B1(\us23/n295 ), .A0N(\us23/n34 ), 
        .A1N(\us23/n24 ), .Y(\us23/n293 ) );
  AOI21X1 \us23/U236  ( .A0(\us23/n101 ), .A1(\us23/n150 ), .B0(\us23/n20 ), 
        .Y(\us23/n294 ) );
  AOI211X1 \us23/U235  ( .A0(\us23/n5 ), .A1(\us23/n79 ), .B0(\us23/n293 ), 
        .C0(\us23/n294 ), .Y(\us23/n292 ) );
  INVX1 \us23/U234  ( .A(\us23/n89 ), .Y(\us23/n10 ) );
  OAI22X1 \us23/U233  ( .A0(\us23/n291 ), .A1(\us23/n114 ), .B0(\us23/n292 ), 
        .B1(\us23/n10 ), .Y(\us23/n286 ) );
  INVX1 \us23/U232  ( .A(\us23/n225 ), .Y(\us23/n288 ) );
  NAND2X1 \us23/U231  ( .A(\us23/n200 ), .B(\us23/n284 ), .Y(\us23/n102 ) );
  NOR2X1 \us23/U230  ( .A(\us23/n290 ), .B(\us23/n163 ), .Y(\us23/n184 ) );
  AOI22X1 \us23/U229  ( .A0(\us23/n102 ), .A1(\us23/n69 ), .B0(\us23/n184 ), 
        .B1(\us23/n33 ), .Y(\us23/n289 ) );
  AOI31X1 \us23/U228  ( .A0(\us23/n132 ), .A1(\us23/n288 ), .A2(\us23/n289 ), 
        .B0(\us23/n52 ), .Y(\us23/n287 ) );
  AOI211X1 \us23/U227  ( .A0(\us23/n285 ), .A1(\us23/n55 ), .B0(\us23/n286 ), 
        .C0(\us23/n287 ), .Y(\us23/n263 ) );
  NAND2X1 \us23/U226  ( .A(\us23/n284 ), .B(\us23/n122 ), .Y(\us23/n125 ) );
  NOR2X1 \us23/U225  ( .A(\us23/n199 ), .B(\us23/n4 ), .Y(\us23/n50 ) );
  AOI21X1 \us23/U224  ( .A0(\us23/n200 ), .A1(\us23/n223 ), .B0(\us23/n20 ), 
        .Y(\us23/n283 ) );
  AOI211X1 \us23/U223  ( .A0(\us23/n5 ), .A1(\us23/n125 ), .B0(\us23/n50 ), 
        .C0(\us23/n283 ), .Y(\us23/n282 ) );
  OAI221XL \us23/U222  ( .A0(\us23/n281 ), .A1(\us23/n27 ), .B0(\us23/n4 ), 
        .B1(\us23/n111 ), .C0(\us23/n282 ), .Y(\us23/n265 ) );
  INVX1 \us23/U221  ( .A(\us23/n280 ), .Y(\us23/n247 ) );
  NAND2X1 \us23/U220  ( .A(\us23/n41 ), .B(\us23/n33 ), .Y(\us23/n272 ) );
  OAI221XL \us23/U219  ( .A0(sa23[1]), .A1(\us23/n247 ), .B0(\us23/n4 ), .B1(
        \us23/n189 ), .C0(\us23/n272 ), .Y(\us23/n279 ) );
  NAND2X1 \us23/U218  ( .A(sa23[2]), .B(\us23/n149 ), .Y(\us23/n276 ) );
  XNOR2X1 \us23/U217  ( .A(\us23/n129 ), .B(sa23[1]), .Y(\us23/n155 ) );
  MXI2X1 \us23/U216  ( .A(\us23/n276 ), .B(\us23/n277 ), .S0(\us23/n155 ), .Y(
        \us23/n275 ) );
  OAI22X1 \us23/U215  ( .A0(\us23/n273 ), .A1(\us23/n10 ), .B0(\us23/n274 ), 
        .B1(\us23/n52 ), .Y(\us23/n266 ) );
  NOR2X1 \us23/U214  ( .A(\us23/n20 ), .B(\us23/n226 ), .Y(\us23/n176 ) );
  OAI21XL \us23/U213  ( .A0(\us23/n4 ), .A1(\us23/n271 ), .B0(\us23/n272 ), 
        .Y(\us23/n270 ) );
  OAI31X1 \us23/U212  ( .A0(\us23/n176 ), .A1(\us23/n269 ), .A2(\us23/n270 ), 
        .B0(\us23/n16 ), .Y(\us23/n268 ) );
  INVX1 \us23/U211  ( .A(\us23/n268 ), .Y(\us23/n267 ) );
  AOI211X1 \us23/U210  ( .A0(\us23/n55 ), .A1(\us23/n265 ), .B0(\us23/n266 ), 
        .C0(\us23/n267 ), .Y(\us23/n264 ) );
  MXI2X1 \us23/U209  ( .A(\us23/n263 ), .B(\us23/n264 ), .S0(sa23[6]), .Y(
        sa21_sr[2]) );
  NOR2X1 \us23/U208  ( .A(\us23/n94 ), .B(sa23[1]), .Y(\us23/n211 ) );
  INVX1 \us23/U207  ( .A(\us23/n262 ), .Y(\us23/n261 ) );
  AOI211X1 \us23/U206  ( .A0(\us23/n259 ), .A1(\us23/n24 ), .B0(\us23/n260 ), 
        .C0(\us23/n261 ), .Y(\us23/n255 ) );
  OAI22X1 \us23/U205  ( .A0(\us23/n20 ), .A1(\us23/n68 ), .B0(\us23/n27 ), 
        .B1(\us23/n37 ), .Y(\us23/n257 ) );
  NOR3X1 \us23/U204  ( .A(\us23/n257 ), .B(\us23/n258 ), .C(\us23/n50 ), .Y(
        \us23/n256 ) );
  MXI2X1 \us23/U203  ( .A(\us23/n255 ), .B(\us23/n256 ), .S0(\us23/n252 ), .Y(
        \us23/n254 ) );
  AOI221X1 \us23/U202  ( .A0(\us23/n211 ), .A1(\us23/n5 ), .B0(\us23/n40 ), 
        .B1(sa23[4]), .C0(\us23/n254 ), .Y(\us23/n248 ) );
  INVX1 \us23/U201  ( .A(\us23/n211 ), .Y(\us23/n106 ) );
  NAND2X1 \us23/U200  ( .A(\us23/n200 ), .B(\us23/n106 ), .Y(\us23/n83 ) );
  NAND2X1 \us23/U199  ( .A(\us23/n199 ), .B(\us23/n204 ), .Y(\us23/n169 ) );
  AOI2BB2X1 \us23/U198  ( .B0(\us23/n65 ), .B1(\us23/n24 ), .A0N(\us23/n169 ), 
        .A1N(\us23/n20 ), .Y(\us23/n253 ) );
  OAI221XL \us23/U197  ( .A0(\us23/n172 ), .A1(\us23/n18 ), .B0(\us23/n27 ), 
        .B1(\us23/n83 ), .C0(\us23/n253 ), .Y(\us23/n251 ) );
  MXI2X1 \us23/U196  ( .A(\us23/n250 ), .B(\us23/n251 ), .S0(\us23/n252 ), .Y(
        \us23/n249 ) );
  MXI2X1 \us23/U195  ( .A(\us23/n248 ), .B(\us23/n249 ), .S0(\us23/n234 ), .Y(
        \us23/n228 ) );
  OAI21XL \us23/U194  ( .A0(\us23/n58 ), .A1(\us23/n27 ), .B0(\us23/n247 ), 
        .Y(\us23/n245 ) );
  NOR2X1 \us23/U193  ( .A(sa23[7]), .B(\us23/n145 ), .Y(\us23/n246 ) );
  XNOR2X1 \us23/U192  ( .A(\us23/n69 ), .B(sa23[1]), .Y(\us23/n130 ) );
  MXI2X1 \us23/U191  ( .A(\us23/n245 ), .B(\us23/n246 ), .S0(\us23/n130 ), .Y(
        \us23/n243 ) );
  OAI211X1 \us23/U190  ( .A0(\us23/n4 ), .A1(\us23/n149 ), .B0(\us23/n243 ), 
        .C0(\us23/n244 ), .Y(\us23/n230 ) );
  NOR2X1 \us23/U189  ( .A(\us23/n242 ), .B(\us23/n137 ), .Y(\us23/n70 ) );
  OAI221XL \us23/U188  ( .A0(\us23/n159 ), .A1(\us23/n27 ), .B0(\us23/n20 ), 
        .B1(\us23/n34 ), .C0(\us23/n241 ), .Y(\us23/n231 ) );
  NAND2X1 \us23/U187  ( .A(\us23/n101 ), .B(\us23/n240 ), .Y(\us23/n76 ) );
  AOI21X1 \us23/U186  ( .A0(\us23/n122 ), .A1(\us23/n106 ), .B0(\us23/n129 ), 
        .Y(\us23/n237 ) );
  INVX1 \us23/U185  ( .A(\us23/n239 ), .Y(\us23/n238 ) );
  OAI21XL \us23/U184  ( .A0(\us23/n237 ), .A1(\us23/n43 ), .B0(\us23/n238 ), 
        .Y(\us23/n236 ) );
  OAI221XL \us23/U183  ( .A0(\us23/n18 ), .A1(\us23/n76 ), .B0(\us23/n59 ), 
        .B1(\us23/n27 ), .C0(\us23/n236 ), .Y(\us23/n232 ) );
  AOI2BB2X1 \us23/U182  ( .B0(\us23/n24 ), .B1(\us23/n187 ), .A0N(\us23/n227 ), 
        .A1N(\us23/n20 ), .Y(\us23/n235 ) );
  OAI211X1 \us23/U181  ( .A0(\us23/n27 ), .A1(\us23/n122 ), .B0(\us23/n158 ), 
        .C0(\us23/n235 ), .Y(\us23/n233 ) );
  MX4X1 \us23/U180  ( .A(\us23/n230 ), .B(\us23/n231 ), .C(\us23/n232 ), .D(
        \us23/n233 ), .S0(\us23/n234 ), .S1(sa23[5]), .Y(\us23/n229 ) );
  MX2X1 \us23/U179  ( .A(\us23/n228 ), .B(\us23/n229 ), .S0(sa23[6]), .Y(
        sa21_sr[3]) );
  NOR2BX1 \us23/U178  ( .AN(\us23/n204 ), .B(\us23/n137 ), .Y(\us23/n110 ) );
  INVX1 \us23/U177  ( .A(\us23/n110 ), .Y(\us23/n64 ) );
  AOI22X1 \us23/U176  ( .A0(\us23/n225 ), .A1(\us23/n226 ), .B0(\us23/n6 ), 
        .B1(\us23/n227 ), .Y(\us23/n224 ) );
  OAI221XL \us23/U175  ( .A0(\us23/n27 ), .A1(\us23/n64 ), .B0(\us23/n4 ), 
        .B1(\us23/n83 ), .C0(\us23/n224 ), .Y(\us23/n212 ) );
  NAND2X1 \us23/U174  ( .A(\us23/n34 ), .B(\us23/n204 ), .Y(\us23/n221 ) );
  OAI21XL \us23/U173  ( .A0(\us23/n69 ), .A1(\us23/n223 ), .B0(\us23/n27 ), 
        .Y(\us23/n222 ) );
  NOR2X1 \us23/U172  ( .A(\us23/n217 ), .B(\us23/n42 ), .Y(\us23/n208 ) );
  AOI211X1 \us23/U171  ( .A0(\us23/n208 ), .A1(\us23/n5 ), .B0(\us23/n220 ), 
        .C0(\us23/n173 ), .Y(\us23/n219 ) );
  OAI22X1 \us23/U170  ( .A0(\us23/n218 ), .A1(\us23/n10 ), .B0(\us23/n219 ), 
        .B1(\us23/n114 ), .Y(\us23/n213 ) );
  INVX1 \us23/U169  ( .A(\us23/n135 ), .Y(\us23/n215 ) );
  NOR2X1 \us23/U168  ( .A(\us23/n4 ), .B(\us23/n159 ), .Y(\us23/n31 ) );
  INVX1 \us23/U167  ( .A(\us23/n31 ), .Y(\us23/n196 ) );
  AOI31X1 \us23/U166  ( .A0(\us23/n215 ), .A1(\us23/n196 ), .A2(\us23/n216 ), 
        .B0(\us23/n52 ), .Y(\us23/n214 ) );
  AOI211X1 \us23/U165  ( .A0(\us23/n55 ), .A1(\us23/n212 ), .B0(\us23/n213 ), 
        .C0(\us23/n214 ), .Y(\us23/n190 ) );
  INVX1 \us23/U164  ( .A(\us23/n207 ), .Y(\us23/n192 ) );
  NOR2X1 \us23/U163  ( .A(\us23/n25 ), .B(\us23/n98 ), .Y(\us23/n32 ) );
  OAI22X1 \us23/U162  ( .A0(\us23/n28 ), .A1(\us23/n4 ), .B0(\us23/n188 ), 
        .B1(\us23/n27 ), .Y(\us23/n206 ) );
  NAND2X1 \us23/U161  ( .A(\us23/n204 ), .B(\us23/n80 ), .Y(\us23/n118 ) );
  INVX1 \us23/U160  ( .A(\us23/n118 ), .Y(\us23/n123 ) );
  NAND2X1 \us23/U159  ( .A(\us23/n94 ), .B(\us23/n79 ), .Y(\us23/n203 ) );
  OAI2BB1X1 \us23/U158  ( .A0N(\us23/n199 ), .A1N(\us23/n200 ), .B0(\us23/n33 ), .Y(\us23/n195 ) );
  INVX1 \us23/U157  ( .A(\us23/n55 ), .Y(\us23/n12 ) );
  AOI31X1 \us23/U156  ( .A0(\us23/n195 ), .A1(\us23/n196 ), .A2(\us23/n197 ), 
        .B0(\us23/n12 ), .Y(\us23/n194 ) );
  AOI211X1 \us23/U155  ( .A0(\us23/n89 ), .A1(\us23/n192 ), .B0(\us23/n193 ), 
        .C0(\us23/n194 ), .Y(\us23/n191 ) );
  MXI2X1 \us23/U154  ( .A(\us23/n190 ), .B(\us23/n191 ), .S0(sa23[6]), .Y(
        sa21_sr[4]) );
  OAI21XL \us23/U153  ( .A0(\us23/n69 ), .A1(\us23/n189 ), .B0(\us23/n27 ), 
        .Y(\us23/n186 ) );
  INVX1 \us23/U152  ( .A(\us23/n183 ), .Y(\us23/n180 ) );
  NAND2X1 \us23/U151  ( .A(\us23/n74 ), .B(\us23/n182 ), .Y(\us23/n181 ) );
  AOI211X1 \us23/U150  ( .A0(\us23/n179 ), .A1(\us23/n24 ), .B0(\us23/n180 ), 
        .C0(\us23/n181 ), .Y(\us23/n165 ) );
  INVX1 \us23/U149  ( .A(\us23/n178 ), .Y(\us23/n175 ) );
  AOI211X1 \us23/U148  ( .A0(\us23/n175 ), .A1(\us23/n5 ), .B0(\us23/n176 ), 
        .C0(\us23/n177 ), .Y(\us23/n174 ) );
  OAI221XL \us23/U147  ( .A0(\us23/n159 ), .A1(\us23/n27 ), .B0(\us23/n145 ), 
        .B1(\us23/n20 ), .C0(\us23/n174 ), .Y(\us23/n167 ) );
  MXI2X1 \us23/U146  ( .A(\us23/n40 ), .B(\us23/n173 ), .S0(\us23/n96 ), .Y(
        \us23/n170 ) );
  AOI22X1 \us23/U145  ( .A0(\us23/n137 ), .A1(\us23/n24 ), .B0(\us23/n172 ), 
        .B1(\us23/n6 ), .Y(\us23/n171 ) );
  OAI211X1 \us23/U144  ( .A0(\us23/n20 ), .A1(\us23/n169 ), .B0(\us23/n170 ), 
        .C0(\us23/n171 ), .Y(\us23/n168 ) );
  AOI22X1 \us23/U143  ( .A0(\us23/n89 ), .A1(\us23/n167 ), .B0(\us23/n55 ), 
        .B1(\us23/n168 ), .Y(\us23/n166 ) );
  OAI221XL \us23/U142  ( .A0(\us23/n164 ), .A1(\us23/n114 ), .B0(\us23/n165 ), 
        .B1(\us23/n52 ), .C0(\us23/n166 ), .Y(\us23/n138 ) );
  OAI21XL \us23/U141  ( .A0(\us23/n41 ), .A1(\us23/n163 ), .B0(\us23/n69 ), 
        .Y(\us23/n162 ) );
  AOI221X1 \us23/U140  ( .A0(\us23/n159 ), .A1(\us23/n24 ), .B0(\us23/n160 ), 
        .B1(\us23/n33 ), .C0(\us23/n161 ), .Y(\us23/n140 ) );
  OAI21XL \us23/U139  ( .A0(\us23/n157 ), .A1(\us23/n20 ), .B0(\us23/n158 ), 
        .Y(\us23/n156 ) );
  NOR2X1 \us23/U138  ( .A(\us23/n4 ), .B(\us23/n136 ), .Y(\us23/n153 ) );
  NOR2X1 \us23/U137  ( .A(\us23/n145 ), .B(\us23/n69 ), .Y(\us23/n154 ) );
  MXI2X1 \us23/U136  ( .A(\us23/n153 ), .B(\us23/n154 ), .S0(\us23/n155 ), .Y(
        \us23/n152 ) );
  OAI221XL \us23/U135  ( .A0(\us23/n110 ), .A1(\us23/n18 ), .B0(\us23/n20 ), 
        .B1(\us23/n151 ), .C0(\us23/n152 ), .Y(\us23/n143 ) );
  AOI21X1 \us23/U134  ( .A0(\us23/n149 ), .A1(\us23/n150 ), .B0(\us23/n18 ), 
        .Y(\us23/n148 ) );
  AOI2BB1X1 \us23/U133  ( .A0N(\us23/n147 ), .A1N(\us23/n27 ), .B0(\us23/n148 ), .Y(\us23/n146 ) );
  OAI221XL \us23/U132  ( .A0(\us23/n145 ), .A1(\us23/n20 ), .B0(\us23/n4 ), 
        .B1(\us23/n34 ), .C0(\us23/n146 ), .Y(\us23/n144 ) );
  AOI22X1 \us23/U131  ( .A0(\us23/n89 ), .A1(\us23/n143 ), .B0(\us23/n14 ), 
        .B1(\us23/n144 ), .Y(\us23/n142 ) );
  OAI221XL \us23/U130  ( .A0(\us23/n140 ), .A1(\us23/n12 ), .B0(\us23/n141 ), 
        .B1(\us23/n114 ), .C0(\us23/n142 ), .Y(\us23/n139 ) );
  MX2X1 \us23/U129  ( .A(\us23/n138 ), .B(\us23/n139 ), .S0(sa23[6]), .Y(
        sa21_sr[5]) );
  INVX1 \us23/U128  ( .A(\us23/n70 ), .Y(\us23/n133 ) );
  OAI22X1 \us23/U127  ( .A0(\us23/n4 ), .A1(\us23/n136 ), .B0(\us23/n137 ), 
        .B1(\us23/n27 ), .Y(\us23/n134 ) );
  AOI211X1 \us23/U126  ( .A0(\us23/n133 ), .A1(\us23/n69 ), .B0(\us23/n134 ), 
        .C0(\us23/n135 ), .Y(\us23/n112 ) );
  INVX1 \us23/U125  ( .A(\us23/n132 ), .Y(\us23/n131 ) );
  OAI21XL \us23/U124  ( .A0(\us23/n18 ), .A1(\us23/n37 ), .B0(\us23/n128 ), 
        .Y(\us23/n127 ) );
  OAI221XL \us23/U123  ( .A0(\us23/n18 ), .A1(\us23/n105 ), .B0(\us23/n123 ), 
        .B1(\us23/n27 ), .C0(\us23/n124 ), .Y(\us23/n116 ) );
  NAND2X1 \us23/U122  ( .A(\us23/n121 ), .B(\us23/n122 ), .Y(\us23/n30 ) );
  OAI221XL \us23/U121  ( .A0(\us23/n18 ), .A1(\us23/n118 ), .B0(\us23/n27 ), 
        .B1(\us23/n30 ), .C0(\us23/n119 ), .Y(\us23/n117 ) );
  AOI22X1 \us23/U120  ( .A0(\us23/n89 ), .A1(\us23/n116 ), .B0(\us23/n55 ), 
        .B1(\us23/n117 ), .Y(\us23/n115 ) );
  OAI221XL \us23/U119  ( .A0(\us23/n112 ), .A1(\us23/n52 ), .B0(\us23/n113 ), 
        .B1(\us23/n114 ), .C0(\us23/n115 ), .Y(\us23/n84 ) );
  OAI22X1 \us23/U118  ( .A0(\us23/n110 ), .A1(\us23/n4 ), .B0(\us23/n20 ), 
        .B1(\us23/n21 ), .Y(\us23/n108 ) );
  AOI21X1 \us23/U117  ( .A0(sa23[1]), .A1(\us23/n58 ), .B0(\us23/n27 ), .Y(
        \us23/n109 ) );
  AOI211X1 \us23/U116  ( .A0(\us23/n5 ), .A1(\us23/n107 ), .B0(\us23/n108 ), 
        .C0(\us23/n109 ), .Y(\us23/n86 ) );
  OAI22X1 \us23/U115  ( .A0(\us23/n45 ), .A1(\us23/n4 ), .B0(sa23[4]), .B1(
        \us23/n18 ), .Y(\us23/n103 ) );
  AOI21X1 \us23/U114  ( .A0(\us23/n105 ), .A1(\us23/n106 ), .B0(\us23/n20 ), 
        .Y(\us23/n104 ) );
  AOI211X1 \us23/U113  ( .A0(\us23/n33 ), .A1(\us23/n102 ), .B0(\us23/n103 ), 
        .C0(\us23/n104 ), .Y(\us23/n87 ) );
  NAND2X1 \us23/U112  ( .A(\us23/n100 ), .B(\us23/n101 ), .Y(\us23/n62 ) );
  OAI221XL \us23/U111  ( .A0(\us23/n27 ), .A1(\us23/n62 ), .B0(\us23/n4 ), 
        .B1(\us23/n21 ), .C0(\us23/n97 ), .Y(\us23/n90 ) );
  NOR3X1 \us23/U110  ( .A(\us23/n4 ), .B(\us23/n95 ), .C(\us23/n96 ), .Y(
        \us23/n67 ) );
  AOI31X1 \us23/U109  ( .A0(\us23/n79 ), .A1(\us23/n94 ), .A2(\us23/n6 ), .B0(
        \us23/n67 ), .Y(\us23/n93 ) );
  OAI221XL \us23/U108  ( .A0(\us23/n73 ), .A1(\us23/n27 ), .B0(\us23/n92 ), 
        .B1(\us23/n20 ), .C0(\us23/n93 ), .Y(\us23/n91 ) );
  AOI22X1 \us23/U107  ( .A0(\us23/n89 ), .A1(\us23/n90 ), .B0(\us23/n16 ), 
        .B1(\us23/n91 ), .Y(\us23/n88 ) );
  OAI221XL \us23/U106  ( .A0(\us23/n86 ), .A1(\us23/n52 ), .B0(\us23/n87 ), 
        .B1(\us23/n12 ), .C0(\us23/n88 ), .Y(\us23/n85 ) );
  MX2X1 \us23/U105  ( .A(\us23/n84 ), .B(\us23/n85 ), .S0(sa23[6]), .Y(
        sa21_sr[6]) );
  INVX1 \us23/U104  ( .A(\us23/n81 ), .Y(\us23/n77 ) );
  AOI21X1 \us23/U103  ( .A0(\us23/n79 ), .A1(\us23/n80 ), .B0(\us23/n27 ), .Y(
        \us23/n78 ) );
  AOI211X1 \us23/U102  ( .A0(\us23/n5 ), .A1(\us23/n76 ), .B0(\us23/n77 ), 
        .C0(\us23/n78 ), .Y(\us23/n51 ) );
  OAI211X1 \us23/U101  ( .A0(\us23/n73 ), .A1(\us23/n27 ), .B0(\us23/n74 ), 
        .C0(\us23/n75 ), .Y(\us23/n72 ) );
  AOI21X1 \us23/U100  ( .A0(\us23/n68 ), .A1(\us23/n69 ), .B0(\us23/n6 ), .Y(
        \us23/n63 ) );
  INVX1 \us23/U99  ( .A(\us23/n67 ), .Y(\us23/n66 ) );
  OAI221XL \us23/U98  ( .A0(\us23/n63 ), .A1(\us23/n64 ), .B0(\us23/n65 ), 
        .B1(\us23/n27 ), .C0(\us23/n66 ), .Y(\us23/n56 ) );
  AOI2BB2X1 \us23/U97  ( .B0(\us23/n61 ), .B1(\us23/n24 ), .A0N(\us23/n62 ), 
        .A1N(\us23/n20 ), .Y(\us23/n60 ) );
  OAI221XL \us23/U96  ( .A0(\us23/n58 ), .A1(\us23/n18 ), .B0(\us23/n59 ), 
        .B1(\us23/n27 ), .C0(\us23/n60 ), .Y(\us23/n57 ) );
  AOI22X1 \us23/U95  ( .A0(\us23/n55 ), .A1(\us23/n56 ), .B0(\us23/n16 ), .B1(
        \us23/n57 ), .Y(\us23/n54 ) );
  OAI221XL \us23/U94  ( .A0(\us23/n51 ), .A1(\us23/n52 ), .B0(\us23/n53 ), 
        .B1(\us23/n10 ), .C0(\us23/n54 ), .Y(\us23/n7 ) );
  INVX1 \us23/U93  ( .A(\us23/n50 ), .Y(\us23/n49 ) );
  OAI221XL \us23/U92  ( .A0(\us23/n47 ), .A1(\us23/n18 ), .B0(\us23/n27 ), 
        .B1(\us23/n48 ), .C0(\us23/n49 ), .Y(\us23/n46 ) );
  NOR2X1 \us23/U91  ( .A(\us23/n41 ), .B(\us23/n42 ), .Y(\us23/n38 ) );
  INVX1 \us23/U90  ( .A(\us23/n40 ), .Y(\us23/n39 ) );
  INVX1 \us23/U89  ( .A(\us23/n32 ), .Y(\us23/n26 ) );
  AOI21X1 \us23/U88  ( .A0(\us23/n5 ), .A1(\us23/n30 ), .B0(\us23/n31 ), .Y(
        \us23/n29 ) );
  OAI221XL \us23/U87  ( .A0(\us23/n26 ), .A1(\us23/n27 ), .B0(\us23/n28 ), 
        .B1(\us23/n20 ), .C0(\us23/n29 ), .Y(\us23/n15 ) );
  OAI221XL \us23/U86  ( .A0(\us23/n18 ), .A1(\us23/n19 ), .B0(\us23/n20 ), 
        .B1(\us23/n21 ), .C0(\us23/n22 ), .Y(\us23/n17 ) );
  AOI22X1 \us23/U85  ( .A0(\us23/n14 ), .A1(\us23/n15 ), .B0(\us23/n16 ), .B1(
        \us23/n17 ), .Y(\us23/n13 ) );
  OAI221XL \us23/U84  ( .A0(\us23/n9 ), .A1(\us23/n10 ), .B0(\us23/n11 ), .B1(
        \us23/n12 ), .C0(\us23/n13 ), .Y(\us23/n8 ) );
  MX2X1 \us23/U83  ( .A(\us23/n7 ), .B(\us23/n8 ), .S0(sa23[6]), .Y(sa21_sr[7]) );
  NOR2X4 \us23/U82  ( .A(\us23/n129 ), .B(sa23[2]), .Y(\us23/n43 ) );
  CLKINVX3 \us23/U81  ( .A(\us23/n14 ), .Y(\us23/n52 ) );
  OAI22XL \us23/U80  ( .A0(\us23/n201 ), .A1(\us23/n52 ), .B0(\us23/n202 ), 
        .B1(\us23/n114 ), .Y(\us23/n193 ) );
  CLKINVX3 \us23/U79  ( .A(sa23[5]), .Y(\us23/n252 ) );
  NOR2X2 \us23/U78  ( .A(\us23/n252 ), .B(\us23/n234 ), .Y(\us23/n55 ) );
  CLKINVX3 \us23/U77  ( .A(sa23[7]), .Y(\us23/n129 ) );
  NOR2X4 \us23/U76  ( .A(\us23/n129 ), .B(\us23/n69 ), .Y(\us23/n24 ) );
  AOI22XL \us23/U75  ( .A0(\us23/n70 ), .A1(\us23/n24 ), .B0(\us23/n96 ), .B1(
        \us23/n129 ), .Y(\us23/n241 ) );
  NOR2X2 \us23/U74  ( .A(\us23/n252 ), .B(sa23[0]), .Y(\us23/n89 ) );
  CLKINVX3 \us23/U73  ( .A(sa23[0]), .Y(\us23/n234 ) );
  NOR2X4 \us23/U72  ( .A(\us23/n69 ), .B(sa23[7]), .Y(\us23/n33 ) );
  INVX12 \us23/U71  ( .A(\us23/n33 ), .Y(\us23/n27 ) );
  CLKINVX3 \us23/U70  ( .A(\us23/n1 ), .Y(\us23/n6 ) );
  CLKINVX3 \us23/U69  ( .A(\us23/n1 ), .Y(\us23/n5 ) );
  INVXL \us23/U68  ( .A(\us23/n24 ), .Y(\us23/n36 ) );
  INVX4 \us23/U67  ( .A(\us23/n3 ), .Y(\us23/n4 ) );
  INVXL \us23/U66  ( .A(\us23/n36 ), .Y(\us23/n3 ) );
  INVX4 \us23/U65  ( .A(sa23[1]), .Y(\us23/n226 ) );
  INVX4 \us23/U64  ( .A(\us23/n43 ), .Y(\us23/n20 ) );
  AOI221X4 \us23/U63  ( .A0(\us23/n24 ), .A1(\us23/n82 ), .B0(\us23/n43 ), 
        .B1(\us23/n295 ), .C0(\us23/n173 ), .Y(\us23/n346 ) );
  AOI221X4 \us23/U62  ( .A0(\us23/n5 ), .A1(\us23/n96 ), .B0(\us23/n43 ), .B1(
        \us23/n239 ), .C0(\us23/n340 ), .Y(\us23/n336 ) );
  AOI222X4 \us23/U61  ( .A0(\us23/n59 ), .A1(\us23/n43 ), .B0(\us23/n6 ), .B1(
        \us23/n221 ), .C0(\us23/n222 ), .C1(\us23/n187 ), .Y(\us23/n218 ) );
  AOI222X4 \us23/U60  ( .A0(\us23/n123 ), .A1(\us23/n43 ), .B0(sa23[2]), .B1(
        \us23/n203 ), .C0(\us23/n6 ), .C1(\us23/n71 ), .Y(\us23/n202 ) );
  AOI221X4 \us23/U59  ( .A0(\us23/n314 ), .A1(\us23/n43 ), .B0(\us23/n160 ), 
        .B1(\us23/n24 ), .C0(\us23/n315 ), .Y(\us23/n307 ) );
  AOI221X4 \us23/U58  ( .A0(\us23/n43 ), .A1(\us23/n208 ), .B0(\us23/n76 ), 
        .B1(\us23/n24 ), .C0(\us23/n209 ), .Y(\us23/n207 ) );
  AOI221X4 \us23/U57  ( .A0(\us23/n43 ), .A1(\us23/n205 ), .B0(\us23/n32 ), 
        .B1(\us23/n6 ), .C0(\us23/n206 ), .Y(\us23/n201 ) );
  AOI221X4 \us23/U56  ( .A0(\us23/n43 ), .A1(\us23/n44 ), .B0(\us23/n45 ), 
        .B1(\us23/n24 ), .C0(\us23/n46 ), .Y(\us23/n9 ) );
  AOI22XL \us23/U55  ( .A0(\us23/n217 ), .A1(\us23/n43 ), .B0(\us23/n33 ), 
        .B1(\us23/n47 ), .Y(\us23/n216 ) );
  AOI22XL \us23/U54  ( .A0(\us23/n98 ), .A1(\us23/n43 ), .B0(\us23/n6 ), .B1(
        \us23/n99 ), .Y(\us23/n97 ) );
  AOI22XL \us23/U53  ( .A0(\us23/n82 ), .A1(\us23/n43 ), .B0(\us23/n83 ), .B1(
        \us23/n24 ), .Y(\us23/n81 ) );
  AOI2BB2XL \us23/U52  ( .B0(\us23/n43 ), .B1(\us23/n94 ), .A0N(\us23/n120 ), 
        .A1N(\us23/n4 ), .Y(\us23/n119 ) );
  AOI222X4 \us23/U51  ( .A0(\us23/n125 ), .A1(\us23/n33 ), .B0(\us23/n145 ), 
        .B1(\us23/n40 ), .C0(\us23/n43 ), .C1(\us23/n184 ), .Y(\us23/n183 ) );
  AOI22XL \us23/U50  ( .A0(\us23/n43 ), .A1(\us23/n303 ), .B0(\us23/n24 ), 
        .B1(\us23/n96 ), .Y(\us23/n358 ) );
  AOI22XL \us23/U49  ( .A0(\us23/n43 ), .A1(\us23/n100 ), .B0(\us23/n24 ), 
        .B1(\us23/n125 ), .Y(\us23/n124 ) );
  AOI21XL \us23/U48  ( .A0(\us23/n159 ), .A1(\us23/n43 ), .B0(\us23/n40 ), .Y(
        \us23/n262 ) );
  AOI22XL \us23/U47  ( .A0(\us23/n40 ), .A1(\us23/n94 ), .B0(\us23/n43 ), .B1(
        \us23/n187 ), .Y(\us23/n244 ) );
  AOI22XL \us23/U46  ( .A0(\us23/n184 ), .A1(\us23/n5 ), .B0(\us23/n198 ), 
        .B1(\us23/n43 ), .Y(\us23/n197 ) );
  NOR2XL \us23/U45  ( .A(\us23/n33 ), .B(\us23/n2 ), .Y(\us23/n302 ) );
  MXI2XL \us23/U44  ( .A(\us23/n2 ), .B(\us23/n6 ), .S0(\us23/n28 ), .Y(
        \us23/n311 ) );
  INVXL \us23/U43  ( .A(\us23/n20 ), .Y(\us23/n2 ) );
  INVX4 \us23/U42  ( .A(\us23/n6 ), .Y(\us23/n18 ) );
  AOI21XL \us23/U41  ( .A0(\us23/n18 ), .A1(\us23/n162 ), .B0(\us23/n25 ), .Y(
        \us23/n161 ) );
  INVX4 \us23/U40  ( .A(sa23[2]), .Y(\us23/n69 ) );
  NOR2X4 \us23/U39  ( .A(\us23/n226 ), .B(\us23/n4 ), .Y(\us23/n40 ) );
  CLKINVX3 \us23/U38  ( .A(sa23[3]), .Y(\us23/n136 ) );
  NOR2X2 \us23/U37  ( .A(\us23/n136 ), .B(sa23[4]), .Y(\us23/n145 ) );
  CLKINVX3 \us23/U36  ( .A(sa23[4]), .Y(\us23/n58 ) );
  NOR2X2 \us23/U35  ( .A(\us23/n58 ), .B(sa23[3]), .Y(\us23/n159 ) );
  NOR2X2 \us23/U34  ( .A(\us23/n136 ), .B(\us23/n58 ), .Y(\us23/n259 ) );
  NOR2X2 \us23/U33  ( .A(sa23[4]), .B(sa23[3]), .Y(\us23/n278 ) );
  NOR2X2 \us23/U32  ( .A(\us23/n259 ), .B(\us23/n278 ), .Y(\us23/n47 ) );
  CLKINVX3 \us23/U31  ( .A(\us23/n259 ), .Y(\us23/n44 ) );
  NOR2X2 \us23/U30  ( .A(\us23/n44 ), .B(sa23[1]), .Y(\us23/n137 ) );
  AOI21XL \us23/U29  ( .A0(\us23/n44 ), .A1(\us23/n111 ), .B0(\us23/n4 ), .Y(
        \us23/n177 ) );
  AOI22XL \us23/U28  ( .A0(\us23/n23 ), .A1(\us23/n24 ), .B0(\us23/n25 ), .B1(
        sa23[2]), .Y(\us23/n22 ) );
  AOI22XL \us23/U27  ( .A0(\us23/n33 ), .A1(sa23[3]), .B0(\us23/n24 ), .B1(
        \us23/n58 ), .Y(\us23/n277 ) );
  NAND2XL \us23/U26  ( .A(\us23/n198 ), .B(\us23/n24 ), .Y(\us23/n132 ) );
  OAI2BB2XL \us23/U25  ( .B0(\us23/n20 ), .B1(\us23/n111 ), .A0N(\us23/n125 ), 
        .A1N(\us23/n24 ), .Y(\us23/n220 ) );
  NAND2XL \us23/U24  ( .A(\us23/n111 ), .B(\us23/n101 ), .Y(\us23/n21 ) );
  NAND2XL \us23/U23  ( .A(\us23/n111 ), .B(\us23/n300 ), .Y(\us23/n187 ) );
  NAND2XL \us23/U22  ( .A(\us23/n111 ), .B(\us23/n121 ), .Y(\us23/n303 ) );
  AOI221XL \us23/U21  ( .A0(\us23/n43 ), .A1(\us23/n151 ), .B0(\us23/n25 ), 
        .B1(\us23/n69 ), .C0(\us23/n275 ), .Y(\us23/n274 ) );
  NOR2BXL \us23/U20  ( .AN(\us23/n101 ), .B(\us23/n25 ), .Y(\us23/n172 ) );
  NAND2X2 \us23/U19  ( .A(\us23/n58 ), .B(\us23/n226 ), .Y(\us23/n34 ) );
  OAI222X1 \us23/U18  ( .A0(\us23/n27 ), .A1(\us23/n34 ), .B0(\us23/n69 ), 
        .B1(\us23/n205 ), .C0(\us23/n20 ), .C1(\us23/n79 ), .Y(\us23/n260 ) );
  OAI222X1 \us23/U17  ( .A0(\us23/n20 ), .A1(\us23/n99 ), .B0(\us23/n27 ), 
        .B1(\us23/n101 ), .C0(\us23/n184 ), .C1(\us23/n4 ), .Y(\us23/n250 ) );
  OAI222X1 \us23/U16  ( .A0(\us23/n4 ), .A1(\us23/n37 ), .B0(\us23/n38 ), .B1(
        \us23/n20 ), .C0(sa23[4]), .C1(\us23/n39 ), .Y(\us23/n35 ) );
  AOI221X1 \us23/U15  ( .A0(\us23/n5 ), .A1(\us23/n19 ), .B0(\us23/n33 ), .B1(
        \us23/n34 ), .C0(\us23/n35 ), .Y(\us23/n11 ) );
  OR2X2 \us23/U14  ( .A(sa23[2]), .B(sa23[7]), .Y(\us23/n1 ) );
  AOI221XL \us23/U13  ( .A0(\us23/n59 ), .A1(\us23/n33 ), .B0(\us23/n43 ), 
        .B1(\us23/n126 ), .C0(\us23/n127 ), .Y(\us23/n113 ) );
  AOI221XL \us23/U12  ( .A0(\us23/n70 ), .A1(\us23/n43 ), .B0(\us23/n24 ), 
        .B1(\us23/n71 ), .C0(\us23/n72 ), .Y(\us23/n53 ) );
  AOI221X1 \us23/U11  ( .A0(\us23/n313 ), .A1(\us23/n5 ), .B0(\us23/n23 ), 
        .B1(\us23/n2 ), .C0(\us23/n328 ), .Y(\us23/n320 ) );
  AOI222XL \us23/U10  ( .A0(\us23/n185 ), .A1(\us23/n43 ), .B0(\us23/n186 ), 
        .B1(\us23/n187 ), .C0(\us23/n6 ), .C1(\us23/n188 ), .Y(\us23/n164 ) );
  AOI221X1 \us23/U9  ( .A0(\us23/n40 ), .A1(\us23/n136 ), .B0(\us23/n33 ), 
        .B1(\us23/n178 ), .C0(\us23/n338 ), .Y(\us23/n337 ) );
  AOI222XL \us23/U8  ( .A0(\us23/n278 ), .A1(\us23/n24 ), .B0(\us23/n42 ), 
        .B1(\us23/n33 ), .C0(\us23/n43 ), .C1(\us23/n136 ), .Y(\us23/n351 ) );
  AOI31X1 \us23/U7  ( .A0(sa23[2]), .A1(\us23/n58 ), .A2(sa23[1]), .B0(
        \us23/n40 ), .Y(\us23/n350 ) );
  AOI31X1 \us23/U6  ( .A0(\us23/n44 ), .A1(\us23/n129 ), .A2(\us23/n130 ), 
        .B0(\us23/n131 ), .Y(\us23/n128 ) );
  AOI221X1 \us23/U5  ( .A0(\us23/n278 ), .A1(\us23/n40 ), .B0(\us23/n185 ), 
        .B1(\us23/n2 ), .C0(\us23/n279 ), .Y(\us23/n273 ) );
  OAI32X1 \us23/U4  ( .A0(\us23/n18 ), .A1(sa23[1]), .A2(\us23/n159 ), .B0(
        sa23[4]), .B1(\us23/n182 ), .Y(\us23/n318 ) );
  AOI221X1 \us23/U3  ( .A0(\us23/n40 ), .A1(\us23/n136 ), .B0(\us23/n33 ), 
        .B1(\us23/n47 ), .C0(\us23/n156 ), .Y(\us23/n141 ) );
  OAI32X1 \us23/U2  ( .A0(\us23/n210 ), .A1(\us23/n145 ), .A2(\us23/n18 ), 
        .B0(\us23/n27 ), .B1(\us23/n211 ), .Y(\us23/n209 ) );
  AOI31XL \us23/U1  ( .A0(\us23/n79 ), .A1(\us23/n44 ), .A2(\us23/n2 ), .B0(
        \us23/n280 ), .Y(\us23/n339 ) );
  NAND2X1 \us30/U366  ( .A(\us30/n47 ), .B(\us30/n226 ), .Y(\us30/n189 ) );
  NOR2X1 \us30/U365  ( .A(\us30/n226 ), .B(sa30[3]), .Y(\us30/n242 ) );
  INVX1 \us30/U364  ( .A(\us30/n242 ), .Y(\us30/n205 ) );
  AND2X1 \us30/U363  ( .A(\us30/n189 ), .B(\us30/n205 ), .Y(\us30/n65 ) );
  NOR2X1 \us30/U362  ( .A(\us30/n226 ), .B(\us30/n47 ), .Y(\us30/n45 ) );
  NOR2X1 \us30/U361  ( .A(\us30/n259 ), .B(\us30/n45 ), .Y(\us30/n73 ) );
  NAND2BX1 \us30/U360  ( .AN(\us30/n73 ), .B(\us30/n6 ), .Y(\us30/n158 ) );
  NOR2X1 \us30/U359  ( .A(\us30/n226 ), .B(\us30/n159 ), .Y(\us30/n95 ) );
  INVX1 \us30/U358  ( .A(\us30/n95 ), .Y(\us30/n111 ) );
  NOR2X1 \us30/U357  ( .A(\us30/n145 ), .B(sa30[1]), .Y(\us30/n42 ) );
  INVX1 \us30/U356  ( .A(\us30/n42 ), .Y(\us30/n121 ) );
  INVX1 \us30/U355  ( .A(\us30/n47 ), .Y(\us30/n96 ) );
  OAI211X1 \us30/U354  ( .A0(\us30/n65 ), .A1(\us30/n27 ), .B0(\us30/n158 ), 
        .C0(\us30/n358 ), .Y(\us30/n355 ) );
  NOR2X1 \us30/U353  ( .A(\us30/n226 ), .B(\us30/n145 ), .Y(\us30/n59 ) );
  NOR2X1 \us30/U352  ( .A(\us30/n96 ), .B(\us30/n59 ), .Y(\us30/n271 ) );
  NOR2X1 \us30/U351  ( .A(\us30/n226 ), .B(\us30/n278 ), .Y(\us30/n217 ) );
  INVX1 \us30/U350  ( .A(\us30/n217 ), .Y(\us30/n150 ) );
  NAND2X1 \us30/U349  ( .A(\us30/n44 ), .B(\us30/n150 ), .Y(\us30/n147 ) );
  NAND2X1 \us30/U348  ( .A(sa30[4]), .B(\us30/n226 ), .Y(\us30/n101 ) );
  INVX1 \us30/U347  ( .A(\us30/n159 ), .Y(\us30/n188 ) );
  NOR2X1 \us30/U346  ( .A(\us30/n188 ), .B(\us30/n226 ), .Y(\us30/n25 ) );
  INVX1 \us30/U345  ( .A(\us30/n172 ), .Y(\us30/n107 ) );
  AOI22X1 \us30/U344  ( .A0(\us30/n33 ), .A1(\us30/n147 ), .B0(\us30/n24 ), 
        .B1(\us30/n107 ), .Y(\us30/n357 ) );
  OAI221XL \us30/U343  ( .A0(\us30/n18 ), .A1(\us30/n121 ), .B0(\us30/n271 ), 
        .B1(\us30/n20 ), .C0(\us30/n357 ), .Y(\us30/n356 ) );
  MXI2X1 \us30/U342  ( .A(\us30/n355 ), .B(\us30/n356 ), .S0(\us30/n252 ), .Y(
        \us30/n331 ) );
  INVX1 \us30/U341  ( .A(\us30/n59 ), .Y(\us30/n79 ) );
  AND2X1 \us30/U340  ( .A(\us30/n101 ), .B(\us30/n79 ), .Y(\us30/n325 ) );
  XNOR2X1 \us30/U339  ( .A(sa30[5]), .B(\us30/n226 ), .Y(\us30/n352 ) );
  NOR2X1 \us30/U338  ( .A(\us30/n226 ), .B(\us30/n136 ), .Y(\us30/n281 ) );
  INVX1 \us30/U337  ( .A(\us30/n281 ), .Y(\us30/n19 ) );
  NAND2X1 \us30/U336  ( .A(\us30/n145 ), .B(\us30/n226 ), .Y(\us30/n223 ) );
  AOI21X1 \us30/U335  ( .A0(\us30/n19 ), .A1(\us30/n223 ), .B0(\us30/n27 ), 
        .Y(\us30/n354 ) );
  AOI31X1 \us30/U334  ( .A0(\us30/n6 ), .A1(\us30/n352 ), .A2(\us30/n259 ), 
        .B0(\us30/n354 ), .Y(\us30/n353 ) );
  OAI221XL \us30/U333  ( .A0(\us30/n20 ), .A1(\us30/n34 ), .B0(\us30/n325 ), 
        .B1(\us30/n4 ), .C0(\us30/n353 ), .Y(\us30/n347 ) );
  INVX1 \us30/U332  ( .A(\us30/n352 ), .Y(\us30/n349 ) );
  NAND2X1 \us30/U331  ( .A(\us30/n278 ), .B(\us30/n6 ), .Y(\us30/n74 ) );
  OAI211X1 \us30/U330  ( .A0(\us30/n349 ), .A1(\us30/n74 ), .B0(\us30/n350 ), 
        .C0(\us30/n351 ), .Y(\us30/n348 ) );
  MXI2X1 \us30/U329  ( .A(\us30/n347 ), .B(\us30/n348 ), .S0(\us30/n252 ), .Y(
        \us30/n332 ) );
  NOR2X1 \us30/U328  ( .A(\us30/n44 ), .B(\us30/n226 ), .Y(\us30/n157 ) );
  INVX1 \us30/U327  ( .A(\us30/n157 ), .Y(\us30/n240 ) );
  NAND2X1 \us30/U326  ( .A(\us30/n240 ), .B(\us30/n189 ), .Y(\us30/n68 ) );
  NOR2X1 \us30/U325  ( .A(\us30/n20 ), .B(\us30/n159 ), .Y(\us30/n225 ) );
  NOR2X1 \us30/U324  ( .A(\us30/n225 ), .B(\us30/n40 ), .Y(\us30/n345 ) );
  INVX1 \us30/U323  ( .A(\us30/n278 ), .Y(\us30/n94 ) );
  NAND2X1 \us30/U322  ( .A(\us30/n94 ), .B(\us30/n226 ), .Y(\us30/n199 ) );
  NAND2X1 \us30/U321  ( .A(\us30/n199 ), .B(\us30/n205 ), .Y(\us30/n82 ) );
  NAND2X1 \us30/U320  ( .A(\us30/n19 ), .B(\us30/n199 ), .Y(\us30/n295 ) );
  NOR2X1 \us30/U319  ( .A(\us30/n226 ), .B(\us30/n259 ), .Y(\us30/n210 ) );
  NOR2X1 \us30/U318  ( .A(\us30/n27 ), .B(\us30/n210 ), .Y(\us30/n173 ) );
  MXI2X1 \us30/U317  ( .A(\us30/n345 ), .B(\us30/n346 ), .S0(\us30/n252 ), .Y(
        \us30/n342 ) );
  NOR2X1 \us30/U316  ( .A(sa30[1]), .B(sa30[3]), .Y(\us30/n163 ) );
  INVX1 \us30/U315  ( .A(\us30/n163 ), .Y(\us30/n37 ) );
  INVX1 \us30/U314  ( .A(\us30/n173 ), .Y(\us30/n344 ) );
  AOI21X1 \us30/U313  ( .A0(\us30/n240 ), .A1(\us30/n37 ), .B0(\us30/n344 ), 
        .Y(\us30/n343 ) );
  AOI211X1 \us30/U312  ( .A0(\us30/n5 ), .A1(\us30/n68 ), .B0(\us30/n342 ), 
        .C0(\us30/n343 ), .Y(\us30/n333 ) );
  NOR2X1 \us30/U311  ( .A(\us30/n18 ), .B(\us30/n226 ), .Y(\us30/n258 ) );
  NAND2X1 \us30/U310  ( .A(\us30/n278 ), .B(sa30[1]), .Y(\us30/n204 ) );
  NOR2X1 \us30/U309  ( .A(\us30/n188 ), .B(sa30[1]), .Y(\us30/n179 ) );
  INVX1 \us30/U308  ( .A(\us30/n179 ), .Y(\us30/n330 ) );
  NAND2X1 \us30/U307  ( .A(\us30/n204 ), .B(\us30/n330 ), .Y(\us30/n239 ) );
  NOR2X1 \us30/U306  ( .A(\us30/n136 ), .B(sa30[1]), .Y(\us30/n299 ) );
  NOR2X1 \us30/U305  ( .A(\us30/n299 ), .B(\us30/n210 ), .Y(\us30/n341 ) );
  OAI32X1 \us30/U304  ( .A0(\us30/n27 ), .A1(\us30/n278 ), .A2(\us30/n95 ), 
        .B0(\us30/n341 ), .B1(\us30/n4 ), .Y(\us30/n340 ) );
  INVX1 \us30/U303  ( .A(\us30/n45 ), .Y(\us30/n126 ) );
  NAND2X1 \us30/U302  ( .A(\us30/n126 ), .B(\us30/n101 ), .Y(\us30/n178 ) );
  NOR2X1 \us30/U301  ( .A(\us30/n18 ), .B(\us30/n136 ), .Y(\us30/n280 ) );
  OAI21XL \us30/U300  ( .A0(\us30/n4 ), .A1(\us30/n121 ), .B0(\us30/n339 ), 
        .Y(\us30/n338 ) );
  MXI2X1 \us30/U299  ( .A(\us30/n336 ), .B(\us30/n337 ), .S0(\us30/n252 ), .Y(
        \us30/n335 ) );
  NOR2X1 \us30/U298  ( .A(\us30/n258 ), .B(\us30/n335 ), .Y(\us30/n334 ) );
  MX4X1 \us30/U297  ( .A(\us30/n331 ), .B(\us30/n332 ), .C(\us30/n333 ), .D(
        \us30/n334 ), .S0(sa30[6]), .S1(\us30/n234 ), .Y(sa31_sr[0]) );
  INVX1 \us30/U296  ( .A(\us30/n299 ), .Y(\us30/n80 ) );
  NOR2X1 \us30/U295  ( .A(\us30/n111 ), .B(\us30/n18 ), .Y(\us30/n269 ) );
  INVX1 \us30/U294  ( .A(\us30/n269 ), .Y(\us30/n75 ) );
  OAI221XL \us30/U293  ( .A0(\us30/n18 ), .A1(\us30/n330 ), .B0(\us30/n20 ), 
        .B1(\us30/n80 ), .C0(\us30/n75 ), .Y(\us30/n329 ) );
  AOI221X1 \us30/U292  ( .A0(\us30/n325 ), .A1(\us30/n33 ), .B0(\us30/n24 ), 
        .B1(\us30/n303 ), .C0(\us30/n329 ), .Y(\us30/n319 ) );
  NOR2X1 \us30/U291  ( .A(\us30/n234 ), .B(sa30[5]), .Y(\us30/n14 ) );
  NOR2X1 \us30/U290  ( .A(\us30/n25 ), .B(\us30/n299 ), .Y(\us30/n313 ) );
  NAND2X1 \us30/U289  ( .A(\us30/n44 ), .B(\us30/n226 ), .Y(\us30/n300 ) );
  AND2X1 \us30/U288  ( .A(\us30/n300 ), .B(\us30/n240 ), .Y(\us30/n23 ) );
  OAI32X1 \us30/U287  ( .A0(\us30/n4 ), .A1(\us30/n145 ), .A2(\us30/n210 ), 
        .B0(\us30/n137 ), .B1(\us30/n27 ), .Y(\us30/n328 ) );
  NOR2X1 \us30/U286  ( .A(sa30[0]), .B(sa30[5]), .Y(\us30/n16 ) );
  INVX1 \us30/U285  ( .A(\us30/n16 ), .Y(\us30/n114 ) );
  INVX1 \us30/U284  ( .A(\us30/n145 ), .Y(\us30/n149 ) );
  NOR2X1 \us30/U283  ( .A(\us30/n47 ), .B(sa30[1]), .Y(\us30/n98 ) );
  INVX1 \us30/U282  ( .A(\us30/n98 ), .Y(\us30/n284 ) );
  OAI21XL \us30/U281  ( .A0(\us30/n69 ), .A1(\us30/n284 ), .B0(\us30/n27 ), 
        .Y(\us30/n327 ) );
  AOI31X1 \us30/U280  ( .A0(\us30/n111 ), .A1(\us30/n149 ), .A2(\us30/n327 ), 
        .B0(\us30/n225 ), .Y(\us30/n326 ) );
  OAI21XL \us30/U279  ( .A0(\us30/n325 ), .A1(\us30/n18 ), .B0(\us30/n326 ), 
        .Y(\us30/n322 ) );
  NAND2X1 \us30/U278  ( .A(\us30/n19 ), .B(\us30/n189 ), .Y(\us30/n71 ) );
  NOR2X1 \us30/U277  ( .A(\us30/n71 ), .B(\us30/n18 ), .Y(\us30/n135 ) );
  AOI21X1 \us30/U276  ( .A0(\us30/n40 ), .A1(sa30[4]), .B0(\us30/n135 ), .Y(
        \us30/n324 ) );
  OAI221XL \us30/U275  ( .A0(\us30/n47 ), .A1(\us30/n27 ), .B0(\us30/n65 ), 
        .B1(\us30/n20 ), .C0(\us30/n324 ), .Y(\us30/n323 ) );
  AOI22X1 \us30/U274  ( .A0(\us30/n55 ), .A1(\us30/n322 ), .B0(\us30/n89 ), 
        .B1(\us30/n323 ), .Y(\us30/n321 ) );
  OAI221XL \us30/U273  ( .A0(\us30/n319 ), .A1(\us30/n52 ), .B0(\us30/n320 ), 
        .B1(\us30/n114 ), .C0(\us30/n321 ), .Y(\us30/n304 ) );
  NOR2X1 \us30/U272  ( .A(\us30/n226 ), .B(\us30/n58 ), .Y(\us30/n290 ) );
  INVX1 \us30/U271  ( .A(\us30/n290 ), .Y(\us30/n200 ) );
  NAND2X1 \us30/U270  ( .A(\us30/n34 ), .B(\us30/n200 ), .Y(\us30/n120 ) );
  INVX1 \us30/U269  ( .A(\us30/n210 ), .Y(\us30/n100 ) );
  OAI221XL \us30/U268  ( .A0(\us30/n20 ), .A1(\us30/n100 ), .B0(sa30[3]), .B1(
        \us30/n4 ), .C0(\us30/n262 ), .Y(\us30/n317 ) );
  INVX1 \us30/U267  ( .A(\us30/n258 ), .Y(\us30/n182 ) );
  AOI211X1 \us30/U266  ( .A0(\us30/n33 ), .A1(\us30/n120 ), .B0(\us30/n317 ), 
        .C0(\us30/n318 ), .Y(\us30/n306 ) );
  NAND2X1 \us30/U265  ( .A(\us30/n100 ), .B(\us30/n199 ), .Y(\us30/n151 ) );
  INVX1 \us30/U264  ( .A(\us30/n151 ), .Y(\us30/n314 ) );
  NOR2X1 \us30/U263  ( .A(\us30/n45 ), .B(\us30/n163 ), .Y(\us30/n160 ) );
  INVX1 \us30/U262  ( .A(\us30/n295 ), .Y(\us30/n92 ) );
  AOI21X1 \us30/U261  ( .A0(sa30[1]), .A1(\us30/n58 ), .B0(\us30/n98 ), .Y(
        \us30/n316 ) );
  OAI22X1 \us30/U260  ( .A0(\us30/n92 ), .A1(\us30/n18 ), .B0(\us30/n316 ), 
        .B1(\us30/n27 ), .Y(\us30/n315 ) );
  NOR2X1 \us30/U259  ( .A(\us30/n149 ), .B(\us30/n226 ), .Y(\us30/n41 ) );
  INVX1 \us30/U258  ( .A(\us30/n41 ), .Y(\us30/n105 ) );
  NAND2X1 \us30/U257  ( .A(\us30/n284 ), .B(\us30/n105 ), .Y(\us30/n227 ) );
  AOI21X1 \us30/U256  ( .A0(\us30/n313 ), .A1(\us30/n33 ), .B0(\us30/n269 ), 
        .Y(\us30/n312 ) );
  OAI221XL \us30/U255  ( .A0(\us30/n149 ), .A1(\us30/n20 ), .B0(\us30/n4 ), 
        .B1(\us30/n227 ), .C0(\us30/n312 ), .Y(\us30/n309 ) );
  AOI21X1 \us30/U254  ( .A0(\us30/n226 ), .A1(\us30/n188 ), .B0(\us30/n242 ), 
        .Y(\us30/n185 ) );
  INVX1 \us30/U253  ( .A(\us30/n185 ), .Y(\us30/n48 ) );
  AND2X1 \us30/U252  ( .A(\us30/n223 ), .B(\us30/n240 ), .Y(\us30/n28 ) );
  OAI221XL \us30/U251  ( .A0(\us30/n27 ), .A1(\us30/n44 ), .B0(\us30/n4 ), 
        .B1(\us30/n48 ), .C0(\us30/n311 ), .Y(\us30/n310 ) );
  AOI22X1 \us30/U250  ( .A0(\us30/n89 ), .A1(\us30/n309 ), .B0(\us30/n55 ), 
        .B1(\us30/n310 ), .Y(\us30/n308 ) );
  OAI221XL \us30/U249  ( .A0(\us30/n306 ), .A1(\us30/n52 ), .B0(\us30/n307 ), 
        .B1(\us30/n114 ), .C0(\us30/n308 ), .Y(\us30/n305 ) );
  MX2X1 \us30/U248  ( .A(\us30/n304 ), .B(\us30/n305 ), .S0(sa30[6]), .Y(
        sa31_sr[1]) );
  INVX1 \us30/U247  ( .A(\us30/n187 ), .Y(\us30/n61 ) );
  MXI2X1 \us30/U246  ( .A(\us30/n303 ), .B(\us30/n61 ), .S0(\us30/n69 ), .Y(
        \us30/n301 ) );
  MXI2X1 \us30/U245  ( .A(\us30/n301 ), .B(\us30/n147 ), .S0(\us30/n302 ), .Y(
        \us30/n285 ) );
  NAND2X1 \us30/U244  ( .A(\us30/n200 ), .B(\us30/n300 ), .Y(\us30/n99 ) );
  INVX1 \us30/U243  ( .A(\us30/n99 ), .Y(\us30/n296 ) );
  NOR2X1 \us30/U242  ( .A(\us30/n299 ), .B(\us30/n242 ), .Y(\us30/n298 ) );
  NAND2X1 \us30/U241  ( .A(sa30[1]), .B(\us30/n47 ), .Y(\us30/n122 ) );
  NOR2X1 \us30/U240  ( .A(\us30/n159 ), .B(\us30/n217 ), .Y(\us30/n198 ) );
  OAI221XL \us30/U239  ( .A0(\us30/n298 ), .A1(\us30/n27 ), .B0(\us30/n20 ), 
        .B1(\us30/n122 ), .C0(\us30/n132 ), .Y(\us30/n297 ) );
  AOI221X1 \us30/U238  ( .A0(\us30/n225 ), .A1(\us30/n226 ), .B0(\us30/n296 ), 
        .B1(\us30/n6 ), .C0(\us30/n297 ), .Y(\us30/n291 ) );
  OAI2BB2X1 \us30/U237  ( .B0(\us30/n27 ), .B1(\us30/n295 ), .A0N(\us30/n34 ), 
        .A1N(\us30/n24 ), .Y(\us30/n293 ) );
  AOI21X1 \us30/U236  ( .A0(\us30/n101 ), .A1(\us30/n150 ), .B0(\us30/n20 ), 
        .Y(\us30/n294 ) );
  AOI211X1 \us30/U235  ( .A0(\us30/n5 ), .A1(\us30/n79 ), .B0(\us30/n293 ), 
        .C0(\us30/n294 ), .Y(\us30/n292 ) );
  INVX1 \us30/U234  ( .A(\us30/n89 ), .Y(\us30/n10 ) );
  OAI22X1 \us30/U233  ( .A0(\us30/n291 ), .A1(\us30/n114 ), .B0(\us30/n292 ), 
        .B1(\us30/n10 ), .Y(\us30/n286 ) );
  INVX1 \us30/U232  ( .A(\us30/n225 ), .Y(\us30/n288 ) );
  NAND2X1 \us30/U231  ( .A(\us30/n200 ), .B(\us30/n284 ), .Y(\us30/n102 ) );
  NOR2X1 \us30/U230  ( .A(\us30/n290 ), .B(\us30/n163 ), .Y(\us30/n184 ) );
  AOI22X1 \us30/U229  ( .A0(\us30/n102 ), .A1(\us30/n69 ), .B0(\us30/n184 ), 
        .B1(\us30/n33 ), .Y(\us30/n289 ) );
  AOI31X1 \us30/U228  ( .A0(\us30/n132 ), .A1(\us30/n288 ), .A2(\us30/n289 ), 
        .B0(\us30/n52 ), .Y(\us30/n287 ) );
  AOI211X1 \us30/U227  ( .A0(\us30/n285 ), .A1(\us30/n55 ), .B0(\us30/n286 ), 
        .C0(\us30/n287 ), .Y(\us30/n263 ) );
  NAND2X1 \us30/U226  ( .A(\us30/n284 ), .B(\us30/n122 ), .Y(\us30/n125 ) );
  NOR2X1 \us30/U225  ( .A(\us30/n199 ), .B(\us30/n4 ), .Y(\us30/n50 ) );
  AOI21X1 \us30/U224  ( .A0(\us30/n200 ), .A1(\us30/n223 ), .B0(\us30/n20 ), 
        .Y(\us30/n283 ) );
  AOI211X1 \us30/U223  ( .A0(\us30/n5 ), .A1(\us30/n125 ), .B0(\us30/n50 ), 
        .C0(\us30/n283 ), .Y(\us30/n282 ) );
  OAI221XL \us30/U222  ( .A0(\us30/n281 ), .A1(\us30/n27 ), .B0(\us30/n4 ), 
        .B1(\us30/n111 ), .C0(\us30/n282 ), .Y(\us30/n265 ) );
  INVX1 \us30/U221  ( .A(\us30/n280 ), .Y(\us30/n247 ) );
  NAND2X1 \us30/U220  ( .A(\us30/n41 ), .B(\us30/n33 ), .Y(\us30/n272 ) );
  OAI221XL \us30/U219  ( .A0(sa30[1]), .A1(\us30/n247 ), .B0(\us30/n4 ), .B1(
        \us30/n189 ), .C0(\us30/n272 ), .Y(\us30/n279 ) );
  NAND2X1 \us30/U218  ( .A(sa30[2]), .B(\us30/n149 ), .Y(\us30/n276 ) );
  XNOR2X1 \us30/U217  ( .A(\us30/n129 ), .B(sa30[1]), .Y(\us30/n155 ) );
  MXI2X1 \us30/U216  ( .A(\us30/n276 ), .B(\us30/n277 ), .S0(\us30/n155 ), .Y(
        \us30/n275 ) );
  OAI22X1 \us30/U215  ( .A0(\us30/n273 ), .A1(\us30/n10 ), .B0(\us30/n274 ), 
        .B1(\us30/n52 ), .Y(\us30/n266 ) );
  NOR2X1 \us30/U214  ( .A(\us30/n20 ), .B(\us30/n226 ), .Y(\us30/n176 ) );
  OAI21XL \us30/U213  ( .A0(\us30/n4 ), .A1(\us30/n271 ), .B0(\us30/n272 ), 
        .Y(\us30/n270 ) );
  OAI31X1 \us30/U212  ( .A0(\us30/n176 ), .A1(\us30/n269 ), .A2(\us30/n270 ), 
        .B0(\us30/n16 ), .Y(\us30/n268 ) );
  INVX1 \us30/U211  ( .A(\us30/n268 ), .Y(\us30/n267 ) );
  AOI211X1 \us30/U210  ( .A0(\us30/n55 ), .A1(\us30/n265 ), .B0(\us30/n266 ), 
        .C0(\us30/n267 ), .Y(\us30/n264 ) );
  MXI2X1 \us30/U209  ( .A(\us30/n263 ), .B(\us30/n264 ), .S0(sa30[6]), .Y(
        sa31_sr[2]) );
  NOR2X1 \us30/U208  ( .A(\us30/n94 ), .B(sa30[1]), .Y(\us30/n211 ) );
  INVX1 \us30/U207  ( .A(\us30/n262 ), .Y(\us30/n261 ) );
  AOI211X1 \us30/U206  ( .A0(\us30/n259 ), .A1(\us30/n24 ), .B0(\us30/n260 ), 
        .C0(\us30/n261 ), .Y(\us30/n255 ) );
  OAI22X1 \us30/U205  ( .A0(\us30/n20 ), .A1(\us30/n68 ), .B0(\us30/n27 ), 
        .B1(\us30/n37 ), .Y(\us30/n257 ) );
  NOR3X1 \us30/U204  ( .A(\us30/n257 ), .B(\us30/n258 ), .C(\us30/n50 ), .Y(
        \us30/n256 ) );
  MXI2X1 \us30/U203  ( .A(\us30/n255 ), .B(\us30/n256 ), .S0(\us30/n252 ), .Y(
        \us30/n254 ) );
  AOI221X1 \us30/U202  ( .A0(\us30/n211 ), .A1(\us30/n5 ), .B0(\us30/n40 ), 
        .B1(sa30[4]), .C0(\us30/n254 ), .Y(\us30/n248 ) );
  INVX1 \us30/U201  ( .A(\us30/n211 ), .Y(\us30/n106 ) );
  NAND2X1 \us30/U200  ( .A(\us30/n200 ), .B(\us30/n106 ), .Y(\us30/n83 ) );
  NAND2X1 \us30/U199  ( .A(\us30/n199 ), .B(\us30/n204 ), .Y(\us30/n169 ) );
  AOI2BB2X1 \us30/U198  ( .B0(\us30/n65 ), .B1(\us30/n24 ), .A0N(\us30/n169 ), 
        .A1N(\us30/n20 ), .Y(\us30/n253 ) );
  OAI221XL \us30/U197  ( .A0(\us30/n172 ), .A1(\us30/n18 ), .B0(\us30/n27 ), 
        .B1(\us30/n83 ), .C0(\us30/n253 ), .Y(\us30/n251 ) );
  MXI2X1 \us30/U196  ( .A(\us30/n250 ), .B(\us30/n251 ), .S0(\us30/n252 ), .Y(
        \us30/n249 ) );
  MXI2X1 \us30/U195  ( .A(\us30/n248 ), .B(\us30/n249 ), .S0(\us30/n234 ), .Y(
        \us30/n228 ) );
  OAI21XL \us30/U194  ( .A0(\us30/n58 ), .A1(\us30/n27 ), .B0(\us30/n247 ), 
        .Y(\us30/n245 ) );
  NOR2X1 \us30/U193  ( .A(sa30[7]), .B(\us30/n145 ), .Y(\us30/n246 ) );
  XNOR2X1 \us30/U192  ( .A(\us30/n69 ), .B(sa30[1]), .Y(\us30/n130 ) );
  MXI2X1 \us30/U191  ( .A(\us30/n245 ), .B(\us30/n246 ), .S0(\us30/n130 ), .Y(
        \us30/n243 ) );
  OAI211X1 \us30/U190  ( .A0(\us30/n4 ), .A1(\us30/n149 ), .B0(\us30/n243 ), 
        .C0(\us30/n244 ), .Y(\us30/n230 ) );
  NOR2X1 \us30/U189  ( .A(\us30/n242 ), .B(\us30/n137 ), .Y(\us30/n70 ) );
  OAI221XL \us30/U188  ( .A0(\us30/n159 ), .A1(\us30/n27 ), .B0(\us30/n20 ), 
        .B1(\us30/n34 ), .C0(\us30/n241 ), .Y(\us30/n231 ) );
  NAND2X1 \us30/U187  ( .A(\us30/n101 ), .B(\us30/n240 ), .Y(\us30/n76 ) );
  AOI21X1 \us30/U186  ( .A0(\us30/n122 ), .A1(\us30/n106 ), .B0(\us30/n129 ), 
        .Y(\us30/n237 ) );
  INVX1 \us30/U185  ( .A(\us30/n239 ), .Y(\us30/n238 ) );
  OAI21XL \us30/U184  ( .A0(\us30/n237 ), .A1(\us30/n43 ), .B0(\us30/n238 ), 
        .Y(\us30/n236 ) );
  OAI221XL \us30/U183  ( .A0(\us30/n18 ), .A1(\us30/n76 ), .B0(\us30/n59 ), 
        .B1(\us30/n27 ), .C0(\us30/n236 ), .Y(\us30/n232 ) );
  AOI2BB2X1 \us30/U182  ( .B0(\us30/n24 ), .B1(\us30/n187 ), .A0N(\us30/n227 ), 
        .A1N(\us30/n20 ), .Y(\us30/n235 ) );
  OAI211X1 \us30/U181  ( .A0(\us30/n27 ), .A1(\us30/n122 ), .B0(\us30/n158 ), 
        .C0(\us30/n235 ), .Y(\us30/n233 ) );
  MX4X1 \us30/U180  ( .A(\us30/n230 ), .B(\us30/n231 ), .C(\us30/n232 ), .D(
        \us30/n233 ), .S0(\us30/n234 ), .S1(sa30[5]), .Y(\us30/n229 ) );
  MX2X1 \us30/U179  ( .A(\us30/n228 ), .B(\us30/n229 ), .S0(sa30[6]), .Y(
        sa31_sr[3]) );
  NOR2BX1 \us30/U178  ( .AN(\us30/n204 ), .B(\us30/n137 ), .Y(\us30/n110 ) );
  INVX1 \us30/U177  ( .A(\us30/n110 ), .Y(\us30/n64 ) );
  AOI22X1 \us30/U176  ( .A0(\us30/n225 ), .A1(\us30/n226 ), .B0(\us30/n6 ), 
        .B1(\us30/n227 ), .Y(\us30/n224 ) );
  OAI221XL \us30/U175  ( .A0(\us30/n27 ), .A1(\us30/n64 ), .B0(\us30/n4 ), 
        .B1(\us30/n83 ), .C0(\us30/n224 ), .Y(\us30/n212 ) );
  NAND2X1 \us30/U174  ( .A(\us30/n34 ), .B(\us30/n204 ), .Y(\us30/n221 ) );
  OAI21XL \us30/U173  ( .A0(\us30/n69 ), .A1(\us30/n223 ), .B0(\us30/n27 ), 
        .Y(\us30/n222 ) );
  NOR2X1 \us30/U172  ( .A(\us30/n217 ), .B(\us30/n42 ), .Y(\us30/n208 ) );
  AOI211X1 \us30/U171  ( .A0(\us30/n208 ), .A1(\us30/n5 ), .B0(\us30/n220 ), 
        .C0(\us30/n173 ), .Y(\us30/n219 ) );
  OAI22X1 \us30/U170  ( .A0(\us30/n218 ), .A1(\us30/n10 ), .B0(\us30/n219 ), 
        .B1(\us30/n114 ), .Y(\us30/n213 ) );
  INVX1 \us30/U169  ( .A(\us30/n135 ), .Y(\us30/n215 ) );
  NOR2X1 \us30/U168  ( .A(\us30/n4 ), .B(\us30/n159 ), .Y(\us30/n31 ) );
  INVX1 \us30/U167  ( .A(\us30/n31 ), .Y(\us30/n196 ) );
  AOI31X1 \us30/U166  ( .A0(\us30/n215 ), .A1(\us30/n196 ), .A2(\us30/n216 ), 
        .B0(\us30/n52 ), .Y(\us30/n214 ) );
  AOI211X1 \us30/U165  ( .A0(\us30/n55 ), .A1(\us30/n212 ), .B0(\us30/n213 ), 
        .C0(\us30/n214 ), .Y(\us30/n190 ) );
  INVX1 \us30/U164  ( .A(\us30/n207 ), .Y(\us30/n192 ) );
  NOR2X1 \us30/U163  ( .A(\us30/n25 ), .B(\us30/n98 ), .Y(\us30/n32 ) );
  OAI22X1 \us30/U162  ( .A0(\us30/n28 ), .A1(\us30/n4 ), .B0(\us30/n188 ), 
        .B1(\us30/n27 ), .Y(\us30/n206 ) );
  NAND2X1 \us30/U161  ( .A(\us30/n204 ), .B(\us30/n80 ), .Y(\us30/n118 ) );
  INVX1 \us30/U160  ( .A(\us30/n118 ), .Y(\us30/n123 ) );
  NAND2X1 \us30/U159  ( .A(\us30/n94 ), .B(\us30/n79 ), .Y(\us30/n203 ) );
  OAI2BB1X1 \us30/U158  ( .A0N(\us30/n199 ), .A1N(\us30/n200 ), .B0(\us30/n33 ), .Y(\us30/n195 ) );
  INVX1 \us30/U157  ( .A(\us30/n55 ), .Y(\us30/n12 ) );
  AOI31X1 \us30/U156  ( .A0(\us30/n195 ), .A1(\us30/n196 ), .A2(\us30/n197 ), 
        .B0(\us30/n12 ), .Y(\us30/n194 ) );
  AOI211X1 \us30/U155  ( .A0(\us30/n89 ), .A1(\us30/n192 ), .B0(\us30/n193 ), 
        .C0(\us30/n194 ), .Y(\us30/n191 ) );
  MXI2X1 \us30/U154  ( .A(\us30/n190 ), .B(\us30/n191 ), .S0(sa30[6]), .Y(
        sa31_sr[4]) );
  OAI21XL \us30/U153  ( .A0(\us30/n69 ), .A1(\us30/n189 ), .B0(\us30/n27 ), 
        .Y(\us30/n186 ) );
  INVX1 \us30/U152  ( .A(\us30/n183 ), .Y(\us30/n180 ) );
  NAND2X1 \us30/U151  ( .A(\us30/n74 ), .B(\us30/n182 ), .Y(\us30/n181 ) );
  AOI211X1 \us30/U150  ( .A0(\us30/n179 ), .A1(\us30/n24 ), .B0(\us30/n180 ), 
        .C0(\us30/n181 ), .Y(\us30/n165 ) );
  INVX1 \us30/U149  ( .A(\us30/n178 ), .Y(\us30/n175 ) );
  AOI211X1 \us30/U148  ( .A0(\us30/n175 ), .A1(\us30/n5 ), .B0(\us30/n176 ), 
        .C0(\us30/n177 ), .Y(\us30/n174 ) );
  OAI221XL \us30/U147  ( .A0(\us30/n159 ), .A1(\us30/n27 ), .B0(\us30/n145 ), 
        .B1(\us30/n20 ), .C0(\us30/n174 ), .Y(\us30/n167 ) );
  MXI2X1 \us30/U146  ( .A(\us30/n40 ), .B(\us30/n173 ), .S0(\us30/n96 ), .Y(
        \us30/n170 ) );
  AOI22X1 \us30/U145  ( .A0(\us30/n137 ), .A1(\us30/n24 ), .B0(\us30/n172 ), 
        .B1(\us30/n6 ), .Y(\us30/n171 ) );
  OAI211X1 \us30/U144  ( .A0(\us30/n20 ), .A1(\us30/n169 ), .B0(\us30/n170 ), 
        .C0(\us30/n171 ), .Y(\us30/n168 ) );
  AOI22X1 \us30/U143  ( .A0(\us30/n89 ), .A1(\us30/n167 ), .B0(\us30/n55 ), 
        .B1(\us30/n168 ), .Y(\us30/n166 ) );
  OAI221XL \us30/U142  ( .A0(\us30/n164 ), .A1(\us30/n114 ), .B0(\us30/n165 ), 
        .B1(\us30/n52 ), .C0(\us30/n166 ), .Y(\us30/n138 ) );
  OAI21XL \us30/U141  ( .A0(\us30/n41 ), .A1(\us30/n163 ), .B0(\us30/n69 ), 
        .Y(\us30/n162 ) );
  AOI221X1 \us30/U140  ( .A0(\us30/n159 ), .A1(\us30/n24 ), .B0(\us30/n160 ), 
        .B1(\us30/n33 ), .C0(\us30/n161 ), .Y(\us30/n140 ) );
  OAI21XL \us30/U139  ( .A0(\us30/n157 ), .A1(\us30/n20 ), .B0(\us30/n158 ), 
        .Y(\us30/n156 ) );
  NOR2X1 \us30/U138  ( .A(\us30/n4 ), .B(\us30/n136 ), .Y(\us30/n153 ) );
  NOR2X1 \us30/U137  ( .A(\us30/n145 ), .B(\us30/n69 ), .Y(\us30/n154 ) );
  MXI2X1 \us30/U136  ( .A(\us30/n153 ), .B(\us30/n154 ), .S0(\us30/n155 ), .Y(
        \us30/n152 ) );
  OAI221XL \us30/U135  ( .A0(\us30/n110 ), .A1(\us30/n18 ), .B0(\us30/n20 ), 
        .B1(\us30/n151 ), .C0(\us30/n152 ), .Y(\us30/n143 ) );
  AOI21X1 \us30/U134  ( .A0(\us30/n149 ), .A1(\us30/n150 ), .B0(\us30/n18 ), 
        .Y(\us30/n148 ) );
  AOI2BB1X1 \us30/U133  ( .A0N(\us30/n147 ), .A1N(\us30/n27 ), .B0(\us30/n148 ), .Y(\us30/n146 ) );
  OAI221XL \us30/U132  ( .A0(\us30/n145 ), .A1(\us30/n20 ), .B0(\us30/n4 ), 
        .B1(\us30/n34 ), .C0(\us30/n146 ), .Y(\us30/n144 ) );
  AOI22X1 \us30/U131  ( .A0(\us30/n89 ), .A1(\us30/n143 ), .B0(\us30/n14 ), 
        .B1(\us30/n144 ), .Y(\us30/n142 ) );
  OAI221XL \us30/U130  ( .A0(\us30/n140 ), .A1(\us30/n12 ), .B0(\us30/n141 ), 
        .B1(\us30/n114 ), .C0(\us30/n142 ), .Y(\us30/n139 ) );
  MX2X1 \us30/U129  ( .A(\us30/n138 ), .B(\us30/n139 ), .S0(sa30[6]), .Y(
        sa31_sr[5]) );
  INVX1 \us30/U128  ( .A(\us30/n70 ), .Y(\us30/n133 ) );
  OAI22X1 \us30/U127  ( .A0(\us30/n4 ), .A1(\us30/n136 ), .B0(\us30/n137 ), 
        .B1(\us30/n27 ), .Y(\us30/n134 ) );
  AOI211X1 \us30/U126  ( .A0(\us30/n133 ), .A1(\us30/n69 ), .B0(\us30/n134 ), 
        .C0(\us30/n135 ), .Y(\us30/n112 ) );
  INVX1 \us30/U125  ( .A(\us30/n132 ), .Y(\us30/n131 ) );
  OAI21XL \us30/U124  ( .A0(\us30/n18 ), .A1(\us30/n37 ), .B0(\us30/n128 ), 
        .Y(\us30/n127 ) );
  OAI221XL \us30/U123  ( .A0(\us30/n18 ), .A1(\us30/n105 ), .B0(\us30/n123 ), 
        .B1(\us30/n27 ), .C0(\us30/n124 ), .Y(\us30/n116 ) );
  NAND2X1 \us30/U122  ( .A(\us30/n121 ), .B(\us30/n122 ), .Y(\us30/n30 ) );
  OAI221XL \us30/U121  ( .A0(\us30/n18 ), .A1(\us30/n118 ), .B0(\us30/n27 ), 
        .B1(\us30/n30 ), .C0(\us30/n119 ), .Y(\us30/n117 ) );
  AOI22X1 \us30/U120  ( .A0(\us30/n89 ), .A1(\us30/n116 ), .B0(\us30/n55 ), 
        .B1(\us30/n117 ), .Y(\us30/n115 ) );
  OAI221XL \us30/U119  ( .A0(\us30/n112 ), .A1(\us30/n52 ), .B0(\us30/n113 ), 
        .B1(\us30/n114 ), .C0(\us30/n115 ), .Y(\us30/n84 ) );
  OAI22X1 \us30/U118  ( .A0(\us30/n110 ), .A1(\us30/n4 ), .B0(\us30/n20 ), 
        .B1(\us30/n21 ), .Y(\us30/n108 ) );
  AOI21X1 \us30/U117  ( .A0(sa30[1]), .A1(\us30/n58 ), .B0(\us30/n27 ), .Y(
        \us30/n109 ) );
  AOI211X1 \us30/U116  ( .A0(\us30/n5 ), .A1(\us30/n107 ), .B0(\us30/n108 ), 
        .C0(\us30/n109 ), .Y(\us30/n86 ) );
  OAI22X1 \us30/U115  ( .A0(\us30/n45 ), .A1(\us30/n4 ), .B0(sa30[4]), .B1(
        \us30/n18 ), .Y(\us30/n103 ) );
  AOI21X1 \us30/U114  ( .A0(\us30/n105 ), .A1(\us30/n106 ), .B0(\us30/n20 ), 
        .Y(\us30/n104 ) );
  AOI211X1 \us30/U113  ( .A0(\us30/n33 ), .A1(\us30/n102 ), .B0(\us30/n103 ), 
        .C0(\us30/n104 ), .Y(\us30/n87 ) );
  NAND2X1 \us30/U112  ( .A(\us30/n100 ), .B(\us30/n101 ), .Y(\us30/n62 ) );
  OAI221XL \us30/U111  ( .A0(\us30/n27 ), .A1(\us30/n62 ), .B0(\us30/n4 ), 
        .B1(\us30/n21 ), .C0(\us30/n97 ), .Y(\us30/n90 ) );
  NOR3X1 \us30/U110  ( .A(\us30/n4 ), .B(\us30/n95 ), .C(\us30/n96 ), .Y(
        \us30/n67 ) );
  AOI31X1 \us30/U109  ( .A0(\us30/n79 ), .A1(\us30/n94 ), .A2(\us30/n6 ), .B0(
        \us30/n67 ), .Y(\us30/n93 ) );
  OAI221XL \us30/U108  ( .A0(\us30/n73 ), .A1(\us30/n27 ), .B0(\us30/n92 ), 
        .B1(\us30/n20 ), .C0(\us30/n93 ), .Y(\us30/n91 ) );
  AOI22X1 \us30/U107  ( .A0(\us30/n89 ), .A1(\us30/n90 ), .B0(\us30/n16 ), 
        .B1(\us30/n91 ), .Y(\us30/n88 ) );
  OAI221XL \us30/U106  ( .A0(\us30/n86 ), .A1(\us30/n52 ), .B0(\us30/n87 ), 
        .B1(\us30/n12 ), .C0(\us30/n88 ), .Y(\us30/n85 ) );
  MX2X1 \us30/U105  ( .A(\us30/n84 ), .B(\us30/n85 ), .S0(sa30[6]), .Y(
        sa31_sr[6]) );
  INVX1 \us30/U104  ( .A(\us30/n81 ), .Y(\us30/n77 ) );
  AOI21X1 \us30/U103  ( .A0(\us30/n79 ), .A1(\us30/n80 ), .B0(\us30/n27 ), .Y(
        \us30/n78 ) );
  AOI211X1 \us30/U102  ( .A0(\us30/n5 ), .A1(\us30/n76 ), .B0(\us30/n77 ), 
        .C0(\us30/n78 ), .Y(\us30/n51 ) );
  OAI211X1 \us30/U101  ( .A0(\us30/n73 ), .A1(\us30/n27 ), .B0(\us30/n74 ), 
        .C0(\us30/n75 ), .Y(\us30/n72 ) );
  AOI21X1 \us30/U100  ( .A0(\us30/n68 ), .A1(\us30/n69 ), .B0(\us30/n6 ), .Y(
        \us30/n63 ) );
  INVX1 \us30/U99  ( .A(\us30/n67 ), .Y(\us30/n66 ) );
  OAI221XL \us30/U98  ( .A0(\us30/n63 ), .A1(\us30/n64 ), .B0(\us30/n65 ), 
        .B1(\us30/n27 ), .C0(\us30/n66 ), .Y(\us30/n56 ) );
  AOI2BB2X1 \us30/U97  ( .B0(\us30/n61 ), .B1(\us30/n24 ), .A0N(\us30/n62 ), 
        .A1N(\us30/n20 ), .Y(\us30/n60 ) );
  OAI221XL \us30/U96  ( .A0(\us30/n58 ), .A1(\us30/n18 ), .B0(\us30/n59 ), 
        .B1(\us30/n27 ), .C0(\us30/n60 ), .Y(\us30/n57 ) );
  AOI22X1 \us30/U95  ( .A0(\us30/n55 ), .A1(\us30/n56 ), .B0(\us30/n16 ), .B1(
        \us30/n57 ), .Y(\us30/n54 ) );
  OAI221XL \us30/U94  ( .A0(\us30/n51 ), .A1(\us30/n52 ), .B0(\us30/n53 ), 
        .B1(\us30/n10 ), .C0(\us30/n54 ), .Y(\us30/n7 ) );
  INVX1 \us30/U93  ( .A(\us30/n50 ), .Y(\us30/n49 ) );
  OAI221XL \us30/U92  ( .A0(\us30/n47 ), .A1(\us30/n18 ), .B0(\us30/n27 ), 
        .B1(\us30/n48 ), .C0(\us30/n49 ), .Y(\us30/n46 ) );
  NOR2X1 \us30/U91  ( .A(\us30/n41 ), .B(\us30/n42 ), .Y(\us30/n38 ) );
  INVX1 \us30/U90  ( .A(\us30/n40 ), .Y(\us30/n39 ) );
  INVX1 \us30/U89  ( .A(\us30/n32 ), .Y(\us30/n26 ) );
  AOI21X1 \us30/U88  ( .A0(\us30/n5 ), .A1(\us30/n30 ), .B0(\us30/n31 ), .Y(
        \us30/n29 ) );
  OAI221XL \us30/U87  ( .A0(\us30/n26 ), .A1(\us30/n27 ), .B0(\us30/n28 ), 
        .B1(\us30/n20 ), .C0(\us30/n29 ), .Y(\us30/n15 ) );
  OAI221XL \us30/U86  ( .A0(\us30/n18 ), .A1(\us30/n19 ), .B0(\us30/n20 ), 
        .B1(\us30/n21 ), .C0(\us30/n22 ), .Y(\us30/n17 ) );
  AOI22X1 \us30/U85  ( .A0(\us30/n14 ), .A1(\us30/n15 ), .B0(\us30/n16 ), .B1(
        \us30/n17 ), .Y(\us30/n13 ) );
  OAI221XL \us30/U84  ( .A0(\us30/n9 ), .A1(\us30/n10 ), .B0(\us30/n11 ), .B1(
        \us30/n12 ), .C0(\us30/n13 ), .Y(\us30/n8 ) );
  MX2X1 \us30/U83  ( .A(\us30/n7 ), .B(\us30/n8 ), .S0(sa30[6]), .Y(sa31_sr[7]) );
  NOR2X4 \us30/U82  ( .A(\us30/n129 ), .B(sa30[2]), .Y(\us30/n43 ) );
  CLKINVX3 \us30/U81  ( .A(\us30/n14 ), .Y(\us30/n52 ) );
  OAI22XL \us30/U80  ( .A0(\us30/n201 ), .A1(\us30/n52 ), .B0(\us30/n202 ), 
        .B1(\us30/n114 ), .Y(\us30/n193 ) );
  CLKINVX3 \us30/U79  ( .A(sa30[5]), .Y(\us30/n252 ) );
  NOR2X2 \us30/U78  ( .A(\us30/n252 ), .B(\us30/n234 ), .Y(\us30/n55 ) );
  CLKINVX3 \us30/U77  ( .A(sa30[7]), .Y(\us30/n129 ) );
  NOR2X4 \us30/U76  ( .A(\us30/n129 ), .B(\us30/n69 ), .Y(\us30/n24 ) );
  AOI22XL \us30/U75  ( .A0(\us30/n70 ), .A1(\us30/n24 ), .B0(\us30/n96 ), .B1(
        \us30/n129 ), .Y(\us30/n241 ) );
  NOR2X2 \us30/U74  ( .A(\us30/n252 ), .B(sa30[0]), .Y(\us30/n89 ) );
  CLKINVX3 \us30/U73  ( .A(sa30[0]), .Y(\us30/n234 ) );
  NOR2X4 \us30/U72  ( .A(\us30/n69 ), .B(sa30[7]), .Y(\us30/n33 ) );
  INVX12 \us30/U71  ( .A(\us30/n33 ), .Y(\us30/n27 ) );
  CLKINVX3 \us30/U70  ( .A(\us30/n1 ), .Y(\us30/n6 ) );
  CLKINVX3 \us30/U69  ( .A(\us30/n1 ), .Y(\us30/n5 ) );
  INVXL \us30/U68  ( .A(\us30/n24 ), .Y(\us30/n36 ) );
  INVX4 \us30/U67  ( .A(\us30/n3 ), .Y(\us30/n4 ) );
  INVXL \us30/U66  ( .A(\us30/n36 ), .Y(\us30/n3 ) );
  INVX4 \us30/U65  ( .A(sa30[1]), .Y(\us30/n226 ) );
  INVX4 \us30/U64  ( .A(\us30/n43 ), .Y(\us30/n20 ) );
  AOI221X4 \us30/U63  ( .A0(\us30/n24 ), .A1(\us30/n82 ), .B0(\us30/n43 ), 
        .B1(\us30/n295 ), .C0(\us30/n173 ), .Y(\us30/n346 ) );
  AOI221X4 \us30/U62  ( .A0(\us30/n5 ), .A1(\us30/n96 ), .B0(\us30/n43 ), .B1(
        \us30/n239 ), .C0(\us30/n340 ), .Y(\us30/n336 ) );
  AOI222X4 \us30/U61  ( .A0(\us30/n59 ), .A1(\us30/n43 ), .B0(\us30/n6 ), .B1(
        \us30/n221 ), .C0(\us30/n222 ), .C1(\us30/n187 ), .Y(\us30/n218 ) );
  AOI222X4 \us30/U60  ( .A0(\us30/n123 ), .A1(\us30/n43 ), .B0(sa30[2]), .B1(
        \us30/n203 ), .C0(\us30/n6 ), .C1(\us30/n71 ), .Y(\us30/n202 ) );
  AOI221X4 \us30/U59  ( .A0(\us30/n314 ), .A1(\us30/n43 ), .B0(\us30/n160 ), 
        .B1(\us30/n24 ), .C0(\us30/n315 ), .Y(\us30/n307 ) );
  AOI221X4 \us30/U58  ( .A0(\us30/n43 ), .A1(\us30/n208 ), .B0(\us30/n76 ), 
        .B1(\us30/n24 ), .C0(\us30/n209 ), .Y(\us30/n207 ) );
  AOI221X4 \us30/U57  ( .A0(\us30/n43 ), .A1(\us30/n205 ), .B0(\us30/n32 ), 
        .B1(\us30/n6 ), .C0(\us30/n206 ), .Y(\us30/n201 ) );
  AOI221X4 \us30/U56  ( .A0(\us30/n43 ), .A1(\us30/n44 ), .B0(\us30/n45 ), 
        .B1(\us30/n24 ), .C0(\us30/n46 ), .Y(\us30/n9 ) );
  AOI22XL \us30/U55  ( .A0(\us30/n217 ), .A1(\us30/n43 ), .B0(\us30/n33 ), 
        .B1(\us30/n47 ), .Y(\us30/n216 ) );
  AOI22XL \us30/U54  ( .A0(\us30/n98 ), .A1(\us30/n43 ), .B0(\us30/n6 ), .B1(
        \us30/n99 ), .Y(\us30/n97 ) );
  AOI22XL \us30/U53  ( .A0(\us30/n82 ), .A1(\us30/n43 ), .B0(\us30/n83 ), .B1(
        \us30/n24 ), .Y(\us30/n81 ) );
  AOI2BB2XL \us30/U52  ( .B0(\us30/n43 ), .B1(\us30/n94 ), .A0N(\us30/n120 ), 
        .A1N(\us30/n4 ), .Y(\us30/n119 ) );
  AOI222X4 \us30/U51  ( .A0(\us30/n125 ), .A1(\us30/n33 ), .B0(\us30/n145 ), 
        .B1(\us30/n40 ), .C0(\us30/n43 ), .C1(\us30/n184 ), .Y(\us30/n183 ) );
  AOI22XL \us30/U50  ( .A0(\us30/n43 ), .A1(\us30/n303 ), .B0(\us30/n24 ), 
        .B1(\us30/n96 ), .Y(\us30/n358 ) );
  AOI22XL \us30/U49  ( .A0(\us30/n43 ), .A1(\us30/n100 ), .B0(\us30/n24 ), 
        .B1(\us30/n125 ), .Y(\us30/n124 ) );
  AOI21XL \us30/U48  ( .A0(\us30/n159 ), .A1(\us30/n43 ), .B0(\us30/n40 ), .Y(
        \us30/n262 ) );
  AOI22XL \us30/U47  ( .A0(\us30/n40 ), .A1(\us30/n94 ), .B0(\us30/n43 ), .B1(
        \us30/n187 ), .Y(\us30/n244 ) );
  AOI22XL \us30/U46  ( .A0(\us30/n184 ), .A1(\us30/n5 ), .B0(\us30/n198 ), 
        .B1(\us30/n43 ), .Y(\us30/n197 ) );
  NOR2XL \us30/U45  ( .A(\us30/n33 ), .B(\us30/n2 ), .Y(\us30/n302 ) );
  MXI2XL \us30/U44  ( .A(\us30/n2 ), .B(\us30/n6 ), .S0(\us30/n28 ), .Y(
        \us30/n311 ) );
  INVXL \us30/U43  ( .A(\us30/n20 ), .Y(\us30/n2 ) );
  INVX4 \us30/U42  ( .A(\us30/n6 ), .Y(\us30/n18 ) );
  AOI21XL \us30/U41  ( .A0(\us30/n18 ), .A1(\us30/n162 ), .B0(\us30/n25 ), .Y(
        \us30/n161 ) );
  INVX4 \us30/U40  ( .A(sa30[2]), .Y(\us30/n69 ) );
  NOR2X4 \us30/U39  ( .A(\us30/n226 ), .B(\us30/n4 ), .Y(\us30/n40 ) );
  CLKINVX3 \us30/U38  ( .A(sa30[3]), .Y(\us30/n136 ) );
  NOR2X2 \us30/U37  ( .A(\us30/n136 ), .B(sa30[4]), .Y(\us30/n145 ) );
  CLKINVX3 \us30/U36  ( .A(sa30[4]), .Y(\us30/n58 ) );
  NOR2X2 \us30/U35  ( .A(\us30/n58 ), .B(sa30[3]), .Y(\us30/n159 ) );
  NOR2X2 \us30/U34  ( .A(\us30/n136 ), .B(\us30/n58 ), .Y(\us30/n259 ) );
  NOR2X2 \us30/U33  ( .A(sa30[4]), .B(sa30[3]), .Y(\us30/n278 ) );
  NOR2X2 \us30/U32  ( .A(\us30/n259 ), .B(\us30/n278 ), .Y(\us30/n47 ) );
  CLKINVX3 \us30/U31  ( .A(\us30/n259 ), .Y(\us30/n44 ) );
  NOR2X2 \us30/U30  ( .A(\us30/n44 ), .B(sa30[1]), .Y(\us30/n137 ) );
  AOI21XL \us30/U29  ( .A0(\us30/n44 ), .A1(\us30/n111 ), .B0(\us30/n4 ), .Y(
        \us30/n177 ) );
  AOI22XL \us30/U28  ( .A0(\us30/n23 ), .A1(\us30/n24 ), .B0(\us30/n25 ), .B1(
        sa30[2]), .Y(\us30/n22 ) );
  AOI22XL \us30/U27  ( .A0(\us30/n33 ), .A1(sa30[3]), .B0(\us30/n24 ), .B1(
        \us30/n58 ), .Y(\us30/n277 ) );
  NAND2XL \us30/U26  ( .A(\us30/n198 ), .B(\us30/n24 ), .Y(\us30/n132 ) );
  OAI2BB2XL \us30/U25  ( .B0(\us30/n20 ), .B1(\us30/n111 ), .A0N(\us30/n125 ), 
        .A1N(\us30/n24 ), .Y(\us30/n220 ) );
  NAND2XL \us30/U24  ( .A(\us30/n111 ), .B(\us30/n101 ), .Y(\us30/n21 ) );
  NAND2XL \us30/U23  ( .A(\us30/n111 ), .B(\us30/n300 ), .Y(\us30/n187 ) );
  NAND2XL \us30/U22  ( .A(\us30/n111 ), .B(\us30/n121 ), .Y(\us30/n303 ) );
  AOI221XL \us30/U21  ( .A0(\us30/n43 ), .A1(\us30/n151 ), .B0(\us30/n25 ), 
        .B1(\us30/n69 ), .C0(\us30/n275 ), .Y(\us30/n274 ) );
  NOR2BXL \us30/U20  ( .AN(\us30/n101 ), .B(\us30/n25 ), .Y(\us30/n172 ) );
  NAND2X2 \us30/U19  ( .A(\us30/n58 ), .B(\us30/n226 ), .Y(\us30/n34 ) );
  OAI222X1 \us30/U18  ( .A0(\us30/n27 ), .A1(\us30/n34 ), .B0(\us30/n69 ), 
        .B1(\us30/n205 ), .C0(\us30/n20 ), .C1(\us30/n79 ), .Y(\us30/n260 ) );
  OAI222X1 \us30/U17  ( .A0(\us30/n20 ), .A1(\us30/n99 ), .B0(\us30/n27 ), 
        .B1(\us30/n101 ), .C0(\us30/n184 ), .C1(\us30/n4 ), .Y(\us30/n250 ) );
  OAI222X1 \us30/U16  ( .A0(\us30/n4 ), .A1(\us30/n37 ), .B0(\us30/n38 ), .B1(
        \us30/n20 ), .C0(sa30[4]), .C1(\us30/n39 ), .Y(\us30/n35 ) );
  AOI221X1 \us30/U15  ( .A0(\us30/n5 ), .A1(\us30/n19 ), .B0(\us30/n33 ), .B1(
        \us30/n34 ), .C0(\us30/n35 ), .Y(\us30/n11 ) );
  OR2X2 \us30/U14  ( .A(sa30[2]), .B(sa30[7]), .Y(\us30/n1 ) );
  AOI221XL \us30/U13  ( .A0(\us30/n70 ), .A1(\us30/n43 ), .B0(\us30/n24 ), 
        .B1(\us30/n71 ), .C0(\us30/n72 ), .Y(\us30/n53 ) );
  AOI221XL \us30/U12  ( .A0(\us30/n59 ), .A1(\us30/n33 ), .B0(\us30/n43 ), 
        .B1(\us30/n126 ), .C0(\us30/n127 ), .Y(\us30/n113 ) );
  AOI222XL \us30/U11  ( .A0(\us30/n185 ), .A1(\us30/n43 ), .B0(\us30/n186 ), 
        .B1(\us30/n187 ), .C0(\us30/n6 ), .C1(\us30/n188 ), .Y(\us30/n164 ) );
  AOI221X1 \us30/U10  ( .A0(\us30/n313 ), .A1(\us30/n5 ), .B0(\us30/n23 ), 
        .B1(\us30/n2 ), .C0(\us30/n328 ), .Y(\us30/n320 ) );
  AOI221X1 \us30/U9  ( .A0(\us30/n40 ), .A1(\us30/n136 ), .B0(\us30/n33 ), 
        .B1(\us30/n178 ), .C0(\us30/n338 ), .Y(\us30/n337 ) );
  AOI222XL \us30/U8  ( .A0(\us30/n278 ), .A1(\us30/n24 ), .B0(\us30/n42 ), 
        .B1(\us30/n33 ), .C0(\us30/n43 ), .C1(\us30/n136 ), .Y(\us30/n351 ) );
  AOI31X1 \us30/U7  ( .A0(sa30[2]), .A1(\us30/n58 ), .A2(sa30[1]), .B0(
        \us30/n40 ), .Y(\us30/n350 ) );
  AOI31X1 \us30/U6  ( .A0(\us30/n44 ), .A1(\us30/n129 ), .A2(\us30/n130 ), 
        .B0(\us30/n131 ), .Y(\us30/n128 ) );
  AOI221X1 \us30/U5  ( .A0(\us30/n40 ), .A1(\us30/n136 ), .B0(\us30/n33 ), 
        .B1(\us30/n47 ), .C0(\us30/n156 ), .Y(\us30/n141 ) );
  OAI32X1 \us30/U4  ( .A0(\us30/n18 ), .A1(sa30[1]), .A2(\us30/n159 ), .B0(
        sa30[4]), .B1(\us30/n182 ), .Y(\us30/n318 ) );
  OAI32X1 \us30/U3  ( .A0(\us30/n210 ), .A1(\us30/n145 ), .A2(\us30/n18 ), 
        .B0(\us30/n27 ), .B1(\us30/n211 ), .Y(\us30/n209 ) );
  AOI221X1 \us30/U2  ( .A0(\us30/n278 ), .A1(\us30/n40 ), .B0(\us30/n185 ), 
        .B1(\us30/n2 ), .C0(\us30/n279 ), .Y(\us30/n273 ) );
  AOI31XL \us30/U1  ( .A0(\us30/n79 ), .A1(\us30/n44 ), .A2(\us30/n2 ), .B0(
        \us30/n280 ), .Y(\us30/n339 ) );
  NAND2X1 \us31/U366  ( .A(\us31/n47 ), .B(\us31/n226 ), .Y(\us31/n189 ) );
  NOR2X1 \us31/U365  ( .A(\us31/n226 ), .B(sa31[3]), .Y(\us31/n242 ) );
  INVX1 \us31/U364  ( .A(\us31/n242 ), .Y(\us31/n205 ) );
  AND2X1 \us31/U363  ( .A(\us31/n189 ), .B(\us31/n205 ), .Y(\us31/n65 ) );
  NOR2X1 \us31/U362  ( .A(\us31/n226 ), .B(\us31/n47 ), .Y(\us31/n45 ) );
  NOR2X1 \us31/U361  ( .A(\us31/n259 ), .B(\us31/n45 ), .Y(\us31/n73 ) );
  NAND2BX1 \us31/U360  ( .AN(\us31/n73 ), .B(\us31/n6 ), .Y(\us31/n158 ) );
  NOR2X1 \us31/U359  ( .A(\us31/n226 ), .B(\us31/n159 ), .Y(\us31/n95 ) );
  INVX1 \us31/U358  ( .A(\us31/n95 ), .Y(\us31/n111 ) );
  NOR2X1 \us31/U357  ( .A(\us31/n145 ), .B(sa31[1]), .Y(\us31/n42 ) );
  INVX1 \us31/U356  ( .A(\us31/n42 ), .Y(\us31/n121 ) );
  INVX1 \us31/U355  ( .A(\us31/n47 ), .Y(\us31/n96 ) );
  OAI211X1 \us31/U354  ( .A0(\us31/n65 ), .A1(\us31/n27 ), .B0(\us31/n158 ), 
        .C0(\us31/n358 ), .Y(\us31/n355 ) );
  NOR2X1 \us31/U353  ( .A(\us31/n226 ), .B(\us31/n145 ), .Y(\us31/n59 ) );
  NOR2X1 \us31/U352  ( .A(\us31/n96 ), .B(\us31/n59 ), .Y(\us31/n271 ) );
  NOR2X1 \us31/U351  ( .A(\us31/n226 ), .B(\us31/n278 ), .Y(\us31/n217 ) );
  INVX1 \us31/U350  ( .A(\us31/n217 ), .Y(\us31/n150 ) );
  NAND2X1 \us31/U349  ( .A(\us31/n44 ), .B(\us31/n150 ), .Y(\us31/n147 ) );
  NAND2X1 \us31/U348  ( .A(sa31[4]), .B(\us31/n226 ), .Y(\us31/n101 ) );
  INVX1 \us31/U347  ( .A(\us31/n159 ), .Y(\us31/n188 ) );
  NOR2X1 \us31/U346  ( .A(\us31/n188 ), .B(\us31/n226 ), .Y(\us31/n25 ) );
  INVX1 \us31/U345  ( .A(\us31/n172 ), .Y(\us31/n107 ) );
  AOI22X1 \us31/U344  ( .A0(\us31/n33 ), .A1(\us31/n147 ), .B0(\us31/n24 ), 
        .B1(\us31/n107 ), .Y(\us31/n357 ) );
  OAI221XL \us31/U343  ( .A0(\us31/n18 ), .A1(\us31/n121 ), .B0(\us31/n271 ), 
        .B1(\us31/n20 ), .C0(\us31/n357 ), .Y(\us31/n356 ) );
  MXI2X1 \us31/U342  ( .A(\us31/n355 ), .B(\us31/n356 ), .S0(\us31/n252 ), .Y(
        \us31/n331 ) );
  INVX1 \us31/U341  ( .A(\us31/n59 ), .Y(\us31/n79 ) );
  AND2X1 \us31/U340  ( .A(\us31/n101 ), .B(\us31/n79 ), .Y(\us31/n325 ) );
  XNOR2X1 \us31/U339  ( .A(sa31[5]), .B(\us31/n226 ), .Y(\us31/n352 ) );
  NOR2X1 \us31/U338  ( .A(\us31/n226 ), .B(\us31/n136 ), .Y(\us31/n281 ) );
  INVX1 \us31/U337  ( .A(\us31/n281 ), .Y(\us31/n19 ) );
  NAND2X1 \us31/U336  ( .A(\us31/n145 ), .B(\us31/n226 ), .Y(\us31/n223 ) );
  AOI21X1 \us31/U335  ( .A0(\us31/n19 ), .A1(\us31/n223 ), .B0(\us31/n27 ), 
        .Y(\us31/n354 ) );
  AOI31X1 \us31/U334  ( .A0(\us31/n6 ), .A1(\us31/n352 ), .A2(\us31/n259 ), 
        .B0(\us31/n354 ), .Y(\us31/n353 ) );
  OAI221XL \us31/U333  ( .A0(\us31/n20 ), .A1(\us31/n34 ), .B0(\us31/n325 ), 
        .B1(\us31/n4 ), .C0(\us31/n353 ), .Y(\us31/n347 ) );
  INVX1 \us31/U332  ( .A(\us31/n352 ), .Y(\us31/n349 ) );
  NAND2X1 \us31/U331  ( .A(\us31/n278 ), .B(\us31/n6 ), .Y(\us31/n74 ) );
  OAI211X1 \us31/U330  ( .A0(\us31/n349 ), .A1(\us31/n74 ), .B0(\us31/n350 ), 
        .C0(\us31/n351 ), .Y(\us31/n348 ) );
  MXI2X1 \us31/U329  ( .A(\us31/n347 ), .B(\us31/n348 ), .S0(\us31/n252 ), .Y(
        \us31/n332 ) );
  NOR2X1 \us31/U328  ( .A(\us31/n44 ), .B(\us31/n226 ), .Y(\us31/n157 ) );
  INVX1 \us31/U327  ( .A(\us31/n157 ), .Y(\us31/n240 ) );
  NAND2X1 \us31/U326  ( .A(\us31/n240 ), .B(\us31/n189 ), .Y(\us31/n68 ) );
  NOR2X1 \us31/U325  ( .A(\us31/n20 ), .B(\us31/n159 ), .Y(\us31/n225 ) );
  NOR2X1 \us31/U324  ( .A(\us31/n225 ), .B(\us31/n40 ), .Y(\us31/n345 ) );
  INVX1 \us31/U323  ( .A(\us31/n278 ), .Y(\us31/n94 ) );
  NAND2X1 \us31/U322  ( .A(\us31/n94 ), .B(\us31/n226 ), .Y(\us31/n199 ) );
  NAND2X1 \us31/U321  ( .A(\us31/n199 ), .B(\us31/n205 ), .Y(\us31/n82 ) );
  NAND2X1 \us31/U320  ( .A(\us31/n19 ), .B(\us31/n199 ), .Y(\us31/n295 ) );
  NOR2X1 \us31/U319  ( .A(\us31/n226 ), .B(\us31/n259 ), .Y(\us31/n210 ) );
  NOR2X1 \us31/U318  ( .A(\us31/n27 ), .B(\us31/n210 ), .Y(\us31/n173 ) );
  MXI2X1 \us31/U317  ( .A(\us31/n345 ), .B(\us31/n346 ), .S0(\us31/n252 ), .Y(
        \us31/n342 ) );
  NOR2X1 \us31/U316  ( .A(sa31[1]), .B(sa31[3]), .Y(\us31/n163 ) );
  INVX1 \us31/U315  ( .A(\us31/n163 ), .Y(\us31/n37 ) );
  INVX1 \us31/U314  ( .A(\us31/n173 ), .Y(\us31/n344 ) );
  AOI21X1 \us31/U313  ( .A0(\us31/n240 ), .A1(\us31/n37 ), .B0(\us31/n344 ), 
        .Y(\us31/n343 ) );
  AOI211X1 \us31/U312  ( .A0(\us31/n5 ), .A1(\us31/n68 ), .B0(\us31/n342 ), 
        .C0(\us31/n343 ), .Y(\us31/n333 ) );
  NOR2X1 \us31/U311  ( .A(\us31/n18 ), .B(\us31/n226 ), .Y(\us31/n258 ) );
  NAND2X1 \us31/U310  ( .A(\us31/n278 ), .B(sa31[1]), .Y(\us31/n204 ) );
  NOR2X1 \us31/U309  ( .A(\us31/n188 ), .B(sa31[1]), .Y(\us31/n179 ) );
  INVX1 \us31/U308  ( .A(\us31/n179 ), .Y(\us31/n330 ) );
  NAND2X1 \us31/U307  ( .A(\us31/n204 ), .B(\us31/n330 ), .Y(\us31/n239 ) );
  NOR2X1 \us31/U306  ( .A(\us31/n136 ), .B(sa31[1]), .Y(\us31/n299 ) );
  NOR2X1 \us31/U305  ( .A(\us31/n299 ), .B(\us31/n210 ), .Y(\us31/n341 ) );
  OAI32X1 \us31/U304  ( .A0(\us31/n27 ), .A1(\us31/n278 ), .A2(\us31/n95 ), 
        .B0(\us31/n341 ), .B1(\us31/n4 ), .Y(\us31/n340 ) );
  INVX1 \us31/U303  ( .A(\us31/n45 ), .Y(\us31/n126 ) );
  NAND2X1 \us31/U302  ( .A(\us31/n126 ), .B(\us31/n101 ), .Y(\us31/n178 ) );
  NOR2X1 \us31/U301  ( .A(\us31/n18 ), .B(\us31/n136 ), .Y(\us31/n280 ) );
  OAI21XL \us31/U300  ( .A0(\us31/n4 ), .A1(\us31/n121 ), .B0(\us31/n339 ), 
        .Y(\us31/n338 ) );
  MXI2X1 \us31/U299  ( .A(\us31/n336 ), .B(\us31/n337 ), .S0(\us31/n252 ), .Y(
        \us31/n335 ) );
  NOR2X1 \us31/U298  ( .A(\us31/n258 ), .B(\us31/n335 ), .Y(\us31/n334 ) );
  MX4X1 \us31/U297  ( .A(\us31/n331 ), .B(\us31/n332 ), .C(\us31/n333 ), .D(
        \us31/n334 ), .S0(sa31[6]), .S1(\us31/n234 ), .Y(sa32_sr[0]) );
  INVX1 \us31/U296  ( .A(\us31/n299 ), .Y(\us31/n80 ) );
  NOR2X1 \us31/U295  ( .A(\us31/n111 ), .B(\us31/n18 ), .Y(\us31/n269 ) );
  INVX1 \us31/U294  ( .A(\us31/n269 ), .Y(\us31/n75 ) );
  OAI221XL \us31/U293  ( .A0(\us31/n18 ), .A1(\us31/n330 ), .B0(\us31/n20 ), 
        .B1(\us31/n80 ), .C0(\us31/n75 ), .Y(\us31/n329 ) );
  AOI221X1 \us31/U292  ( .A0(\us31/n325 ), .A1(\us31/n33 ), .B0(\us31/n24 ), 
        .B1(\us31/n303 ), .C0(\us31/n329 ), .Y(\us31/n319 ) );
  NOR2X1 \us31/U291  ( .A(\us31/n234 ), .B(sa31[5]), .Y(\us31/n14 ) );
  NOR2X1 \us31/U290  ( .A(\us31/n25 ), .B(\us31/n299 ), .Y(\us31/n313 ) );
  NAND2X1 \us31/U289  ( .A(\us31/n44 ), .B(\us31/n226 ), .Y(\us31/n300 ) );
  AND2X1 \us31/U288  ( .A(\us31/n300 ), .B(\us31/n240 ), .Y(\us31/n23 ) );
  OAI32X1 \us31/U287  ( .A0(\us31/n4 ), .A1(\us31/n145 ), .A2(\us31/n210 ), 
        .B0(\us31/n137 ), .B1(\us31/n27 ), .Y(\us31/n328 ) );
  NOR2X1 \us31/U286  ( .A(sa31[0]), .B(sa31[5]), .Y(\us31/n16 ) );
  INVX1 \us31/U285  ( .A(\us31/n16 ), .Y(\us31/n114 ) );
  INVX1 \us31/U284  ( .A(\us31/n145 ), .Y(\us31/n149 ) );
  NOR2X1 \us31/U283  ( .A(\us31/n47 ), .B(sa31[1]), .Y(\us31/n98 ) );
  INVX1 \us31/U282  ( .A(\us31/n98 ), .Y(\us31/n284 ) );
  OAI21XL \us31/U281  ( .A0(\us31/n69 ), .A1(\us31/n284 ), .B0(\us31/n27 ), 
        .Y(\us31/n327 ) );
  AOI31X1 \us31/U280  ( .A0(\us31/n111 ), .A1(\us31/n149 ), .A2(\us31/n327 ), 
        .B0(\us31/n225 ), .Y(\us31/n326 ) );
  OAI21XL \us31/U279  ( .A0(\us31/n325 ), .A1(\us31/n18 ), .B0(\us31/n326 ), 
        .Y(\us31/n322 ) );
  NAND2X1 \us31/U278  ( .A(\us31/n19 ), .B(\us31/n189 ), .Y(\us31/n71 ) );
  NOR2X1 \us31/U277  ( .A(\us31/n71 ), .B(\us31/n18 ), .Y(\us31/n135 ) );
  AOI21X1 \us31/U276  ( .A0(\us31/n40 ), .A1(sa31[4]), .B0(\us31/n135 ), .Y(
        \us31/n324 ) );
  OAI221XL \us31/U275  ( .A0(\us31/n47 ), .A1(\us31/n27 ), .B0(\us31/n65 ), 
        .B1(\us31/n20 ), .C0(\us31/n324 ), .Y(\us31/n323 ) );
  AOI22X1 \us31/U274  ( .A0(\us31/n55 ), .A1(\us31/n322 ), .B0(\us31/n89 ), 
        .B1(\us31/n323 ), .Y(\us31/n321 ) );
  OAI221XL \us31/U273  ( .A0(\us31/n319 ), .A1(\us31/n52 ), .B0(\us31/n320 ), 
        .B1(\us31/n114 ), .C0(\us31/n321 ), .Y(\us31/n304 ) );
  NOR2X1 \us31/U272  ( .A(\us31/n226 ), .B(\us31/n58 ), .Y(\us31/n290 ) );
  INVX1 \us31/U271  ( .A(\us31/n290 ), .Y(\us31/n200 ) );
  NAND2X1 \us31/U270  ( .A(\us31/n34 ), .B(\us31/n200 ), .Y(\us31/n120 ) );
  INVX1 \us31/U269  ( .A(\us31/n210 ), .Y(\us31/n100 ) );
  OAI221XL \us31/U268  ( .A0(\us31/n20 ), .A1(\us31/n100 ), .B0(sa31[3]), .B1(
        \us31/n4 ), .C0(\us31/n262 ), .Y(\us31/n317 ) );
  INVX1 \us31/U267  ( .A(\us31/n258 ), .Y(\us31/n182 ) );
  AOI211X1 \us31/U266  ( .A0(\us31/n33 ), .A1(\us31/n120 ), .B0(\us31/n317 ), 
        .C0(\us31/n318 ), .Y(\us31/n306 ) );
  NAND2X1 \us31/U265  ( .A(\us31/n100 ), .B(\us31/n199 ), .Y(\us31/n151 ) );
  INVX1 \us31/U264  ( .A(\us31/n151 ), .Y(\us31/n314 ) );
  NOR2X1 \us31/U263  ( .A(\us31/n45 ), .B(\us31/n163 ), .Y(\us31/n160 ) );
  INVX1 \us31/U262  ( .A(\us31/n295 ), .Y(\us31/n92 ) );
  AOI21X1 \us31/U261  ( .A0(sa31[1]), .A1(\us31/n58 ), .B0(\us31/n98 ), .Y(
        \us31/n316 ) );
  OAI22X1 \us31/U260  ( .A0(\us31/n92 ), .A1(\us31/n18 ), .B0(\us31/n316 ), 
        .B1(\us31/n27 ), .Y(\us31/n315 ) );
  NOR2X1 \us31/U259  ( .A(\us31/n149 ), .B(\us31/n226 ), .Y(\us31/n41 ) );
  INVX1 \us31/U258  ( .A(\us31/n41 ), .Y(\us31/n105 ) );
  NAND2X1 \us31/U257  ( .A(\us31/n284 ), .B(\us31/n105 ), .Y(\us31/n227 ) );
  AOI21X1 \us31/U256  ( .A0(\us31/n313 ), .A1(\us31/n33 ), .B0(\us31/n269 ), 
        .Y(\us31/n312 ) );
  OAI221XL \us31/U255  ( .A0(\us31/n149 ), .A1(\us31/n20 ), .B0(\us31/n4 ), 
        .B1(\us31/n227 ), .C0(\us31/n312 ), .Y(\us31/n309 ) );
  AOI21X1 \us31/U254  ( .A0(\us31/n226 ), .A1(\us31/n188 ), .B0(\us31/n242 ), 
        .Y(\us31/n185 ) );
  INVX1 \us31/U253  ( .A(\us31/n185 ), .Y(\us31/n48 ) );
  AND2X1 \us31/U252  ( .A(\us31/n223 ), .B(\us31/n240 ), .Y(\us31/n28 ) );
  OAI221XL \us31/U251  ( .A0(\us31/n27 ), .A1(\us31/n44 ), .B0(\us31/n4 ), 
        .B1(\us31/n48 ), .C0(\us31/n311 ), .Y(\us31/n310 ) );
  AOI22X1 \us31/U250  ( .A0(\us31/n89 ), .A1(\us31/n309 ), .B0(\us31/n55 ), 
        .B1(\us31/n310 ), .Y(\us31/n308 ) );
  OAI221XL \us31/U249  ( .A0(\us31/n306 ), .A1(\us31/n52 ), .B0(\us31/n307 ), 
        .B1(\us31/n114 ), .C0(\us31/n308 ), .Y(\us31/n305 ) );
  MX2X1 \us31/U248  ( .A(\us31/n304 ), .B(\us31/n305 ), .S0(sa31[6]), .Y(
        sa32_sr[1]) );
  INVX1 \us31/U247  ( .A(\us31/n187 ), .Y(\us31/n61 ) );
  MXI2X1 \us31/U246  ( .A(\us31/n303 ), .B(\us31/n61 ), .S0(\us31/n69 ), .Y(
        \us31/n301 ) );
  MXI2X1 \us31/U245  ( .A(\us31/n301 ), .B(\us31/n147 ), .S0(\us31/n302 ), .Y(
        \us31/n285 ) );
  NAND2X1 \us31/U244  ( .A(\us31/n200 ), .B(\us31/n300 ), .Y(\us31/n99 ) );
  INVX1 \us31/U243  ( .A(\us31/n99 ), .Y(\us31/n296 ) );
  NOR2X1 \us31/U242  ( .A(\us31/n299 ), .B(\us31/n242 ), .Y(\us31/n298 ) );
  NAND2X1 \us31/U241  ( .A(sa31[1]), .B(\us31/n47 ), .Y(\us31/n122 ) );
  NOR2X1 \us31/U240  ( .A(\us31/n159 ), .B(\us31/n217 ), .Y(\us31/n198 ) );
  OAI221XL \us31/U239  ( .A0(\us31/n298 ), .A1(\us31/n27 ), .B0(\us31/n20 ), 
        .B1(\us31/n122 ), .C0(\us31/n132 ), .Y(\us31/n297 ) );
  AOI221X1 \us31/U238  ( .A0(\us31/n225 ), .A1(\us31/n226 ), .B0(\us31/n296 ), 
        .B1(\us31/n6 ), .C0(\us31/n297 ), .Y(\us31/n291 ) );
  OAI2BB2X1 \us31/U237  ( .B0(\us31/n27 ), .B1(\us31/n295 ), .A0N(\us31/n34 ), 
        .A1N(\us31/n24 ), .Y(\us31/n293 ) );
  AOI21X1 \us31/U236  ( .A0(\us31/n101 ), .A1(\us31/n150 ), .B0(\us31/n20 ), 
        .Y(\us31/n294 ) );
  AOI211X1 \us31/U235  ( .A0(\us31/n5 ), .A1(\us31/n79 ), .B0(\us31/n293 ), 
        .C0(\us31/n294 ), .Y(\us31/n292 ) );
  INVX1 \us31/U234  ( .A(\us31/n89 ), .Y(\us31/n10 ) );
  OAI22X1 \us31/U233  ( .A0(\us31/n291 ), .A1(\us31/n114 ), .B0(\us31/n292 ), 
        .B1(\us31/n10 ), .Y(\us31/n286 ) );
  INVX1 \us31/U232  ( .A(\us31/n225 ), .Y(\us31/n288 ) );
  NAND2X1 \us31/U231  ( .A(\us31/n200 ), .B(\us31/n284 ), .Y(\us31/n102 ) );
  NOR2X1 \us31/U230  ( .A(\us31/n290 ), .B(\us31/n163 ), .Y(\us31/n184 ) );
  AOI22X1 \us31/U229  ( .A0(\us31/n102 ), .A1(\us31/n69 ), .B0(\us31/n184 ), 
        .B1(\us31/n33 ), .Y(\us31/n289 ) );
  AOI31X1 \us31/U228  ( .A0(\us31/n132 ), .A1(\us31/n288 ), .A2(\us31/n289 ), 
        .B0(\us31/n52 ), .Y(\us31/n287 ) );
  AOI211X1 \us31/U227  ( .A0(\us31/n285 ), .A1(\us31/n55 ), .B0(\us31/n286 ), 
        .C0(\us31/n287 ), .Y(\us31/n263 ) );
  NAND2X1 \us31/U226  ( .A(\us31/n284 ), .B(\us31/n122 ), .Y(\us31/n125 ) );
  NOR2X1 \us31/U225  ( .A(\us31/n199 ), .B(\us31/n4 ), .Y(\us31/n50 ) );
  AOI21X1 \us31/U224  ( .A0(\us31/n200 ), .A1(\us31/n223 ), .B0(\us31/n20 ), 
        .Y(\us31/n283 ) );
  AOI211X1 \us31/U223  ( .A0(\us31/n5 ), .A1(\us31/n125 ), .B0(\us31/n50 ), 
        .C0(\us31/n283 ), .Y(\us31/n282 ) );
  OAI221XL \us31/U222  ( .A0(\us31/n281 ), .A1(\us31/n27 ), .B0(\us31/n4 ), 
        .B1(\us31/n111 ), .C0(\us31/n282 ), .Y(\us31/n265 ) );
  INVX1 \us31/U221  ( .A(\us31/n280 ), .Y(\us31/n247 ) );
  NAND2X1 \us31/U220  ( .A(\us31/n41 ), .B(\us31/n33 ), .Y(\us31/n272 ) );
  OAI221XL \us31/U219  ( .A0(sa31[1]), .A1(\us31/n247 ), .B0(\us31/n4 ), .B1(
        \us31/n189 ), .C0(\us31/n272 ), .Y(\us31/n279 ) );
  NAND2X1 \us31/U218  ( .A(sa31[2]), .B(\us31/n149 ), .Y(\us31/n276 ) );
  XNOR2X1 \us31/U217  ( .A(\us31/n129 ), .B(sa31[1]), .Y(\us31/n155 ) );
  MXI2X1 \us31/U216  ( .A(\us31/n276 ), .B(\us31/n277 ), .S0(\us31/n155 ), .Y(
        \us31/n275 ) );
  OAI22X1 \us31/U215  ( .A0(\us31/n273 ), .A1(\us31/n10 ), .B0(\us31/n274 ), 
        .B1(\us31/n52 ), .Y(\us31/n266 ) );
  NOR2X1 \us31/U214  ( .A(\us31/n20 ), .B(\us31/n226 ), .Y(\us31/n176 ) );
  OAI21XL \us31/U213  ( .A0(\us31/n4 ), .A1(\us31/n271 ), .B0(\us31/n272 ), 
        .Y(\us31/n270 ) );
  OAI31X1 \us31/U212  ( .A0(\us31/n176 ), .A1(\us31/n269 ), .A2(\us31/n270 ), 
        .B0(\us31/n16 ), .Y(\us31/n268 ) );
  INVX1 \us31/U211  ( .A(\us31/n268 ), .Y(\us31/n267 ) );
  AOI211X1 \us31/U210  ( .A0(\us31/n55 ), .A1(\us31/n265 ), .B0(\us31/n266 ), 
        .C0(\us31/n267 ), .Y(\us31/n264 ) );
  MXI2X1 \us31/U209  ( .A(\us31/n263 ), .B(\us31/n264 ), .S0(sa31[6]), .Y(
        sa32_sr[2]) );
  NOR2X1 \us31/U208  ( .A(\us31/n94 ), .B(sa31[1]), .Y(\us31/n211 ) );
  INVX1 \us31/U207  ( .A(\us31/n262 ), .Y(\us31/n261 ) );
  AOI211X1 \us31/U206  ( .A0(\us31/n259 ), .A1(\us31/n24 ), .B0(\us31/n260 ), 
        .C0(\us31/n261 ), .Y(\us31/n255 ) );
  OAI22X1 \us31/U205  ( .A0(\us31/n20 ), .A1(\us31/n68 ), .B0(\us31/n27 ), 
        .B1(\us31/n37 ), .Y(\us31/n257 ) );
  NOR3X1 \us31/U204  ( .A(\us31/n257 ), .B(\us31/n258 ), .C(\us31/n50 ), .Y(
        \us31/n256 ) );
  MXI2X1 \us31/U203  ( .A(\us31/n255 ), .B(\us31/n256 ), .S0(\us31/n252 ), .Y(
        \us31/n254 ) );
  AOI221X1 \us31/U202  ( .A0(\us31/n211 ), .A1(\us31/n5 ), .B0(\us31/n40 ), 
        .B1(sa31[4]), .C0(\us31/n254 ), .Y(\us31/n248 ) );
  INVX1 \us31/U201  ( .A(\us31/n211 ), .Y(\us31/n106 ) );
  NAND2X1 \us31/U200  ( .A(\us31/n200 ), .B(\us31/n106 ), .Y(\us31/n83 ) );
  NAND2X1 \us31/U199  ( .A(\us31/n199 ), .B(\us31/n204 ), .Y(\us31/n169 ) );
  AOI2BB2X1 \us31/U198  ( .B0(\us31/n65 ), .B1(\us31/n24 ), .A0N(\us31/n169 ), 
        .A1N(\us31/n20 ), .Y(\us31/n253 ) );
  OAI221XL \us31/U197  ( .A0(\us31/n172 ), .A1(\us31/n18 ), .B0(\us31/n27 ), 
        .B1(\us31/n83 ), .C0(\us31/n253 ), .Y(\us31/n251 ) );
  MXI2X1 \us31/U196  ( .A(\us31/n250 ), .B(\us31/n251 ), .S0(\us31/n252 ), .Y(
        \us31/n249 ) );
  MXI2X1 \us31/U195  ( .A(\us31/n248 ), .B(\us31/n249 ), .S0(\us31/n234 ), .Y(
        \us31/n228 ) );
  OAI21XL \us31/U194  ( .A0(\us31/n58 ), .A1(\us31/n27 ), .B0(\us31/n247 ), 
        .Y(\us31/n245 ) );
  NOR2X1 \us31/U193  ( .A(sa31[7]), .B(\us31/n145 ), .Y(\us31/n246 ) );
  XNOR2X1 \us31/U192  ( .A(\us31/n69 ), .B(sa31[1]), .Y(\us31/n130 ) );
  MXI2X1 \us31/U191  ( .A(\us31/n245 ), .B(\us31/n246 ), .S0(\us31/n130 ), .Y(
        \us31/n243 ) );
  OAI211X1 \us31/U190  ( .A0(\us31/n4 ), .A1(\us31/n149 ), .B0(\us31/n243 ), 
        .C0(\us31/n244 ), .Y(\us31/n230 ) );
  NOR2X1 \us31/U189  ( .A(\us31/n242 ), .B(\us31/n137 ), .Y(\us31/n70 ) );
  OAI221XL \us31/U188  ( .A0(\us31/n159 ), .A1(\us31/n27 ), .B0(\us31/n20 ), 
        .B1(\us31/n34 ), .C0(\us31/n241 ), .Y(\us31/n231 ) );
  NAND2X1 \us31/U187  ( .A(\us31/n101 ), .B(\us31/n240 ), .Y(\us31/n76 ) );
  AOI21X1 \us31/U186  ( .A0(\us31/n122 ), .A1(\us31/n106 ), .B0(\us31/n129 ), 
        .Y(\us31/n237 ) );
  INVX1 \us31/U185  ( .A(\us31/n239 ), .Y(\us31/n238 ) );
  OAI21XL \us31/U184  ( .A0(\us31/n237 ), .A1(\us31/n43 ), .B0(\us31/n238 ), 
        .Y(\us31/n236 ) );
  OAI221XL \us31/U183  ( .A0(\us31/n18 ), .A1(\us31/n76 ), .B0(\us31/n59 ), 
        .B1(\us31/n27 ), .C0(\us31/n236 ), .Y(\us31/n232 ) );
  AOI2BB2X1 \us31/U182  ( .B0(\us31/n24 ), .B1(\us31/n187 ), .A0N(\us31/n227 ), 
        .A1N(\us31/n20 ), .Y(\us31/n235 ) );
  OAI211X1 \us31/U181  ( .A0(\us31/n27 ), .A1(\us31/n122 ), .B0(\us31/n158 ), 
        .C0(\us31/n235 ), .Y(\us31/n233 ) );
  MX4X1 \us31/U180  ( .A(\us31/n230 ), .B(\us31/n231 ), .C(\us31/n232 ), .D(
        \us31/n233 ), .S0(\us31/n234 ), .S1(sa31[5]), .Y(\us31/n229 ) );
  MX2X1 \us31/U179  ( .A(\us31/n228 ), .B(\us31/n229 ), .S0(sa31[6]), .Y(
        sa32_sr[3]) );
  NOR2BX1 \us31/U178  ( .AN(\us31/n204 ), .B(\us31/n137 ), .Y(\us31/n110 ) );
  INVX1 \us31/U177  ( .A(\us31/n110 ), .Y(\us31/n64 ) );
  AOI22X1 \us31/U176  ( .A0(\us31/n225 ), .A1(\us31/n226 ), .B0(\us31/n6 ), 
        .B1(\us31/n227 ), .Y(\us31/n224 ) );
  OAI221XL \us31/U175  ( .A0(\us31/n27 ), .A1(\us31/n64 ), .B0(\us31/n4 ), 
        .B1(\us31/n83 ), .C0(\us31/n224 ), .Y(\us31/n212 ) );
  NAND2X1 \us31/U174  ( .A(\us31/n34 ), .B(\us31/n204 ), .Y(\us31/n221 ) );
  OAI21XL \us31/U173  ( .A0(\us31/n69 ), .A1(\us31/n223 ), .B0(\us31/n27 ), 
        .Y(\us31/n222 ) );
  NOR2X1 \us31/U172  ( .A(\us31/n217 ), .B(\us31/n42 ), .Y(\us31/n208 ) );
  AOI211X1 \us31/U171  ( .A0(\us31/n208 ), .A1(\us31/n5 ), .B0(\us31/n220 ), 
        .C0(\us31/n173 ), .Y(\us31/n219 ) );
  OAI22X1 \us31/U170  ( .A0(\us31/n218 ), .A1(\us31/n10 ), .B0(\us31/n219 ), 
        .B1(\us31/n114 ), .Y(\us31/n213 ) );
  INVX1 \us31/U169  ( .A(\us31/n135 ), .Y(\us31/n215 ) );
  NOR2X1 \us31/U168  ( .A(\us31/n4 ), .B(\us31/n159 ), .Y(\us31/n31 ) );
  INVX1 \us31/U167  ( .A(\us31/n31 ), .Y(\us31/n196 ) );
  AOI31X1 \us31/U166  ( .A0(\us31/n215 ), .A1(\us31/n196 ), .A2(\us31/n216 ), 
        .B0(\us31/n52 ), .Y(\us31/n214 ) );
  AOI211X1 \us31/U165  ( .A0(\us31/n55 ), .A1(\us31/n212 ), .B0(\us31/n213 ), 
        .C0(\us31/n214 ), .Y(\us31/n190 ) );
  INVX1 \us31/U164  ( .A(\us31/n207 ), .Y(\us31/n192 ) );
  NOR2X1 \us31/U163  ( .A(\us31/n25 ), .B(\us31/n98 ), .Y(\us31/n32 ) );
  OAI22X1 \us31/U162  ( .A0(\us31/n28 ), .A1(\us31/n4 ), .B0(\us31/n188 ), 
        .B1(\us31/n27 ), .Y(\us31/n206 ) );
  NAND2X1 \us31/U161  ( .A(\us31/n204 ), .B(\us31/n80 ), .Y(\us31/n118 ) );
  INVX1 \us31/U160  ( .A(\us31/n118 ), .Y(\us31/n123 ) );
  NAND2X1 \us31/U159  ( .A(\us31/n94 ), .B(\us31/n79 ), .Y(\us31/n203 ) );
  OAI2BB1X1 \us31/U158  ( .A0N(\us31/n199 ), .A1N(\us31/n200 ), .B0(\us31/n33 ), .Y(\us31/n195 ) );
  INVX1 \us31/U157  ( .A(\us31/n55 ), .Y(\us31/n12 ) );
  AOI31X1 \us31/U156  ( .A0(\us31/n195 ), .A1(\us31/n196 ), .A2(\us31/n197 ), 
        .B0(\us31/n12 ), .Y(\us31/n194 ) );
  AOI211X1 \us31/U155  ( .A0(\us31/n89 ), .A1(\us31/n192 ), .B0(\us31/n193 ), 
        .C0(\us31/n194 ), .Y(\us31/n191 ) );
  MXI2X1 \us31/U154  ( .A(\us31/n190 ), .B(\us31/n191 ), .S0(sa31[6]), .Y(
        sa32_sr[4]) );
  OAI21XL \us31/U153  ( .A0(\us31/n69 ), .A1(\us31/n189 ), .B0(\us31/n27 ), 
        .Y(\us31/n186 ) );
  INVX1 \us31/U152  ( .A(\us31/n183 ), .Y(\us31/n180 ) );
  NAND2X1 \us31/U151  ( .A(\us31/n74 ), .B(\us31/n182 ), .Y(\us31/n181 ) );
  AOI211X1 \us31/U150  ( .A0(\us31/n179 ), .A1(\us31/n24 ), .B0(\us31/n180 ), 
        .C0(\us31/n181 ), .Y(\us31/n165 ) );
  INVX1 \us31/U149  ( .A(\us31/n178 ), .Y(\us31/n175 ) );
  AOI211X1 \us31/U148  ( .A0(\us31/n175 ), .A1(\us31/n5 ), .B0(\us31/n176 ), 
        .C0(\us31/n177 ), .Y(\us31/n174 ) );
  OAI221XL \us31/U147  ( .A0(\us31/n159 ), .A1(\us31/n27 ), .B0(\us31/n145 ), 
        .B1(\us31/n20 ), .C0(\us31/n174 ), .Y(\us31/n167 ) );
  MXI2X1 \us31/U146  ( .A(\us31/n40 ), .B(\us31/n173 ), .S0(\us31/n96 ), .Y(
        \us31/n170 ) );
  AOI22X1 \us31/U145  ( .A0(\us31/n137 ), .A1(\us31/n24 ), .B0(\us31/n172 ), 
        .B1(\us31/n6 ), .Y(\us31/n171 ) );
  OAI211X1 \us31/U144  ( .A0(\us31/n20 ), .A1(\us31/n169 ), .B0(\us31/n170 ), 
        .C0(\us31/n171 ), .Y(\us31/n168 ) );
  AOI22X1 \us31/U143  ( .A0(\us31/n89 ), .A1(\us31/n167 ), .B0(\us31/n55 ), 
        .B1(\us31/n168 ), .Y(\us31/n166 ) );
  OAI221XL \us31/U142  ( .A0(\us31/n164 ), .A1(\us31/n114 ), .B0(\us31/n165 ), 
        .B1(\us31/n52 ), .C0(\us31/n166 ), .Y(\us31/n138 ) );
  OAI21XL \us31/U141  ( .A0(\us31/n41 ), .A1(\us31/n163 ), .B0(\us31/n69 ), 
        .Y(\us31/n162 ) );
  AOI221X1 \us31/U140  ( .A0(\us31/n159 ), .A1(\us31/n24 ), .B0(\us31/n160 ), 
        .B1(\us31/n33 ), .C0(\us31/n161 ), .Y(\us31/n140 ) );
  OAI21XL \us31/U139  ( .A0(\us31/n157 ), .A1(\us31/n20 ), .B0(\us31/n158 ), 
        .Y(\us31/n156 ) );
  NOR2X1 \us31/U138  ( .A(\us31/n4 ), .B(\us31/n136 ), .Y(\us31/n153 ) );
  NOR2X1 \us31/U137  ( .A(\us31/n145 ), .B(\us31/n69 ), .Y(\us31/n154 ) );
  MXI2X1 \us31/U136  ( .A(\us31/n153 ), .B(\us31/n154 ), .S0(\us31/n155 ), .Y(
        \us31/n152 ) );
  OAI221XL \us31/U135  ( .A0(\us31/n110 ), .A1(\us31/n18 ), .B0(\us31/n20 ), 
        .B1(\us31/n151 ), .C0(\us31/n152 ), .Y(\us31/n143 ) );
  AOI21X1 \us31/U134  ( .A0(\us31/n149 ), .A1(\us31/n150 ), .B0(\us31/n18 ), 
        .Y(\us31/n148 ) );
  AOI2BB1X1 \us31/U133  ( .A0N(\us31/n147 ), .A1N(\us31/n27 ), .B0(\us31/n148 ), .Y(\us31/n146 ) );
  OAI221XL \us31/U132  ( .A0(\us31/n145 ), .A1(\us31/n20 ), .B0(\us31/n4 ), 
        .B1(\us31/n34 ), .C0(\us31/n146 ), .Y(\us31/n144 ) );
  AOI22X1 \us31/U131  ( .A0(\us31/n89 ), .A1(\us31/n143 ), .B0(\us31/n14 ), 
        .B1(\us31/n144 ), .Y(\us31/n142 ) );
  OAI221XL \us31/U130  ( .A0(\us31/n140 ), .A1(\us31/n12 ), .B0(\us31/n141 ), 
        .B1(\us31/n114 ), .C0(\us31/n142 ), .Y(\us31/n139 ) );
  MX2X1 \us31/U129  ( .A(\us31/n138 ), .B(\us31/n139 ), .S0(sa31[6]), .Y(
        sa32_sr[5]) );
  INVX1 \us31/U128  ( .A(\us31/n70 ), .Y(\us31/n133 ) );
  OAI22X1 \us31/U127  ( .A0(\us31/n4 ), .A1(\us31/n136 ), .B0(\us31/n137 ), 
        .B1(\us31/n27 ), .Y(\us31/n134 ) );
  AOI211X1 \us31/U126  ( .A0(\us31/n133 ), .A1(\us31/n69 ), .B0(\us31/n134 ), 
        .C0(\us31/n135 ), .Y(\us31/n112 ) );
  INVX1 \us31/U125  ( .A(\us31/n132 ), .Y(\us31/n131 ) );
  OAI21XL \us31/U124  ( .A0(\us31/n18 ), .A1(\us31/n37 ), .B0(\us31/n128 ), 
        .Y(\us31/n127 ) );
  OAI221XL \us31/U123  ( .A0(\us31/n18 ), .A1(\us31/n105 ), .B0(\us31/n123 ), 
        .B1(\us31/n27 ), .C0(\us31/n124 ), .Y(\us31/n116 ) );
  NAND2X1 \us31/U122  ( .A(\us31/n121 ), .B(\us31/n122 ), .Y(\us31/n30 ) );
  OAI221XL \us31/U121  ( .A0(\us31/n18 ), .A1(\us31/n118 ), .B0(\us31/n27 ), 
        .B1(\us31/n30 ), .C0(\us31/n119 ), .Y(\us31/n117 ) );
  AOI22X1 \us31/U120  ( .A0(\us31/n89 ), .A1(\us31/n116 ), .B0(\us31/n55 ), 
        .B1(\us31/n117 ), .Y(\us31/n115 ) );
  OAI221XL \us31/U119  ( .A0(\us31/n112 ), .A1(\us31/n52 ), .B0(\us31/n113 ), 
        .B1(\us31/n114 ), .C0(\us31/n115 ), .Y(\us31/n84 ) );
  OAI22X1 \us31/U118  ( .A0(\us31/n110 ), .A1(\us31/n4 ), .B0(\us31/n20 ), 
        .B1(\us31/n21 ), .Y(\us31/n108 ) );
  AOI21X1 \us31/U117  ( .A0(sa31[1]), .A1(\us31/n58 ), .B0(\us31/n27 ), .Y(
        \us31/n109 ) );
  AOI211X1 \us31/U116  ( .A0(\us31/n5 ), .A1(\us31/n107 ), .B0(\us31/n108 ), 
        .C0(\us31/n109 ), .Y(\us31/n86 ) );
  OAI22X1 \us31/U115  ( .A0(\us31/n45 ), .A1(\us31/n4 ), .B0(sa31[4]), .B1(
        \us31/n18 ), .Y(\us31/n103 ) );
  AOI21X1 \us31/U114  ( .A0(\us31/n105 ), .A1(\us31/n106 ), .B0(\us31/n20 ), 
        .Y(\us31/n104 ) );
  AOI211X1 \us31/U113  ( .A0(\us31/n33 ), .A1(\us31/n102 ), .B0(\us31/n103 ), 
        .C0(\us31/n104 ), .Y(\us31/n87 ) );
  NAND2X1 \us31/U112  ( .A(\us31/n100 ), .B(\us31/n101 ), .Y(\us31/n62 ) );
  OAI221XL \us31/U111  ( .A0(\us31/n27 ), .A1(\us31/n62 ), .B0(\us31/n4 ), 
        .B1(\us31/n21 ), .C0(\us31/n97 ), .Y(\us31/n90 ) );
  NOR3X1 \us31/U110  ( .A(\us31/n4 ), .B(\us31/n95 ), .C(\us31/n96 ), .Y(
        \us31/n67 ) );
  AOI31X1 \us31/U109  ( .A0(\us31/n79 ), .A1(\us31/n94 ), .A2(\us31/n6 ), .B0(
        \us31/n67 ), .Y(\us31/n93 ) );
  OAI221XL \us31/U108  ( .A0(\us31/n73 ), .A1(\us31/n27 ), .B0(\us31/n92 ), 
        .B1(\us31/n20 ), .C0(\us31/n93 ), .Y(\us31/n91 ) );
  AOI22X1 \us31/U107  ( .A0(\us31/n89 ), .A1(\us31/n90 ), .B0(\us31/n16 ), 
        .B1(\us31/n91 ), .Y(\us31/n88 ) );
  OAI221XL \us31/U106  ( .A0(\us31/n86 ), .A1(\us31/n52 ), .B0(\us31/n87 ), 
        .B1(\us31/n12 ), .C0(\us31/n88 ), .Y(\us31/n85 ) );
  MX2X1 \us31/U105  ( .A(\us31/n84 ), .B(\us31/n85 ), .S0(sa31[6]), .Y(
        sa32_sr[6]) );
  INVX1 \us31/U104  ( .A(\us31/n81 ), .Y(\us31/n77 ) );
  AOI21X1 \us31/U103  ( .A0(\us31/n79 ), .A1(\us31/n80 ), .B0(\us31/n27 ), .Y(
        \us31/n78 ) );
  AOI211X1 \us31/U102  ( .A0(\us31/n5 ), .A1(\us31/n76 ), .B0(\us31/n77 ), 
        .C0(\us31/n78 ), .Y(\us31/n51 ) );
  OAI211X1 \us31/U101  ( .A0(\us31/n73 ), .A1(\us31/n27 ), .B0(\us31/n74 ), 
        .C0(\us31/n75 ), .Y(\us31/n72 ) );
  AOI21X1 \us31/U100  ( .A0(\us31/n68 ), .A1(\us31/n69 ), .B0(\us31/n6 ), .Y(
        \us31/n63 ) );
  INVX1 \us31/U99  ( .A(\us31/n67 ), .Y(\us31/n66 ) );
  OAI221XL \us31/U98  ( .A0(\us31/n63 ), .A1(\us31/n64 ), .B0(\us31/n65 ), 
        .B1(\us31/n27 ), .C0(\us31/n66 ), .Y(\us31/n56 ) );
  AOI2BB2X1 \us31/U97  ( .B0(\us31/n61 ), .B1(\us31/n24 ), .A0N(\us31/n62 ), 
        .A1N(\us31/n20 ), .Y(\us31/n60 ) );
  OAI221XL \us31/U96  ( .A0(\us31/n58 ), .A1(\us31/n18 ), .B0(\us31/n59 ), 
        .B1(\us31/n27 ), .C0(\us31/n60 ), .Y(\us31/n57 ) );
  AOI22X1 \us31/U95  ( .A0(\us31/n55 ), .A1(\us31/n56 ), .B0(\us31/n16 ), .B1(
        \us31/n57 ), .Y(\us31/n54 ) );
  OAI221XL \us31/U94  ( .A0(\us31/n51 ), .A1(\us31/n52 ), .B0(\us31/n53 ), 
        .B1(\us31/n10 ), .C0(\us31/n54 ), .Y(\us31/n7 ) );
  INVX1 \us31/U93  ( .A(\us31/n50 ), .Y(\us31/n49 ) );
  OAI221XL \us31/U92  ( .A0(\us31/n47 ), .A1(\us31/n18 ), .B0(\us31/n27 ), 
        .B1(\us31/n48 ), .C0(\us31/n49 ), .Y(\us31/n46 ) );
  NOR2X1 \us31/U91  ( .A(\us31/n41 ), .B(\us31/n42 ), .Y(\us31/n38 ) );
  INVX1 \us31/U90  ( .A(\us31/n40 ), .Y(\us31/n39 ) );
  INVX1 \us31/U89  ( .A(\us31/n32 ), .Y(\us31/n26 ) );
  AOI21X1 \us31/U88  ( .A0(\us31/n5 ), .A1(\us31/n30 ), .B0(\us31/n31 ), .Y(
        \us31/n29 ) );
  OAI221XL \us31/U87  ( .A0(\us31/n26 ), .A1(\us31/n27 ), .B0(\us31/n28 ), 
        .B1(\us31/n20 ), .C0(\us31/n29 ), .Y(\us31/n15 ) );
  OAI221XL \us31/U86  ( .A0(\us31/n18 ), .A1(\us31/n19 ), .B0(\us31/n20 ), 
        .B1(\us31/n21 ), .C0(\us31/n22 ), .Y(\us31/n17 ) );
  AOI22X1 \us31/U85  ( .A0(\us31/n14 ), .A1(\us31/n15 ), .B0(\us31/n16 ), .B1(
        \us31/n17 ), .Y(\us31/n13 ) );
  OAI221XL \us31/U84  ( .A0(\us31/n9 ), .A1(\us31/n10 ), .B0(\us31/n11 ), .B1(
        \us31/n12 ), .C0(\us31/n13 ), .Y(\us31/n8 ) );
  MX2X1 \us31/U83  ( .A(\us31/n7 ), .B(\us31/n8 ), .S0(sa31[6]), .Y(sa32_sr[7]) );
  NOR2X4 \us31/U82  ( .A(\us31/n129 ), .B(sa31[2]), .Y(\us31/n43 ) );
  CLKINVX3 \us31/U81  ( .A(\us31/n14 ), .Y(\us31/n52 ) );
  OAI22XL \us31/U80  ( .A0(\us31/n201 ), .A1(\us31/n52 ), .B0(\us31/n202 ), 
        .B1(\us31/n114 ), .Y(\us31/n193 ) );
  CLKINVX3 \us31/U79  ( .A(sa31[5]), .Y(\us31/n252 ) );
  NOR2X2 \us31/U78  ( .A(\us31/n252 ), .B(\us31/n234 ), .Y(\us31/n55 ) );
  CLKINVX3 \us31/U77  ( .A(sa31[7]), .Y(\us31/n129 ) );
  NOR2X4 \us31/U76  ( .A(\us31/n129 ), .B(\us31/n69 ), .Y(\us31/n24 ) );
  AOI22XL \us31/U75  ( .A0(\us31/n70 ), .A1(\us31/n24 ), .B0(\us31/n96 ), .B1(
        \us31/n129 ), .Y(\us31/n241 ) );
  NOR2X2 \us31/U74  ( .A(\us31/n252 ), .B(sa31[0]), .Y(\us31/n89 ) );
  CLKINVX3 \us31/U73  ( .A(sa31[0]), .Y(\us31/n234 ) );
  NOR2X4 \us31/U72  ( .A(\us31/n69 ), .B(sa31[7]), .Y(\us31/n33 ) );
  INVX12 \us31/U71  ( .A(\us31/n33 ), .Y(\us31/n27 ) );
  CLKINVX3 \us31/U70  ( .A(\us31/n1 ), .Y(\us31/n6 ) );
  CLKINVX3 \us31/U69  ( .A(\us31/n1 ), .Y(\us31/n5 ) );
  INVXL \us31/U68  ( .A(\us31/n24 ), .Y(\us31/n36 ) );
  INVX4 \us31/U67  ( .A(\us31/n3 ), .Y(\us31/n4 ) );
  INVXL \us31/U66  ( .A(\us31/n36 ), .Y(\us31/n3 ) );
  INVX4 \us31/U65  ( .A(sa31[1]), .Y(\us31/n226 ) );
  INVX4 \us31/U64  ( .A(\us31/n43 ), .Y(\us31/n20 ) );
  AOI221X4 \us31/U63  ( .A0(\us31/n24 ), .A1(\us31/n82 ), .B0(\us31/n43 ), 
        .B1(\us31/n295 ), .C0(\us31/n173 ), .Y(\us31/n346 ) );
  AOI221X4 \us31/U62  ( .A0(\us31/n5 ), .A1(\us31/n96 ), .B0(\us31/n43 ), .B1(
        \us31/n239 ), .C0(\us31/n340 ), .Y(\us31/n336 ) );
  AOI222X4 \us31/U61  ( .A0(\us31/n59 ), .A1(\us31/n43 ), .B0(\us31/n6 ), .B1(
        \us31/n221 ), .C0(\us31/n222 ), .C1(\us31/n187 ), .Y(\us31/n218 ) );
  AOI222X4 \us31/U60  ( .A0(\us31/n123 ), .A1(\us31/n43 ), .B0(sa31[2]), .B1(
        \us31/n203 ), .C0(\us31/n6 ), .C1(\us31/n71 ), .Y(\us31/n202 ) );
  AOI221X4 \us31/U59  ( .A0(\us31/n314 ), .A1(\us31/n43 ), .B0(\us31/n160 ), 
        .B1(\us31/n24 ), .C0(\us31/n315 ), .Y(\us31/n307 ) );
  AOI221X4 \us31/U58  ( .A0(\us31/n43 ), .A1(\us31/n208 ), .B0(\us31/n76 ), 
        .B1(\us31/n24 ), .C0(\us31/n209 ), .Y(\us31/n207 ) );
  AOI221X4 \us31/U57  ( .A0(\us31/n43 ), .A1(\us31/n205 ), .B0(\us31/n32 ), 
        .B1(\us31/n6 ), .C0(\us31/n206 ), .Y(\us31/n201 ) );
  AOI221X4 \us31/U56  ( .A0(\us31/n43 ), .A1(\us31/n44 ), .B0(\us31/n45 ), 
        .B1(\us31/n24 ), .C0(\us31/n46 ), .Y(\us31/n9 ) );
  AOI22XL \us31/U55  ( .A0(\us31/n217 ), .A1(\us31/n43 ), .B0(\us31/n33 ), 
        .B1(\us31/n47 ), .Y(\us31/n216 ) );
  AOI22XL \us31/U54  ( .A0(\us31/n98 ), .A1(\us31/n43 ), .B0(\us31/n6 ), .B1(
        \us31/n99 ), .Y(\us31/n97 ) );
  AOI22XL \us31/U53  ( .A0(\us31/n82 ), .A1(\us31/n43 ), .B0(\us31/n83 ), .B1(
        \us31/n24 ), .Y(\us31/n81 ) );
  AOI2BB2XL \us31/U52  ( .B0(\us31/n43 ), .B1(\us31/n94 ), .A0N(\us31/n120 ), 
        .A1N(\us31/n4 ), .Y(\us31/n119 ) );
  AOI222X4 \us31/U51  ( .A0(\us31/n125 ), .A1(\us31/n33 ), .B0(\us31/n145 ), 
        .B1(\us31/n40 ), .C0(\us31/n43 ), .C1(\us31/n184 ), .Y(\us31/n183 ) );
  AOI22XL \us31/U50  ( .A0(\us31/n43 ), .A1(\us31/n303 ), .B0(\us31/n24 ), 
        .B1(\us31/n96 ), .Y(\us31/n358 ) );
  AOI22XL \us31/U49  ( .A0(\us31/n43 ), .A1(\us31/n100 ), .B0(\us31/n24 ), 
        .B1(\us31/n125 ), .Y(\us31/n124 ) );
  AOI21XL \us31/U48  ( .A0(\us31/n159 ), .A1(\us31/n43 ), .B0(\us31/n40 ), .Y(
        \us31/n262 ) );
  AOI22XL \us31/U47  ( .A0(\us31/n40 ), .A1(\us31/n94 ), .B0(\us31/n43 ), .B1(
        \us31/n187 ), .Y(\us31/n244 ) );
  AOI22XL \us31/U46  ( .A0(\us31/n184 ), .A1(\us31/n5 ), .B0(\us31/n198 ), 
        .B1(\us31/n43 ), .Y(\us31/n197 ) );
  NOR2XL \us31/U45  ( .A(\us31/n33 ), .B(\us31/n2 ), .Y(\us31/n302 ) );
  MXI2XL \us31/U44  ( .A(\us31/n2 ), .B(\us31/n6 ), .S0(\us31/n28 ), .Y(
        \us31/n311 ) );
  INVXL \us31/U43  ( .A(\us31/n20 ), .Y(\us31/n2 ) );
  INVX4 \us31/U42  ( .A(\us31/n6 ), .Y(\us31/n18 ) );
  AOI21XL \us31/U41  ( .A0(\us31/n18 ), .A1(\us31/n162 ), .B0(\us31/n25 ), .Y(
        \us31/n161 ) );
  INVX4 \us31/U40  ( .A(sa31[2]), .Y(\us31/n69 ) );
  NOR2X4 \us31/U39  ( .A(\us31/n226 ), .B(\us31/n4 ), .Y(\us31/n40 ) );
  CLKINVX3 \us31/U38  ( .A(sa31[3]), .Y(\us31/n136 ) );
  NOR2X2 \us31/U37  ( .A(\us31/n136 ), .B(sa31[4]), .Y(\us31/n145 ) );
  CLKINVX3 \us31/U36  ( .A(sa31[4]), .Y(\us31/n58 ) );
  NOR2X2 \us31/U35  ( .A(\us31/n58 ), .B(sa31[3]), .Y(\us31/n159 ) );
  NOR2X2 \us31/U34  ( .A(\us31/n136 ), .B(\us31/n58 ), .Y(\us31/n259 ) );
  NOR2X2 \us31/U33  ( .A(sa31[4]), .B(sa31[3]), .Y(\us31/n278 ) );
  NOR2X2 \us31/U32  ( .A(\us31/n259 ), .B(\us31/n278 ), .Y(\us31/n47 ) );
  CLKINVX3 \us31/U31  ( .A(\us31/n259 ), .Y(\us31/n44 ) );
  NOR2X2 \us31/U30  ( .A(\us31/n44 ), .B(sa31[1]), .Y(\us31/n137 ) );
  AOI21XL \us31/U29  ( .A0(\us31/n44 ), .A1(\us31/n111 ), .B0(\us31/n4 ), .Y(
        \us31/n177 ) );
  AOI22XL \us31/U28  ( .A0(\us31/n23 ), .A1(\us31/n24 ), .B0(\us31/n25 ), .B1(
        sa31[2]), .Y(\us31/n22 ) );
  AOI22XL \us31/U27  ( .A0(\us31/n33 ), .A1(sa31[3]), .B0(\us31/n24 ), .B1(
        \us31/n58 ), .Y(\us31/n277 ) );
  NAND2XL \us31/U26  ( .A(\us31/n198 ), .B(\us31/n24 ), .Y(\us31/n132 ) );
  OAI2BB2XL \us31/U25  ( .B0(\us31/n20 ), .B1(\us31/n111 ), .A0N(\us31/n125 ), 
        .A1N(\us31/n24 ), .Y(\us31/n220 ) );
  NAND2XL \us31/U24  ( .A(\us31/n111 ), .B(\us31/n101 ), .Y(\us31/n21 ) );
  NAND2XL \us31/U23  ( .A(\us31/n111 ), .B(\us31/n300 ), .Y(\us31/n187 ) );
  NAND2XL \us31/U22  ( .A(\us31/n111 ), .B(\us31/n121 ), .Y(\us31/n303 ) );
  AOI221XL \us31/U21  ( .A0(\us31/n43 ), .A1(\us31/n151 ), .B0(\us31/n25 ), 
        .B1(\us31/n69 ), .C0(\us31/n275 ), .Y(\us31/n274 ) );
  NOR2BXL \us31/U20  ( .AN(\us31/n101 ), .B(\us31/n25 ), .Y(\us31/n172 ) );
  NAND2X2 \us31/U19  ( .A(\us31/n58 ), .B(\us31/n226 ), .Y(\us31/n34 ) );
  OAI222X1 \us31/U18  ( .A0(\us31/n27 ), .A1(\us31/n34 ), .B0(\us31/n69 ), 
        .B1(\us31/n205 ), .C0(\us31/n20 ), .C1(\us31/n79 ), .Y(\us31/n260 ) );
  OAI222X1 \us31/U17  ( .A0(\us31/n20 ), .A1(\us31/n99 ), .B0(\us31/n27 ), 
        .B1(\us31/n101 ), .C0(\us31/n184 ), .C1(\us31/n4 ), .Y(\us31/n250 ) );
  OAI222X1 \us31/U16  ( .A0(\us31/n4 ), .A1(\us31/n37 ), .B0(\us31/n38 ), .B1(
        \us31/n20 ), .C0(sa31[4]), .C1(\us31/n39 ), .Y(\us31/n35 ) );
  AOI221X1 \us31/U15  ( .A0(\us31/n5 ), .A1(\us31/n19 ), .B0(\us31/n33 ), .B1(
        \us31/n34 ), .C0(\us31/n35 ), .Y(\us31/n11 ) );
  OR2X2 \us31/U14  ( .A(sa31[2]), .B(sa31[7]), .Y(\us31/n1 ) );
  AOI221XL \us31/U13  ( .A0(\us31/n70 ), .A1(\us31/n43 ), .B0(\us31/n24 ), 
        .B1(\us31/n71 ), .C0(\us31/n72 ), .Y(\us31/n53 ) );
  AOI221XL \us31/U12  ( .A0(\us31/n59 ), .A1(\us31/n33 ), .B0(\us31/n43 ), 
        .B1(\us31/n126 ), .C0(\us31/n127 ), .Y(\us31/n113 ) );
  AOI222XL \us31/U11  ( .A0(\us31/n185 ), .A1(\us31/n43 ), .B0(\us31/n186 ), 
        .B1(\us31/n187 ), .C0(\us31/n6 ), .C1(\us31/n188 ), .Y(\us31/n164 ) );
  AOI221X1 \us31/U10  ( .A0(\us31/n313 ), .A1(\us31/n5 ), .B0(\us31/n23 ), 
        .B1(\us31/n2 ), .C0(\us31/n328 ), .Y(\us31/n320 ) );
  AOI221X1 \us31/U9  ( .A0(\us31/n40 ), .A1(\us31/n136 ), .B0(\us31/n33 ), 
        .B1(\us31/n178 ), .C0(\us31/n338 ), .Y(\us31/n337 ) );
  AOI222XL \us31/U8  ( .A0(\us31/n278 ), .A1(\us31/n24 ), .B0(\us31/n42 ), 
        .B1(\us31/n33 ), .C0(\us31/n43 ), .C1(\us31/n136 ), .Y(\us31/n351 ) );
  AOI31X1 \us31/U7  ( .A0(sa31[2]), .A1(\us31/n58 ), .A2(sa31[1]), .B0(
        \us31/n40 ), .Y(\us31/n350 ) );
  AOI31X1 \us31/U6  ( .A0(\us31/n44 ), .A1(\us31/n129 ), .A2(\us31/n130 ), 
        .B0(\us31/n131 ), .Y(\us31/n128 ) );
  AOI221X1 \us31/U5  ( .A0(\us31/n40 ), .A1(\us31/n136 ), .B0(\us31/n33 ), 
        .B1(\us31/n47 ), .C0(\us31/n156 ), .Y(\us31/n141 ) );
  OAI32X1 \us31/U4  ( .A0(\us31/n18 ), .A1(sa31[1]), .A2(\us31/n159 ), .B0(
        sa31[4]), .B1(\us31/n182 ), .Y(\us31/n318 ) );
  OAI32X1 \us31/U3  ( .A0(\us31/n210 ), .A1(\us31/n145 ), .A2(\us31/n18 ), 
        .B0(\us31/n27 ), .B1(\us31/n211 ), .Y(\us31/n209 ) );
  AOI221X1 \us31/U2  ( .A0(\us31/n278 ), .A1(\us31/n40 ), .B0(\us31/n185 ), 
        .B1(\us31/n2 ), .C0(\us31/n279 ), .Y(\us31/n273 ) );
  AOI31XL \us31/U1  ( .A0(\us31/n79 ), .A1(\us31/n44 ), .A2(\us31/n2 ), .B0(
        \us31/n280 ), .Y(\us31/n339 ) );
  NAND2X1 \us32/U366  ( .A(\us32/n47 ), .B(\us32/n226 ), .Y(\us32/n189 ) );
  NOR2X1 \us32/U365  ( .A(\us32/n226 ), .B(sa32[3]), .Y(\us32/n242 ) );
  INVX1 \us32/U364  ( .A(\us32/n242 ), .Y(\us32/n205 ) );
  AND2X1 \us32/U363  ( .A(\us32/n189 ), .B(\us32/n205 ), .Y(\us32/n65 ) );
  NOR2X1 \us32/U362  ( .A(\us32/n226 ), .B(\us32/n47 ), .Y(\us32/n45 ) );
  NOR2X1 \us32/U361  ( .A(\us32/n259 ), .B(\us32/n45 ), .Y(\us32/n73 ) );
  NAND2BX1 \us32/U360  ( .AN(\us32/n73 ), .B(\us32/n6 ), .Y(\us32/n158 ) );
  NOR2X1 \us32/U359  ( .A(\us32/n226 ), .B(\us32/n159 ), .Y(\us32/n95 ) );
  INVX1 \us32/U358  ( .A(\us32/n95 ), .Y(\us32/n111 ) );
  NOR2X1 \us32/U357  ( .A(\us32/n145 ), .B(sa32[1]), .Y(\us32/n42 ) );
  INVX1 \us32/U356  ( .A(\us32/n42 ), .Y(\us32/n121 ) );
  INVX1 \us32/U355  ( .A(\us32/n47 ), .Y(\us32/n96 ) );
  OAI211X1 \us32/U354  ( .A0(\us32/n65 ), .A1(\us32/n27 ), .B0(\us32/n158 ), 
        .C0(\us32/n358 ), .Y(\us32/n355 ) );
  NOR2X1 \us32/U353  ( .A(\us32/n226 ), .B(\us32/n145 ), .Y(\us32/n59 ) );
  NOR2X1 \us32/U352  ( .A(\us32/n96 ), .B(\us32/n59 ), .Y(\us32/n271 ) );
  NOR2X1 \us32/U351  ( .A(\us32/n226 ), .B(\us32/n278 ), .Y(\us32/n217 ) );
  INVX1 \us32/U350  ( .A(\us32/n217 ), .Y(\us32/n150 ) );
  NAND2X1 \us32/U349  ( .A(\us32/n44 ), .B(\us32/n150 ), .Y(\us32/n147 ) );
  NAND2X1 \us32/U348  ( .A(sa32[4]), .B(\us32/n226 ), .Y(\us32/n101 ) );
  INVX1 \us32/U347  ( .A(\us32/n159 ), .Y(\us32/n188 ) );
  NOR2X1 \us32/U346  ( .A(\us32/n188 ), .B(\us32/n226 ), .Y(\us32/n25 ) );
  INVX1 \us32/U345  ( .A(\us32/n172 ), .Y(\us32/n107 ) );
  AOI22X1 \us32/U344  ( .A0(\us32/n33 ), .A1(\us32/n147 ), .B0(\us32/n24 ), 
        .B1(\us32/n107 ), .Y(\us32/n357 ) );
  OAI221XL \us32/U343  ( .A0(\us32/n18 ), .A1(\us32/n121 ), .B0(\us32/n271 ), 
        .B1(\us32/n20 ), .C0(\us32/n357 ), .Y(\us32/n356 ) );
  MXI2X1 \us32/U342  ( .A(\us32/n355 ), .B(\us32/n356 ), .S0(\us32/n252 ), .Y(
        \us32/n331 ) );
  INVX1 \us32/U341  ( .A(\us32/n59 ), .Y(\us32/n79 ) );
  AND2X1 \us32/U340  ( .A(\us32/n101 ), .B(\us32/n79 ), .Y(\us32/n325 ) );
  XNOR2X1 \us32/U339  ( .A(sa32[5]), .B(\us32/n226 ), .Y(\us32/n352 ) );
  NOR2X1 \us32/U338  ( .A(\us32/n226 ), .B(\us32/n136 ), .Y(\us32/n281 ) );
  INVX1 \us32/U337  ( .A(\us32/n281 ), .Y(\us32/n19 ) );
  NAND2X1 \us32/U336  ( .A(\us32/n145 ), .B(\us32/n226 ), .Y(\us32/n223 ) );
  AOI21X1 \us32/U335  ( .A0(\us32/n19 ), .A1(\us32/n223 ), .B0(\us32/n27 ), 
        .Y(\us32/n354 ) );
  AOI31X1 \us32/U334  ( .A0(\us32/n6 ), .A1(\us32/n352 ), .A2(\us32/n259 ), 
        .B0(\us32/n354 ), .Y(\us32/n353 ) );
  OAI221XL \us32/U333  ( .A0(\us32/n20 ), .A1(\us32/n34 ), .B0(\us32/n325 ), 
        .B1(\us32/n4 ), .C0(\us32/n353 ), .Y(\us32/n347 ) );
  INVX1 \us32/U332  ( .A(\us32/n352 ), .Y(\us32/n349 ) );
  NAND2X1 \us32/U331  ( .A(\us32/n278 ), .B(\us32/n6 ), .Y(\us32/n74 ) );
  OAI211X1 \us32/U330  ( .A0(\us32/n349 ), .A1(\us32/n74 ), .B0(\us32/n350 ), 
        .C0(\us32/n351 ), .Y(\us32/n348 ) );
  MXI2X1 \us32/U329  ( .A(\us32/n347 ), .B(\us32/n348 ), .S0(\us32/n252 ), .Y(
        \us32/n332 ) );
  NOR2X1 \us32/U328  ( .A(\us32/n44 ), .B(\us32/n226 ), .Y(\us32/n157 ) );
  INVX1 \us32/U327  ( .A(\us32/n157 ), .Y(\us32/n240 ) );
  NAND2X1 \us32/U326  ( .A(\us32/n240 ), .B(\us32/n189 ), .Y(\us32/n68 ) );
  NOR2X1 \us32/U325  ( .A(\us32/n20 ), .B(\us32/n159 ), .Y(\us32/n225 ) );
  NOR2X1 \us32/U324  ( .A(\us32/n225 ), .B(\us32/n40 ), .Y(\us32/n345 ) );
  INVX1 \us32/U323  ( .A(\us32/n278 ), .Y(\us32/n94 ) );
  NAND2X1 \us32/U322  ( .A(\us32/n94 ), .B(\us32/n226 ), .Y(\us32/n199 ) );
  NAND2X1 \us32/U321  ( .A(\us32/n199 ), .B(\us32/n205 ), .Y(\us32/n82 ) );
  NAND2X1 \us32/U320  ( .A(\us32/n19 ), .B(\us32/n199 ), .Y(\us32/n295 ) );
  NOR2X1 \us32/U319  ( .A(\us32/n226 ), .B(\us32/n259 ), .Y(\us32/n210 ) );
  NOR2X1 \us32/U318  ( .A(\us32/n27 ), .B(\us32/n210 ), .Y(\us32/n173 ) );
  MXI2X1 \us32/U317  ( .A(\us32/n345 ), .B(\us32/n346 ), .S0(\us32/n252 ), .Y(
        \us32/n342 ) );
  NOR2X1 \us32/U316  ( .A(sa32[1]), .B(sa32[3]), .Y(\us32/n163 ) );
  INVX1 \us32/U315  ( .A(\us32/n163 ), .Y(\us32/n37 ) );
  INVX1 \us32/U314  ( .A(\us32/n173 ), .Y(\us32/n344 ) );
  AOI21X1 \us32/U313  ( .A0(\us32/n240 ), .A1(\us32/n37 ), .B0(\us32/n344 ), 
        .Y(\us32/n343 ) );
  AOI211X1 \us32/U312  ( .A0(\us32/n5 ), .A1(\us32/n68 ), .B0(\us32/n342 ), 
        .C0(\us32/n343 ), .Y(\us32/n333 ) );
  NOR2X1 \us32/U311  ( .A(\us32/n18 ), .B(\us32/n226 ), .Y(\us32/n258 ) );
  NAND2X1 \us32/U310  ( .A(\us32/n278 ), .B(sa32[1]), .Y(\us32/n204 ) );
  NOR2X1 \us32/U309  ( .A(\us32/n188 ), .B(sa32[1]), .Y(\us32/n179 ) );
  INVX1 \us32/U308  ( .A(\us32/n179 ), .Y(\us32/n330 ) );
  NAND2X1 \us32/U307  ( .A(\us32/n204 ), .B(\us32/n330 ), .Y(\us32/n239 ) );
  NOR2X1 \us32/U306  ( .A(\us32/n136 ), .B(sa32[1]), .Y(\us32/n299 ) );
  NOR2X1 \us32/U305  ( .A(\us32/n299 ), .B(\us32/n210 ), .Y(\us32/n341 ) );
  OAI32X1 \us32/U304  ( .A0(\us32/n27 ), .A1(\us32/n278 ), .A2(\us32/n95 ), 
        .B0(\us32/n341 ), .B1(\us32/n4 ), .Y(\us32/n340 ) );
  INVX1 \us32/U303  ( .A(\us32/n45 ), .Y(\us32/n126 ) );
  NAND2X1 \us32/U302  ( .A(\us32/n126 ), .B(\us32/n101 ), .Y(\us32/n178 ) );
  NOR2X1 \us32/U301  ( .A(\us32/n18 ), .B(\us32/n136 ), .Y(\us32/n280 ) );
  OAI21XL \us32/U300  ( .A0(\us32/n4 ), .A1(\us32/n121 ), .B0(\us32/n339 ), 
        .Y(\us32/n338 ) );
  MXI2X1 \us32/U299  ( .A(\us32/n336 ), .B(\us32/n337 ), .S0(\us32/n252 ), .Y(
        \us32/n335 ) );
  NOR2X1 \us32/U298  ( .A(\us32/n258 ), .B(\us32/n335 ), .Y(\us32/n334 ) );
  MX4X1 \us32/U297  ( .A(\us32/n331 ), .B(\us32/n332 ), .C(\us32/n333 ), .D(
        \us32/n334 ), .S0(sa32[6]), .S1(\us32/n234 ), .Y(sa33_sr[0]) );
  INVX1 \us32/U296  ( .A(\us32/n299 ), .Y(\us32/n80 ) );
  NOR2X1 \us32/U295  ( .A(\us32/n111 ), .B(\us32/n18 ), .Y(\us32/n269 ) );
  INVX1 \us32/U294  ( .A(\us32/n269 ), .Y(\us32/n75 ) );
  OAI221XL \us32/U293  ( .A0(\us32/n18 ), .A1(\us32/n330 ), .B0(\us32/n20 ), 
        .B1(\us32/n80 ), .C0(\us32/n75 ), .Y(\us32/n329 ) );
  AOI221X1 \us32/U292  ( .A0(\us32/n325 ), .A1(\us32/n33 ), .B0(\us32/n24 ), 
        .B1(\us32/n303 ), .C0(\us32/n329 ), .Y(\us32/n319 ) );
  NOR2X1 \us32/U291  ( .A(\us32/n234 ), .B(sa32[5]), .Y(\us32/n14 ) );
  NOR2X1 \us32/U290  ( .A(\us32/n25 ), .B(\us32/n299 ), .Y(\us32/n313 ) );
  NAND2X1 \us32/U289  ( .A(\us32/n44 ), .B(\us32/n226 ), .Y(\us32/n300 ) );
  AND2X1 \us32/U288  ( .A(\us32/n300 ), .B(\us32/n240 ), .Y(\us32/n23 ) );
  OAI32X1 \us32/U287  ( .A0(\us32/n4 ), .A1(\us32/n145 ), .A2(\us32/n210 ), 
        .B0(\us32/n137 ), .B1(\us32/n27 ), .Y(\us32/n328 ) );
  NOR2X1 \us32/U286  ( .A(sa32[0]), .B(sa32[5]), .Y(\us32/n16 ) );
  INVX1 \us32/U285  ( .A(\us32/n16 ), .Y(\us32/n114 ) );
  INVX1 \us32/U284  ( .A(\us32/n145 ), .Y(\us32/n149 ) );
  NOR2X1 \us32/U283  ( .A(\us32/n47 ), .B(sa32[1]), .Y(\us32/n98 ) );
  INVX1 \us32/U282  ( .A(\us32/n98 ), .Y(\us32/n284 ) );
  OAI21XL \us32/U281  ( .A0(\us32/n69 ), .A1(\us32/n284 ), .B0(\us32/n27 ), 
        .Y(\us32/n327 ) );
  AOI31X1 \us32/U280  ( .A0(\us32/n111 ), .A1(\us32/n149 ), .A2(\us32/n327 ), 
        .B0(\us32/n225 ), .Y(\us32/n326 ) );
  OAI21XL \us32/U279  ( .A0(\us32/n325 ), .A1(\us32/n18 ), .B0(\us32/n326 ), 
        .Y(\us32/n322 ) );
  NAND2X1 \us32/U278  ( .A(\us32/n19 ), .B(\us32/n189 ), .Y(\us32/n71 ) );
  NOR2X1 \us32/U277  ( .A(\us32/n71 ), .B(\us32/n18 ), .Y(\us32/n135 ) );
  AOI21X1 \us32/U276  ( .A0(\us32/n40 ), .A1(sa32[4]), .B0(\us32/n135 ), .Y(
        \us32/n324 ) );
  OAI221XL \us32/U275  ( .A0(\us32/n47 ), .A1(\us32/n27 ), .B0(\us32/n65 ), 
        .B1(\us32/n20 ), .C0(\us32/n324 ), .Y(\us32/n323 ) );
  AOI22X1 \us32/U274  ( .A0(\us32/n55 ), .A1(\us32/n322 ), .B0(\us32/n89 ), 
        .B1(\us32/n323 ), .Y(\us32/n321 ) );
  OAI221XL \us32/U273  ( .A0(\us32/n319 ), .A1(\us32/n52 ), .B0(\us32/n320 ), 
        .B1(\us32/n114 ), .C0(\us32/n321 ), .Y(\us32/n304 ) );
  NOR2X1 \us32/U272  ( .A(\us32/n226 ), .B(\us32/n58 ), .Y(\us32/n290 ) );
  INVX1 \us32/U271  ( .A(\us32/n290 ), .Y(\us32/n200 ) );
  NAND2X1 \us32/U270  ( .A(\us32/n34 ), .B(\us32/n200 ), .Y(\us32/n120 ) );
  INVX1 \us32/U269  ( .A(\us32/n210 ), .Y(\us32/n100 ) );
  OAI221XL \us32/U268  ( .A0(\us32/n20 ), .A1(\us32/n100 ), .B0(sa32[3]), .B1(
        \us32/n4 ), .C0(\us32/n262 ), .Y(\us32/n317 ) );
  INVX1 \us32/U267  ( .A(\us32/n258 ), .Y(\us32/n182 ) );
  AOI211X1 \us32/U266  ( .A0(\us32/n33 ), .A1(\us32/n120 ), .B0(\us32/n317 ), 
        .C0(\us32/n318 ), .Y(\us32/n306 ) );
  NAND2X1 \us32/U265  ( .A(\us32/n100 ), .B(\us32/n199 ), .Y(\us32/n151 ) );
  INVX1 \us32/U264  ( .A(\us32/n151 ), .Y(\us32/n314 ) );
  NOR2X1 \us32/U263  ( .A(\us32/n45 ), .B(\us32/n163 ), .Y(\us32/n160 ) );
  INVX1 \us32/U262  ( .A(\us32/n295 ), .Y(\us32/n92 ) );
  AOI21X1 \us32/U261  ( .A0(sa32[1]), .A1(\us32/n58 ), .B0(\us32/n98 ), .Y(
        \us32/n316 ) );
  OAI22X1 \us32/U260  ( .A0(\us32/n92 ), .A1(\us32/n18 ), .B0(\us32/n316 ), 
        .B1(\us32/n27 ), .Y(\us32/n315 ) );
  NOR2X1 \us32/U259  ( .A(\us32/n149 ), .B(\us32/n226 ), .Y(\us32/n41 ) );
  INVX1 \us32/U258  ( .A(\us32/n41 ), .Y(\us32/n105 ) );
  NAND2X1 \us32/U257  ( .A(\us32/n284 ), .B(\us32/n105 ), .Y(\us32/n227 ) );
  AOI21X1 \us32/U256  ( .A0(\us32/n313 ), .A1(\us32/n33 ), .B0(\us32/n269 ), 
        .Y(\us32/n312 ) );
  OAI221XL \us32/U255  ( .A0(\us32/n149 ), .A1(\us32/n20 ), .B0(\us32/n4 ), 
        .B1(\us32/n227 ), .C0(\us32/n312 ), .Y(\us32/n309 ) );
  AOI21X1 \us32/U254  ( .A0(\us32/n226 ), .A1(\us32/n188 ), .B0(\us32/n242 ), 
        .Y(\us32/n185 ) );
  INVX1 \us32/U253  ( .A(\us32/n185 ), .Y(\us32/n48 ) );
  AND2X1 \us32/U252  ( .A(\us32/n223 ), .B(\us32/n240 ), .Y(\us32/n28 ) );
  OAI221XL \us32/U251  ( .A0(\us32/n27 ), .A1(\us32/n44 ), .B0(\us32/n4 ), 
        .B1(\us32/n48 ), .C0(\us32/n311 ), .Y(\us32/n310 ) );
  AOI22X1 \us32/U250  ( .A0(\us32/n89 ), .A1(\us32/n309 ), .B0(\us32/n55 ), 
        .B1(\us32/n310 ), .Y(\us32/n308 ) );
  OAI221XL \us32/U249  ( .A0(\us32/n306 ), .A1(\us32/n52 ), .B0(\us32/n307 ), 
        .B1(\us32/n114 ), .C0(\us32/n308 ), .Y(\us32/n305 ) );
  MX2X1 \us32/U248  ( .A(\us32/n304 ), .B(\us32/n305 ), .S0(sa32[6]), .Y(
        sa33_sr[1]) );
  INVX1 \us32/U247  ( .A(\us32/n187 ), .Y(\us32/n61 ) );
  MXI2X1 \us32/U246  ( .A(\us32/n303 ), .B(\us32/n61 ), .S0(\us32/n69 ), .Y(
        \us32/n301 ) );
  MXI2X1 \us32/U245  ( .A(\us32/n301 ), .B(\us32/n147 ), .S0(\us32/n302 ), .Y(
        \us32/n285 ) );
  NAND2X1 \us32/U244  ( .A(\us32/n200 ), .B(\us32/n300 ), .Y(\us32/n99 ) );
  INVX1 \us32/U243  ( .A(\us32/n99 ), .Y(\us32/n296 ) );
  NOR2X1 \us32/U242  ( .A(\us32/n299 ), .B(\us32/n242 ), .Y(\us32/n298 ) );
  NAND2X1 \us32/U241  ( .A(sa32[1]), .B(\us32/n47 ), .Y(\us32/n122 ) );
  NOR2X1 \us32/U240  ( .A(\us32/n159 ), .B(\us32/n217 ), .Y(\us32/n198 ) );
  OAI221XL \us32/U239  ( .A0(\us32/n298 ), .A1(\us32/n27 ), .B0(\us32/n20 ), 
        .B1(\us32/n122 ), .C0(\us32/n132 ), .Y(\us32/n297 ) );
  AOI221X1 \us32/U238  ( .A0(\us32/n225 ), .A1(\us32/n226 ), .B0(\us32/n296 ), 
        .B1(\us32/n6 ), .C0(\us32/n297 ), .Y(\us32/n291 ) );
  OAI2BB2X1 \us32/U237  ( .B0(\us32/n27 ), .B1(\us32/n295 ), .A0N(\us32/n34 ), 
        .A1N(\us32/n24 ), .Y(\us32/n293 ) );
  AOI21X1 \us32/U236  ( .A0(\us32/n101 ), .A1(\us32/n150 ), .B0(\us32/n20 ), 
        .Y(\us32/n294 ) );
  AOI211X1 \us32/U235  ( .A0(\us32/n5 ), .A1(\us32/n79 ), .B0(\us32/n293 ), 
        .C0(\us32/n294 ), .Y(\us32/n292 ) );
  INVX1 \us32/U234  ( .A(\us32/n89 ), .Y(\us32/n10 ) );
  OAI22X1 \us32/U233  ( .A0(\us32/n291 ), .A1(\us32/n114 ), .B0(\us32/n292 ), 
        .B1(\us32/n10 ), .Y(\us32/n286 ) );
  INVX1 \us32/U232  ( .A(\us32/n225 ), .Y(\us32/n288 ) );
  NAND2X1 \us32/U231  ( .A(\us32/n200 ), .B(\us32/n284 ), .Y(\us32/n102 ) );
  NOR2X1 \us32/U230  ( .A(\us32/n290 ), .B(\us32/n163 ), .Y(\us32/n184 ) );
  AOI22X1 \us32/U229  ( .A0(\us32/n102 ), .A1(\us32/n69 ), .B0(\us32/n184 ), 
        .B1(\us32/n33 ), .Y(\us32/n289 ) );
  AOI31X1 \us32/U228  ( .A0(\us32/n132 ), .A1(\us32/n288 ), .A2(\us32/n289 ), 
        .B0(\us32/n52 ), .Y(\us32/n287 ) );
  AOI211X1 \us32/U227  ( .A0(\us32/n285 ), .A1(\us32/n55 ), .B0(\us32/n286 ), 
        .C0(\us32/n287 ), .Y(\us32/n263 ) );
  NAND2X1 \us32/U226  ( .A(\us32/n284 ), .B(\us32/n122 ), .Y(\us32/n125 ) );
  NOR2X1 \us32/U225  ( .A(\us32/n199 ), .B(\us32/n4 ), .Y(\us32/n50 ) );
  AOI21X1 \us32/U224  ( .A0(\us32/n200 ), .A1(\us32/n223 ), .B0(\us32/n20 ), 
        .Y(\us32/n283 ) );
  AOI211X1 \us32/U223  ( .A0(\us32/n5 ), .A1(\us32/n125 ), .B0(\us32/n50 ), 
        .C0(\us32/n283 ), .Y(\us32/n282 ) );
  OAI221XL \us32/U222  ( .A0(\us32/n281 ), .A1(\us32/n27 ), .B0(\us32/n4 ), 
        .B1(\us32/n111 ), .C0(\us32/n282 ), .Y(\us32/n265 ) );
  INVX1 \us32/U221  ( .A(\us32/n280 ), .Y(\us32/n247 ) );
  NAND2X1 \us32/U220  ( .A(\us32/n41 ), .B(\us32/n33 ), .Y(\us32/n272 ) );
  OAI221XL \us32/U219  ( .A0(sa32[1]), .A1(\us32/n247 ), .B0(\us32/n4 ), .B1(
        \us32/n189 ), .C0(\us32/n272 ), .Y(\us32/n279 ) );
  NAND2X1 \us32/U218  ( .A(sa32[2]), .B(\us32/n149 ), .Y(\us32/n276 ) );
  XNOR2X1 \us32/U217  ( .A(\us32/n129 ), .B(sa32[1]), .Y(\us32/n155 ) );
  MXI2X1 \us32/U216  ( .A(\us32/n276 ), .B(\us32/n277 ), .S0(\us32/n155 ), .Y(
        \us32/n275 ) );
  OAI22X1 \us32/U215  ( .A0(\us32/n273 ), .A1(\us32/n10 ), .B0(\us32/n274 ), 
        .B1(\us32/n52 ), .Y(\us32/n266 ) );
  NOR2X1 \us32/U214  ( .A(\us32/n20 ), .B(\us32/n226 ), .Y(\us32/n176 ) );
  OAI21XL \us32/U213  ( .A0(\us32/n4 ), .A1(\us32/n271 ), .B0(\us32/n272 ), 
        .Y(\us32/n270 ) );
  OAI31X1 \us32/U212  ( .A0(\us32/n176 ), .A1(\us32/n269 ), .A2(\us32/n270 ), 
        .B0(\us32/n16 ), .Y(\us32/n268 ) );
  INVX1 \us32/U211  ( .A(\us32/n268 ), .Y(\us32/n267 ) );
  AOI211X1 \us32/U210  ( .A0(\us32/n55 ), .A1(\us32/n265 ), .B0(\us32/n266 ), 
        .C0(\us32/n267 ), .Y(\us32/n264 ) );
  MXI2X1 \us32/U209  ( .A(\us32/n263 ), .B(\us32/n264 ), .S0(sa32[6]), .Y(
        sa33_sr[2]) );
  NOR2X1 \us32/U208  ( .A(\us32/n94 ), .B(sa32[1]), .Y(\us32/n211 ) );
  INVX1 \us32/U207  ( .A(\us32/n262 ), .Y(\us32/n261 ) );
  AOI211X1 \us32/U206  ( .A0(\us32/n259 ), .A1(\us32/n24 ), .B0(\us32/n260 ), 
        .C0(\us32/n261 ), .Y(\us32/n255 ) );
  OAI22X1 \us32/U205  ( .A0(\us32/n20 ), .A1(\us32/n68 ), .B0(\us32/n27 ), 
        .B1(\us32/n37 ), .Y(\us32/n257 ) );
  NOR3X1 \us32/U204  ( .A(\us32/n257 ), .B(\us32/n258 ), .C(\us32/n50 ), .Y(
        \us32/n256 ) );
  MXI2X1 \us32/U203  ( .A(\us32/n255 ), .B(\us32/n256 ), .S0(\us32/n252 ), .Y(
        \us32/n254 ) );
  AOI221X1 \us32/U202  ( .A0(\us32/n211 ), .A1(\us32/n5 ), .B0(\us32/n40 ), 
        .B1(sa32[4]), .C0(\us32/n254 ), .Y(\us32/n248 ) );
  INVX1 \us32/U201  ( .A(\us32/n211 ), .Y(\us32/n106 ) );
  NAND2X1 \us32/U200  ( .A(\us32/n200 ), .B(\us32/n106 ), .Y(\us32/n83 ) );
  NAND2X1 \us32/U199  ( .A(\us32/n199 ), .B(\us32/n204 ), .Y(\us32/n169 ) );
  AOI2BB2X1 \us32/U198  ( .B0(\us32/n65 ), .B1(\us32/n24 ), .A0N(\us32/n169 ), 
        .A1N(\us32/n20 ), .Y(\us32/n253 ) );
  OAI221XL \us32/U197  ( .A0(\us32/n172 ), .A1(\us32/n18 ), .B0(\us32/n27 ), 
        .B1(\us32/n83 ), .C0(\us32/n253 ), .Y(\us32/n251 ) );
  MXI2X1 \us32/U196  ( .A(\us32/n250 ), .B(\us32/n251 ), .S0(\us32/n252 ), .Y(
        \us32/n249 ) );
  MXI2X1 \us32/U195  ( .A(\us32/n248 ), .B(\us32/n249 ), .S0(\us32/n234 ), .Y(
        \us32/n228 ) );
  OAI21XL \us32/U194  ( .A0(\us32/n58 ), .A1(\us32/n27 ), .B0(\us32/n247 ), 
        .Y(\us32/n245 ) );
  NOR2X1 \us32/U193  ( .A(sa32[7]), .B(\us32/n145 ), .Y(\us32/n246 ) );
  XNOR2X1 \us32/U192  ( .A(\us32/n69 ), .B(sa32[1]), .Y(\us32/n130 ) );
  MXI2X1 \us32/U191  ( .A(\us32/n245 ), .B(\us32/n246 ), .S0(\us32/n130 ), .Y(
        \us32/n243 ) );
  OAI211X1 \us32/U190  ( .A0(\us32/n4 ), .A1(\us32/n149 ), .B0(\us32/n243 ), 
        .C0(\us32/n244 ), .Y(\us32/n230 ) );
  NOR2X1 \us32/U189  ( .A(\us32/n242 ), .B(\us32/n137 ), .Y(\us32/n70 ) );
  OAI221XL \us32/U188  ( .A0(\us32/n159 ), .A1(\us32/n27 ), .B0(\us32/n20 ), 
        .B1(\us32/n34 ), .C0(\us32/n241 ), .Y(\us32/n231 ) );
  NAND2X1 \us32/U187  ( .A(\us32/n101 ), .B(\us32/n240 ), .Y(\us32/n76 ) );
  AOI21X1 \us32/U186  ( .A0(\us32/n122 ), .A1(\us32/n106 ), .B0(\us32/n129 ), 
        .Y(\us32/n237 ) );
  INVX1 \us32/U185  ( .A(\us32/n239 ), .Y(\us32/n238 ) );
  OAI21XL \us32/U184  ( .A0(\us32/n237 ), .A1(\us32/n43 ), .B0(\us32/n238 ), 
        .Y(\us32/n236 ) );
  OAI221XL \us32/U183  ( .A0(\us32/n18 ), .A1(\us32/n76 ), .B0(\us32/n59 ), 
        .B1(\us32/n27 ), .C0(\us32/n236 ), .Y(\us32/n232 ) );
  AOI2BB2X1 \us32/U182  ( .B0(\us32/n24 ), .B1(\us32/n187 ), .A0N(\us32/n227 ), 
        .A1N(\us32/n20 ), .Y(\us32/n235 ) );
  OAI211X1 \us32/U181  ( .A0(\us32/n27 ), .A1(\us32/n122 ), .B0(\us32/n158 ), 
        .C0(\us32/n235 ), .Y(\us32/n233 ) );
  MX4X1 \us32/U180  ( .A(\us32/n230 ), .B(\us32/n231 ), .C(\us32/n232 ), .D(
        \us32/n233 ), .S0(\us32/n234 ), .S1(sa32[5]), .Y(\us32/n229 ) );
  MX2X1 \us32/U179  ( .A(\us32/n228 ), .B(\us32/n229 ), .S0(sa32[6]), .Y(
        sa33_sr[3]) );
  NOR2BX1 \us32/U178  ( .AN(\us32/n204 ), .B(\us32/n137 ), .Y(\us32/n110 ) );
  INVX1 \us32/U177  ( .A(\us32/n110 ), .Y(\us32/n64 ) );
  AOI22X1 \us32/U176  ( .A0(\us32/n225 ), .A1(\us32/n226 ), .B0(\us32/n6 ), 
        .B1(\us32/n227 ), .Y(\us32/n224 ) );
  OAI221XL \us32/U175  ( .A0(\us32/n27 ), .A1(\us32/n64 ), .B0(\us32/n4 ), 
        .B1(\us32/n83 ), .C0(\us32/n224 ), .Y(\us32/n212 ) );
  NAND2X1 \us32/U174  ( .A(\us32/n34 ), .B(\us32/n204 ), .Y(\us32/n221 ) );
  OAI21XL \us32/U173  ( .A0(\us32/n69 ), .A1(\us32/n223 ), .B0(\us32/n27 ), 
        .Y(\us32/n222 ) );
  NOR2X1 \us32/U172  ( .A(\us32/n217 ), .B(\us32/n42 ), .Y(\us32/n208 ) );
  AOI211X1 \us32/U171  ( .A0(\us32/n208 ), .A1(\us32/n5 ), .B0(\us32/n220 ), 
        .C0(\us32/n173 ), .Y(\us32/n219 ) );
  OAI22X1 \us32/U170  ( .A0(\us32/n218 ), .A1(\us32/n10 ), .B0(\us32/n219 ), 
        .B1(\us32/n114 ), .Y(\us32/n213 ) );
  INVX1 \us32/U169  ( .A(\us32/n135 ), .Y(\us32/n215 ) );
  NOR2X1 \us32/U168  ( .A(\us32/n4 ), .B(\us32/n159 ), .Y(\us32/n31 ) );
  INVX1 \us32/U167  ( .A(\us32/n31 ), .Y(\us32/n196 ) );
  AOI31X1 \us32/U166  ( .A0(\us32/n215 ), .A1(\us32/n196 ), .A2(\us32/n216 ), 
        .B0(\us32/n52 ), .Y(\us32/n214 ) );
  AOI211X1 \us32/U165  ( .A0(\us32/n55 ), .A1(\us32/n212 ), .B0(\us32/n213 ), 
        .C0(\us32/n214 ), .Y(\us32/n190 ) );
  INVX1 \us32/U164  ( .A(\us32/n207 ), .Y(\us32/n192 ) );
  NOR2X1 \us32/U163  ( .A(\us32/n25 ), .B(\us32/n98 ), .Y(\us32/n32 ) );
  OAI22X1 \us32/U162  ( .A0(\us32/n28 ), .A1(\us32/n4 ), .B0(\us32/n188 ), 
        .B1(\us32/n27 ), .Y(\us32/n206 ) );
  NAND2X1 \us32/U161  ( .A(\us32/n204 ), .B(\us32/n80 ), .Y(\us32/n118 ) );
  INVX1 \us32/U160  ( .A(\us32/n118 ), .Y(\us32/n123 ) );
  NAND2X1 \us32/U159  ( .A(\us32/n94 ), .B(\us32/n79 ), .Y(\us32/n203 ) );
  OAI2BB1X1 \us32/U158  ( .A0N(\us32/n199 ), .A1N(\us32/n200 ), .B0(\us32/n33 ), .Y(\us32/n195 ) );
  INVX1 \us32/U157  ( .A(\us32/n55 ), .Y(\us32/n12 ) );
  AOI31X1 \us32/U156  ( .A0(\us32/n195 ), .A1(\us32/n196 ), .A2(\us32/n197 ), 
        .B0(\us32/n12 ), .Y(\us32/n194 ) );
  AOI211X1 \us32/U155  ( .A0(\us32/n89 ), .A1(\us32/n192 ), .B0(\us32/n193 ), 
        .C0(\us32/n194 ), .Y(\us32/n191 ) );
  MXI2X1 \us32/U154  ( .A(\us32/n190 ), .B(\us32/n191 ), .S0(sa32[6]), .Y(
        sa33_sr[4]) );
  OAI21XL \us32/U153  ( .A0(\us32/n69 ), .A1(\us32/n189 ), .B0(\us32/n27 ), 
        .Y(\us32/n186 ) );
  INVX1 \us32/U152  ( .A(\us32/n183 ), .Y(\us32/n180 ) );
  NAND2X1 \us32/U151  ( .A(\us32/n74 ), .B(\us32/n182 ), .Y(\us32/n181 ) );
  AOI211X1 \us32/U150  ( .A0(\us32/n179 ), .A1(\us32/n24 ), .B0(\us32/n180 ), 
        .C0(\us32/n181 ), .Y(\us32/n165 ) );
  INVX1 \us32/U149  ( .A(\us32/n178 ), .Y(\us32/n175 ) );
  AOI211X1 \us32/U148  ( .A0(\us32/n175 ), .A1(\us32/n5 ), .B0(\us32/n176 ), 
        .C0(\us32/n177 ), .Y(\us32/n174 ) );
  OAI221XL \us32/U147  ( .A0(\us32/n159 ), .A1(\us32/n27 ), .B0(\us32/n145 ), 
        .B1(\us32/n20 ), .C0(\us32/n174 ), .Y(\us32/n167 ) );
  MXI2X1 \us32/U146  ( .A(\us32/n40 ), .B(\us32/n173 ), .S0(\us32/n96 ), .Y(
        \us32/n170 ) );
  AOI22X1 \us32/U145  ( .A0(\us32/n137 ), .A1(\us32/n24 ), .B0(\us32/n172 ), 
        .B1(\us32/n6 ), .Y(\us32/n171 ) );
  OAI211X1 \us32/U144  ( .A0(\us32/n20 ), .A1(\us32/n169 ), .B0(\us32/n170 ), 
        .C0(\us32/n171 ), .Y(\us32/n168 ) );
  AOI22X1 \us32/U143  ( .A0(\us32/n89 ), .A1(\us32/n167 ), .B0(\us32/n55 ), 
        .B1(\us32/n168 ), .Y(\us32/n166 ) );
  OAI221XL \us32/U142  ( .A0(\us32/n164 ), .A1(\us32/n114 ), .B0(\us32/n165 ), 
        .B1(\us32/n52 ), .C0(\us32/n166 ), .Y(\us32/n138 ) );
  OAI21XL \us32/U141  ( .A0(\us32/n41 ), .A1(\us32/n163 ), .B0(\us32/n69 ), 
        .Y(\us32/n162 ) );
  AOI221X1 \us32/U140  ( .A0(\us32/n159 ), .A1(\us32/n24 ), .B0(\us32/n160 ), 
        .B1(\us32/n33 ), .C0(\us32/n161 ), .Y(\us32/n140 ) );
  OAI21XL \us32/U139  ( .A0(\us32/n157 ), .A1(\us32/n20 ), .B0(\us32/n158 ), 
        .Y(\us32/n156 ) );
  NOR2X1 \us32/U138  ( .A(\us32/n4 ), .B(\us32/n136 ), .Y(\us32/n153 ) );
  NOR2X1 \us32/U137  ( .A(\us32/n145 ), .B(\us32/n69 ), .Y(\us32/n154 ) );
  MXI2X1 \us32/U136  ( .A(\us32/n153 ), .B(\us32/n154 ), .S0(\us32/n155 ), .Y(
        \us32/n152 ) );
  OAI221XL \us32/U135  ( .A0(\us32/n110 ), .A1(\us32/n18 ), .B0(\us32/n20 ), 
        .B1(\us32/n151 ), .C0(\us32/n152 ), .Y(\us32/n143 ) );
  AOI21X1 \us32/U134  ( .A0(\us32/n149 ), .A1(\us32/n150 ), .B0(\us32/n18 ), 
        .Y(\us32/n148 ) );
  AOI2BB1X1 \us32/U133  ( .A0N(\us32/n147 ), .A1N(\us32/n27 ), .B0(\us32/n148 ), .Y(\us32/n146 ) );
  OAI221XL \us32/U132  ( .A0(\us32/n145 ), .A1(\us32/n20 ), .B0(\us32/n4 ), 
        .B1(\us32/n34 ), .C0(\us32/n146 ), .Y(\us32/n144 ) );
  AOI22X1 \us32/U131  ( .A0(\us32/n89 ), .A1(\us32/n143 ), .B0(\us32/n14 ), 
        .B1(\us32/n144 ), .Y(\us32/n142 ) );
  OAI221XL \us32/U130  ( .A0(\us32/n140 ), .A1(\us32/n12 ), .B0(\us32/n141 ), 
        .B1(\us32/n114 ), .C0(\us32/n142 ), .Y(\us32/n139 ) );
  MX2X1 \us32/U129  ( .A(\us32/n138 ), .B(\us32/n139 ), .S0(sa32[6]), .Y(
        sa33_sr[5]) );
  INVX1 \us32/U128  ( .A(\us32/n70 ), .Y(\us32/n133 ) );
  OAI22X1 \us32/U127  ( .A0(\us32/n4 ), .A1(\us32/n136 ), .B0(\us32/n137 ), 
        .B1(\us32/n27 ), .Y(\us32/n134 ) );
  AOI211X1 \us32/U126  ( .A0(\us32/n133 ), .A1(\us32/n69 ), .B0(\us32/n134 ), 
        .C0(\us32/n135 ), .Y(\us32/n112 ) );
  INVX1 \us32/U125  ( .A(\us32/n132 ), .Y(\us32/n131 ) );
  OAI21XL \us32/U124  ( .A0(\us32/n18 ), .A1(\us32/n37 ), .B0(\us32/n128 ), 
        .Y(\us32/n127 ) );
  OAI221XL \us32/U123  ( .A0(\us32/n18 ), .A1(\us32/n105 ), .B0(\us32/n123 ), 
        .B1(\us32/n27 ), .C0(\us32/n124 ), .Y(\us32/n116 ) );
  NAND2X1 \us32/U122  ( .A(\us32/n121 ), .B(\us32/n122 ), .Y(\us32/n30 ) );
  OAI221XL \us32/U121  ( .A0(\us32/n18 ), .A1(\us32/n118 ), .B0(\us32/n27 ), 
        .B1(\us32/n30 ), .C0(\us32/n119 ), .Y(\us32/n117 ) );
  AOI22X1 \us32/U120  ( .A0(\us32/n89 ), .A1(\us32/n116 ), .B0(\us32/n55 ), 
        .B1(\us32/n117 ), .Y(\us32/n115 ) );
  OAI221XL \us32/U119  ( .A0(\us32/n112 ), .A1(\us32/n52 ), .B0(\us32/n113 ), 
        .B1(\us32/n114 ), .C0(\us32/n115 ), .Y(\us32/n84 ) );
  OAI22X1 \us32/U118  ( .A0(\us32/n110 ), .A1(\us32/n4 ), .B0(\us32/n20 ), 
        .B1(\us32/n21 ), .Y(\us32/n108 ) );
  AOI21X1 \us32/U117  ( .A0(sa32[1]), .A1(\us32/n58 ), .B0(\us32/n27 ), .Y(
        \us32/n109 ) );
  AOI211X1 \us32/U116  ( .A0(\us32/n5 ), .A1(\us32/n107 ), .B0(\us32/n108 ), 
        .C0(\us32/n109 ), .Y(\us32/n86 ) );
  OAI22X1 \us32/U115  ( .A0(\us32/n45 ), .A1(\us32/n4 ), .B0(sa32[4]), .B1(
        \us32/n18 ), .Y(\us32/n103 ) );
  AOI21X1 \us32/U114  ( .A0(\us32/n105 ), .A1(\us32/n106 ), .B0(\us32/n20 ), 
        .Y(\us32/n104 ) );
  AOI211X1 \us32/U113  ( .A0(\us32/n33 ), .A1(\us32/n102 ), .B0(\us32/n103 ), 
        .C0(\us32/n104 ), .Y(\us32/n87 ) );
  NAND2X1 \us32/U112  ( .A(\us32/n100 ), .B(\us32/n101 ), .Y(\us32/n62 ) );
  OAI221XL \us32/U111  ( .A0(\us32/n27 ), .A1(\us32/n62 ), .B0(\us32/n4 ), 
        .B1(\us32/n21 ), .C0(\us32/n97 ), .Y(\us32/n90 ) );
  NOR3X1 \us32/U110  ( .A(\us32/n4 ), .B(\us32/n95 ), .C(\us32/n96 ), .Y(
        \us32/n67 ) );
  AOI31X1 \us32/U109  ( .A0(\us32/n79 ), .A1(\us32/n94 ), .A2(\us32/n6 ), .B0(
        \us32/n67 ), .Y(\us32/n93 ) );
  OAI221XL \us32/U108  ( .A0(\us32/n73 ), .A1(\us32/n27 ), .B0(\us32/n92 ), 
        .B1(\us32/n20 ), .C0(\us32/n93 ), .Y(\us32/n91 ) );
  AOI22X1 \us32/U107  ( .A0(\us32/n89 ), .A1(\us32/n90 ), .B0(\us32/n16 ), 
        .B1(\us32/n91 ), .Y(\us32/n88 ) );
  OAI221XL \us32/U106  ( .A0(\us32/n86 ), .A1(\us32/n52 ), .B0(\us32/n87 ), 
        .B1(\us32/n12 ), .C0(\us32/n88 ), .Y(\us32/n85 ) );
  MX2X1 \us32/U105  ( .A(\us32/n84 ), .B(\us32/n85 ), .S0(sa32[6]), .Y(
        sa33_sr[6]) );
  INVX1 \us32/U104  ( .A(\us32/n81 ), .Y(\us32/n77 ) );
  AOI21X1 \us32/U103  ( .A0(\us32/n79 ), .A1(\us32/n80 ), .B0(\us32/n27 ), .Y(
        \us32/n78 ) );
  AOI211X1 \us32/U102  ( .A0(\us32/n5 ), .A1(\us32/n76 ), .B0(\us32/n77 ), 
        .C0(\us32/n78 ), .Y(\us32/n51 ) );
  OAI211X1 \us32/U101  ( .A0(\us32/n73 ), .A1(\us32/n27 ), .B0(\us32/n74 ), 
        .C0(\us32/n75 ), .Y(\us32/n72 ) );
  AOI21X1 \us32/U100  ( .A0(\us32/n68 ), .A1(\us32/n69 ), .B0(\us32/n6 ), .Y(
        \us32/n63 ) );
  INVX1 \us32/U99  ( .A(\us32/n67 ), .Y(\us32/n66 ) );
  OAI221XL \us32/U98  ( .A0(\us32/n63 ), .A1(\us32/n64 ), .B0(\us32/n65 ), 
        .B1(\us32/n27 ), .C0(\us32/n66 ), .Y(\us32/n56 ) );
  AOI2BB2X1 \us32/U97  ( .B0(\us32/n61 ), .B1(\us32/n24 ), .A0N(\us32/n62 ), 
        .A1N(\us32/n20 ), .Y(\us32/n60 ) );
  OAI221XL \us32/U96  ( .A0(\us32/n58 ), .A1(\us32/n18 ), .B0(\us32/n59 ), 
        .B1(\us32/n27 ), .C0(\us32/n60 ), .Y(\us32/n57 ) );
  AOI22X1 \us32/U95  ( .A0(\us32/n55 ), .A1(\us32/n56 ), .B0(\us32/n16 ), .B1(
        \us32/n57 ), .Y(\us32/n54 ) );
  OAI221XL \us32/U94  ( .A0(\us32/n51 ), .A1(\us32/n52 ), .B0(\us32/n53 ), 
        .B1(\us32/n10 ), .C0(\us32/n54 ), .Y(\us32/n7 ) );
  INVX1 \us32/U93  ( .A(\us32/n50 ), .Y(\us32/n49 ) );
  OAI221XL \us32/U92  ( .A0(\us32/n47 ), .A1(\us32/n18 ), .B0(\us32/n27 ), 
        .B1(\us32/n48 ), .C0(\us32/n49 ), .Y(\us32/n46 ) );
  NOR2X1 \us32/U91  ( .A(\us32/n41 ), .B(\us32/n42 ), .Y(\us32/n38 ) );
  INVX1 \us32/U90  ( .A(\us32/n40 ), .Y(\us32/n39 ) );
  INVX1 \us32/U89  ( .A(\us32/n32 ), .Y(\us32/n26 ) );
  AOI21X1 \us32/U88  ( .A0(\us32/n5 ), .A1(\us32/n30 ), .B0(\us32/n31 ), .Y(
        \us32/n29 ) );
  OAI221XL \us32/U87  ( .A0(\us32/n26 ), .A1(\us32/n27 ), .B0(\us32/n28 ), 
        .B1(\us32/n20 ), .C0(\us32/n29 ), .Y(\us32/n15 ) );
  OAI221XL \us32/U86  ( .A0(\us32/n18 ), .A1(\us32/n19 ), .B0(\us32/n20 ), 
        .B1(\us32/n21 ), .C0(\us32/n22 ), .Y(\us32/n17 ) );
  AOI22X1 \us32/U85  ( .A0(\us32/n14 ), .A1(\us32/n15 ), .B0(\us32/n16 ), .B1(
        \us32/n17 ), .Y(\us32/n13 ) );
  OAI221XL \us32/U84  ( .A0(\us32/n9 ), .A1(\us32/n10 ), .B0(\us32/n11 ), .B1(
        \us32/n12 ), .C0(\us32/n13 ), .Y(\us32/n8 ) );
  MX2X1 \us32/U83  ( .A(\us32/n7 ), .B(\us32/n8 ), .S0(sa32[6]), .Y(sa33_sr[7]) );
  NOR2X4 \us32/U82  ( .A(\us32/n129 ), .B(sa32[2]), .Y(\us32/n43 ) );
  CLKINVX3 \us32/U81  ( .A(\us32/n14 ), .Y(\us32/n52 ) );
  OAI22XL \us32/U80  ( .A0(\us32/n201 ), .A1(\us32/n52 ), .B0(\us32/n202 ), 
        .B1(\us32/n114 ), .Y(\us32/n193 ) );
  CLKINVX3 \us32/U79  ( .A(sa32[5]), .Y(\us32/n252 ) );
  NOR2X2 \us32/U78  ( .A(\us32/n252 ), .B(\us32/n234 ), .Y(\us32/n55 ) );
  CLKINVX3 \us32/U77  ( .A(sa32[7]), .Y(\us32/n129 ) );
  NOR2X4 \us32/U76  ( .A(\us32/n129 ), .B(\us32/n69 ), .Y(\us32/n24 ) );
  AOI22XL \us32/U75  ( .A0(\us32/n70 ), .A1(\us32/n24 ), .B0(\us32/n96 ), .B1(
        \us32/n129 ), .Y(\us32/n241 ) );
  NOR2X2 \us32/U74  ( .A(\us32/n252 ), .B(sa32[0]), .Y(\us32/n89 ) );
  CLKINVX3 \us32/U73  ( .A(sa32[0]), .Y(\us32/n234 ) );
  NOR2X4 \us32/U72  ( .A(\us32/n69 ), .B(sa32[7]), .Y(\us32/n33 ) );
  INVX12 \us32/U71  ( .A(\us32/n33 ), .Y(\us32/n27 ) );
  CLKINVX3 \us32/U70  ( .A(\us32/n1 ), .Y(\us32/n6 ) );
  CLKINVX3 \us32/U69  ( .A(\us32/n1 ), .Y(\us32/n5 ) );
  INVXL \us32/U68  ( .A(\us32/n24 ), .Y(\us32/n36 ) );
  INVX4 \us32/U67  ( .A(\us32/n3 ), .Y(\us32/n4 ) );
  INVXL \us32/U66  ( .A(\us32/n36 ), .Y(\us32/n3 ) );
  INVX4 \us32/U65  ( .A(sa32[1]), .Y(\us32/n226 ) );
  INVX4 \us32/U64  ( .A(\us32/n43 ), .Y(\us32/n20 ) );
  AOI221X4 \us32/U63  ( .A0(\us32/n24 ), .A1(\us32/n82 ), .B0(\us32/n43 ), 
        .B1(\us32/n295 ), .C0(\us32/n173 ), .Y(\us32/n346 ) );
  AOI221X4 \us32/U62  ( .A0(\us32/n5 ), .A1(\us32/n96 ), .B0(\us32/n43 ), .B1(
        \us32/n239 ), .C0(\us32/n340 ), .Y(\us32/n336 ) );
  AOI222X4 \us32/U61  ( .A0(\us32/n59 ), .A1(\us32/n43 ), .B0(\us32/n6 ), .B1(
        \us32/n221 ), .C0(\us32/n222 ), .C1(\us32/n187 ), .Y(\us32/n218 ) );
  AOI222X4 \us32/U60  ( .A0(\us32/n123 ), .A1(\us32/n43 ), .B0(sa32[2]), .B1(
        \us32/n203 ), .C0(\us32/n6 ), .C1(\us32/n71 ), .Y(\us32/n202 ) );
  AOI221X4 \us32/U59  ( .A0(\us32/n314 ), .A1(\us32/n43 ), .B0(\us32/n160 ), 
        .B1(\us32/n24 ), .C0(\us32/n315 ), .Y(\us32/n307 ) );
  AOI221X4 \us32/U58  ( .A0(\us32/n43 ), .A1(\us32/n208 ), .B0(\us32/n76 ), 
        .B1(\us32/n24 ), .C0(\us32/n209 ), .Y(\us32/n207 ) );
  AOI221X4 \us32/U57  ( .A0(\us32/n43 ), .A1(\us32/n205 ), .B0(\us32/n32 ), 
        .B1(\us32/n6 ), .C0(\us32/n206 ), .Y(\us32/n201 ) );
  AOI221X4 \us32/U56  ( .A0(\us32/n43 ), .A1(\us32/n44 ), .B0(\us32/n45 ), 
        .B1(\us32/n24 ), .C0(\us32/n46 ), .Y(\us32/n9 ) );
  AOI22XL \us32/U55  ( .A0(\us32/n217 ), .A1(\us32/n43 ), .B0(\us32/n33 ), 
        .B1(\us32/n47 ), .Y(\us32/n216 ) );
  AOI22XL \us32/U54  ( .A0(\us32/n98 ), .A1(\us32/n43 ), .B0(\us32/n6 ), .B1(
        \us32/n99 ), .Y(\us32/n97 ) );
  AOI22XL \us32/U53  ( .A0(\us32/n82 ), .A1(\us32/n43 ), .B0(\us32/n83 ), .B1(
        \us32/n24 ), .Y(\us32/n81 ) );
  AOI2BB2XL \us32/U52  ( .B0(\us32/n43 ), .B1(\us32/n94 ), .A0N(\us32/n120 ), 
        .A1N(\us32/n4 ), .Y(\us32/n119 ) );
  AOI222X4 \us32/U51  ( .A0(\us32/n125 ), .A1(\us32/n33 ), .B0(\us32/n145 ), 
        .B1(\us32/n40 ), .C0(\us32/n43 ), .C1(\us32/n184 ), .Y(\us32/n183 ) );
  AOI22XL \us32/U50  ( .A0(\us32/n43 ), .A1(\us32/n303 ), .B0(\us32/n24 ), 
        .B1(\us32/n96 ), .Y(\us32/n358 ) );
  AOI22XL \us32/U49  ( .A0(\us32/n43 ), .A1(\us32/n100 ), .B0(\us32/n24 ), 
        .B1(\us32/n125 ), .Y(\us32/n124 ) );
  AOI21XL \us32/U48  ( .A0(\us32/n159 ), .A1(\us32/n43 ), .B0(\us32/n40 ), .Y(
        \us32/n262 ) );
  AOI22XL \us32/U47  ( .A0(\us32/n40 ), .A1(\us32/n94 ), .B0(\us32/n43 ), .B1(
        \us32/n187 ), .Y(\us32/n244 ) );
  AOI22XL \us32/U46  ( .A0(\us32/n184 ), .A1(\us32/n5 ), .B0(\us32/n198 ), 
        .B1(\us32/n43 ), .Y(\us32/n197 ) );
  NOR2XL \us32/U45  ( .A(\us32/n33 ), .B(\us32/n2 ), .Y(\us32/n302 ) );
  MXI2XL \us32/U44  ( .A(\us32/n2 ), .B(\us32/n6 ), .S0(\us32/n28 ), .Y(
        \us32/n311 ) );
  INVXL \us32/U43  ( .A(\us32/n20 ), .Y(\us32/n2 ) );
  INVX4 \us32/U42  ( .A(\us32/n6 ), .Y(\us32/n18 ) );
  AOI21XL \us32/U41  ( .A0(\us32/n18 ), .A1(\us32/n162 ), .B0(\us32/n25 ), .Y(
        \us32/n161 ) );
  INVX4 \us32/U40  ( .A(sa32[2]), .Y(\us32/n69 ) );
  NOR2X4 \us32/U39  ( .A(\us32/n226 ), .B(\us32/n4 ), .Y(\us32/n40 ) );
  CLKINVX3 \us32/U38  ( .A(sa32[3]), .Y(\us32/n136 ) );
  NOR2X2 \us32/U37  ( .A(\us32/n136 ), .B(sa32[4]), .Y(\us32/n145 ) );
  CLKINVX3 \us32/U36  ( .A(sa32[4]), .Y(\us32/n58 ) );
  NOR2X2 \us32/U35  ( .A(\us32/n58 ), .B(sa32[3]), .Y(\us32/n159 ) );
  NOR2X2 \us32/U34  ( .A(\us32/n136 ), .B(\us32/n58 ), .Y(\us32/n259 ) );
  NOR2X2 \us32/U33  ( .A(sa32[4]), .B(sa32[3]), .Y(\us32/n278 ) );
  NOR2X2 \us32/U32  ( .A(\us32/n259 ), .B(\us32/n278 ), .Y(\us32/n47 ) );
  CLKINVX3 \us32/U31  ( .A(\us32/n259 ), .Y(\us32/n44 ) );
  NOR2X2 \us32/U30  ( .A(\us32/n44 ), .B(sa32[1]), .Y(\us32/n137 ) );
  AOI21XL \us32/U29  ( .A0(\us32/n44 ), .A1(\us32/n111 ), .B0(\us32/n4 ), .Y(
        \us32/n177 ) );
  AOI22XL \us32/U28  ( .A0(\us32/n23 ), .A1(\us32/n24 ), .B0(\us32/n25 ), .B1(
        sa32[2]), .Y(\us32/n22 ) );
  AOI22XL \us32/U27  ( .A0(\us32/n33 ), .A1(sa32[3]), .B0(\us32/n24 ), .B1(
        \us32/n58 ), .Y(\us32/n277 ) );
  NAND2XL \us32/U26  ( .A(\us32/n198 ), .B(\us32/n24 ), .Y(\us32/n132 ) );
  OAI2BB2XL \us32/U25  ( .B0(\us32/n20 ), .B1(\us32/n111 ), .A0N(\us32/n125 ), 
        .A1N(\us32/n24 ), .Y(\us32/n220 ) );
  NAND2XL \us32/U24  ( .A(\us32/n111 ), .B(\us32/n101 ), .Y(\us32/n21 ) );
  NAND2XL \us32/U23  ( .A(\us32/n111 ), .B(\us32/n300 ), .Y(\us32/n187 ) );
  NAND2XL \us32/U22  ( .A(\us32/n111 ), .B(\us32/n121 ), .Y(\us32/n303 ) );
  AOI221XL \us32/U21  ( .A0(\us32/n43 ), .A1(\us32/n151 ), .B0(\us32/n25 ), 
        .B1(\us32/n69 ), .C0(\us32/n275 ), .Y(\us32/n274 ) );
  NOR2BXL \us32/U20  ( .AN(\us32/n101 ), .B(\us32/n25 ), .Y(\us32/n172 ) );
  NAND2X2 \us32/U19  ( .A(\us32/n58 ), .B(\us32/n226 ), .Y(\us32/n34 ) );
  OAI222X1 \us32/U18  ( .A0(\us32/n27 ), .A1(\us32/n34 ), .B0(\us32/n69 ), 
        .B1(\us32/n205 ), .C0(\us32/n20 ), .C1(\us32/n79 ), .Y(\us32/n260 ) );
  OAI222X1 \us32/U17  ( .A0(\us32/n20 ), .A1(\us32/n99 ), .B0(\us32/n27 ), 
        .B1(\us32/n101 ), .C0(\us32/n184 ), .C1(\us32/n4 ), .Y(\us32/n250 ) );
  OAI222X1 \us32/U16  ( .A0(\us32/n4 ), .A1(\us32/n37 ), .B0(\us32/n38 ), .B1(
        \us32/n20 ), .C0(sa32[4]), .C1(\us32/n39 ), .Y(\us32/n35 ) );
  AOI221X1 \us32/U15  ( .A0(\us32/n5 ), .A1(\us32/n19 ), .B0(\us32/n33 ), .B1(
        \us32/n34 ), .C0(\us32/n35 ), .Y(\us32/n11 ) );
  OR2X2 \us32/U14  ( .A(sa32[2]), .B(sa32[7]), .Y(\us32/n1 ) );
  AOI221XL \us32/U13  ( .A0(\us32/n70 ), .A1(\us32/n43 ), .B0(\us32/n24 ), 
        .B1(\us32/n71 ), .C0(\us32/n72 ), .Y(\us32/n53 ) );
  AOI221XL \us32/U12  ( .A0(\us32/n59 ), .A1(\us32/n33 ), .B0(\us32/n43 ), 
        .B1(\us32/n126 ), .C0(\us32/n127 ), .Y(\us32/n113 ) );
  AOI222XL \us32/U11  ( .A0(\us32/n185 ), .A1(\us32/n43 ), .B0(\us32/n186 ), 
        .B1(\us32/n187 ), .C0(\us32/n6 ), .C1(\us32/n188 ), .Y(\us32/n164 ) );
  AOI221X1 \us32/U10  ( .A0(\us32/n313 ), .A1(\us32/n5 ), .B0(\us32/n23 ), 
        .B1(\us32/n2 ), .C0(\us32/n328 ), .Y(\us32/n320 ) );
  AOI221X1 \us32/U9  ( .A0(\us32/n40 ), .A1(\us32/n136 ), .B0(\us32/n33 ), 
        .B1(\us32/n178 ), .C0(\us32/n338 ), .Y(\us32/n337 ) );
  AOI222XL \us32/U8  ( .A0(\us32/n278 ), .A1(\us32/n24 ), .B0(\us32/n42 ), 
        .B1(\us32/n33 ), .C0(\us32/n43 ), .C1(\us32/n136 ), .Y(\us32/n351 ) );
  AOI31X1 \us32/U7  ( .A0(sa32[2]), .A1(\us32/n58 ), .A2(sa32[1]), .B0(
        \us32/n40 ), .Y(\us32/n350 ) );
  AOI31X1 \us32/U6  ( .A0(\us32/n44 ), .A1(\us32/n129 ), .A2(\us32/n130 ), 
        .B0(\us32/n131 ), .Y(\us32/n128 ) );
  AOI221X1 \us32/U5  ( .A0(\us32/n40 ), .A1(\us32/n136 ), .B0(\us32/n33 ), 
        .B1(\us32/n47 ), .C0(\us32/n156 ), .Y(\us32/n141 ) );
  OAI32X1 \us32/U4  ( .A0(\us32/n18 ), .A1(sa32[1]), .A2(\us32/n159 ), .B0(
        sa32[4]), .B1(\us32/n182 ), .Y(\us32/n318 ) );
  OAI32X1 \us32/U3  ( .A0(\us32/n210 ), .A1(\us32/n145 ), .A2(\us32/n18 ), 
        .B0(\us32/n27 ), .B1(\us32/n211 ), .Y(\us32/n209 ) );
  AOI221X1 \us32/U2  ( .A0(\us32/n278 ), .A1(\us32/n40 ), .B0(\us32/n185 ), 
        .B1(\us32/n2 ), .C0(\us32/n279 ), .Y(\us32/n273 ) );
  AOI31XL \us32/U1  ( .A0(\us32/n79 ), .A1(\us32/n44 ), .A2(\us32/n2 ), .B0(
        \us32/n280 ), .Y(\us32/n339 ) );
  NAND2X1 \us33/U366  ( .A(\us33/n47 ), .B(\us33/n226 ), .Y(\us33/n189 ) );
  NOR2X1 \us33/U365  ( .A(\us33/n226 ), .B(sa33[3]), .Y(\us33/n242 ) );
  INVX1 \us33/U364  ( .A(\us33/n242 ), .Y(\us33/n205 ) );
  AND2X1 \us33/U363  ( .A(\us33/n189 ), .B(\us33/n205 ), .Y(\us33/n65 ) );
  NOR2X1 \us33/U362  ( .A(\us33/n226 ), .B(\us33/n47 ), .Y(\us33/n45 ) );
  NOR2X1 \us33/U361  ( .A(\us33/n259 ), .B(\us33/n45 ), .Y(\us33/n73 ) );
  NAND2BX1 \us33/U360  ( .AN(\us33/n73 ), .B(\us33/n6 ), .Y(\us33/n158 ) );
  NOR2X1 \us33/U359  ( .A(\us33/n226 ), .B(\us33/n159 ), .Y(\us33/n95 ) );
  INVX1 \us33/U358  ( .A(\us33/n95 ), .Y(\us33/n111 ) );
  NOR2X1 \us33/U357  ( .A(\us33/n145 ), .B(sa33[1]), .Y(\us33/n42 ) );
  INVX1 \us33/U356  ( .A(\us33/n42 ), .Y(\us33/n121 ) );
  INVX1 \us33/U355  ( .A(\us33/n47 ), .Y(\us33/n96 ) );
  OAI211X1 \us33/U354  ( .A0(\us33/n65 ), .A1(\us33/n27 ), .B0(\us33/n158 ), 
        .C0(\us33/n358 ), .Y(\us33/n355 ) );
  NOR2X1 \us33/U353  ( .A(\us33/n226 ), .B(\us33/n145 ), .Y(\us33/n59 ) );
  NOR2X1 \us33/U352  ( .A(\us33/n96 ), .B(\us33/n59 ), .Y(\us33/n271 ) );
  NOR2X1 \us33/U351  ( .A(\us33/n226 ), .B(\us33/n278 ), .Y(\us33/n217 ) );
  INVX1 \us33/U350  ( .A(\us33/n217 ), .Y(\us33/n150 ) );
  NAND2X1 \us33/U349  ( .A(\us33/n44 ), .B(\us33/n150 ), .Y(\us33/n147 ) );
  NAND2X1 \us33/U348  ( .A(sa33[4]), .B(\us33/n226 ), .Y(\us33/n101 ) );
  INVX1 \us33/U347  ( .A(\us33/n159 ), .Y(\us33/n188 ) );
  NOR2X1 \us33/U346  ( .A(\us33/n188 ), .B(\us33/n226 ), .Y(\us33/n25 ) );
  INVX1 \us33/U345  ( .A(\us33/n172 ), .Y(\us33/n107 ) );
  AOI22X1 \us33/U344  ( .A0(\us33/n33 ), .A1(\us33/n147 ), .B0(\us33/n24 ), 
        .B1(\us33/n107 ), .Y(\us33/n357 ) );
  OAI221XL \us33/U343  ( .A0(\us33/n18 ), .A1(\us33/n121 ), .B0(\us33/n271 ), 
        .B1(\us33/n20 ), .C0(\us33/n357 ), .Y(\us33/n356 ) );
  MXI2X1 \us33/U342  ( .A(\us33/n355 ), .B(\us33/n356 ), .S0(\us33/n252 ), .Y(
        \us33/n331 ) );
  INVX1 \us33/U341  ( .A(\us33/n59 ), .Y(\us33/n79 ) );
  AND2X1 \us33/U340  ( .A(\us33/n101 ), .B(\us33/n79 ), .Y(\us33/n325 ) );
  XNOR2X1 \us33/U339  ( .A(sa33[5]), .B(\us33/n226 ), .Y(\us33/n352 ) );
  NOR2X1 \us33/U338  ( .A(\us33/n226 ), .B(\us33/n136 ), .Y(\us33/n281 ) );
  INVX1 \us33/U337  ( .A(\us33/n281 ), .Y(\us33/n19 ) );
  NAND2X1 \us33/U336  ( .A(\us33/n145 ), .B(\us33/n226 ), .Y(\us33/n223 ) );
  AOI21X1 \us33/U335  ( .A0(\us33/n19 ), .A1(\us33/n223 ), .B0(\us33/n27 ), 
        .Y(\us33/n354 ) );
  AOI31X1 \us33/U334  ( .A0(\us33/n6 ), .A1(\us33/n352 ), .A2(\us33/n259 ), 
        .B0(\us33/n354 ), .Y(\us33/n353 ) );
  OAI221XL \us33/U333  ( .A0(\us33/n20 ), .A1(\us33/n34 ), .B0(\us33/n325 ), 
        .B1(\us33/n4 ), .C0(\us33/n353 ), .Y(\us33/n347 ) );
  INVX1 \us33/U332  ( .A(\us33/n352 ), .Y(\us33/n349 ) );
  NAND2X1 \us33/U331  ( .A(\us33/n278 ), .B(\us33/n6 ), .Y(\us33/n74 ) );
  OAI211X1 \us33/U330  ( .A0(\us33/n349 ), .A1(\us33/n74 ), .B0(\us33/n350 ), 
        .C0(\us33/n351 ), .Y(\us33/n348 ) );
  MXI2X1 \us33/U329  ( .A(\us33/n347 ), .B(\us33/n348 ), .S0(\us33/n252 ), .Y(
        \us33/n332 ) );
  NOR2X1 \us33/U328  ( .A(\us33/n44 ), .B(\us33/n226 ), .Y(\us33/n157 ) );
  INVX1 \us33/U327  ( .A(\us33/n157 ), .Y(\us33/n240 ) );
  NAND2X1 \us33/U326  ( .A(\us33/n240 ), .B(\us33/n189 ), .Y(\us33/n68 ) );
  NOR2X1 \us33/U325  ( .A(\us33/n20 ), .B(\us33/n159 ), .Y(\us33/n225 ) );
  NOR2X1 \us33/U324  ( .A(\us33/n225 ), .B(\us33/n40 ), .Y(\us33/n345 ) );
  INVX1 \us33/U323  ( .A(\us33/n278 ), .Y(\us33/n94 ) );
  NAND2X1 \us33/U322  ( .A(\us33/n94 ), .B(\us33/n226 ), .Y(\us33/n199 ) );
  NAND2X1 \us33/U321  ( .A(\us33/n199 ), .B(\us33/n205 ), .Y(\us33/n82 ) );
  NAND2X1 \us33/U320  ( .A(\us33/n19 ), .B(\us33/n199 ), .Y(\us33/n295 ) );
  NOR2X1 \us33/U319  ( .A(\us33/n226 ), .B(\us33/n259 ), .Y(\us33/n210 ) );
  NOR2X1 \us33/U318  ( .A(\us33/n27 ), .B(\us33/n210 ), .Y(\us33/n173 ) );
  MXI2X1 \us33/U317  ( .A(\us33/n345 ), .B(\us33/n346 ), .S0(\us33/n252 ), .Y(
        \us33/n342 ) );
  NOR2X1 \us33/U316  ( .A(sa33[1]), .B(sa33[3]), .Y(\us33/n163 ) );
  INVX1 \us33/U315  ( .A(\us33/n163 ), .Y(\us33/n37 ) );
  INVX1 \us33/U314  ( .A(\us33/n173 ), .Y(\us33/n344 ) );
  AOI21X1 \us33/U313  ( .A0(\us33/n240 ), .A1(\us33/n37 ), .B0(\us33/n344 ), 
        .Y(\us33/n343 ) );
  AOI211X1 \us33/U312  ( .A0(\us33/n5 ), .A1(\us33/n68 ), .B0(\us33/n342 ), 
        .C0(\us33/n343 ), .Y(\us33/n333 ) );
  NOR2X1 \us33/U311  ( .A(\us33/n18 ), .B(\us33/n226 ), .Y(\us33/n258 ) );
  NAND2X1 \us33/U310  ( .A(\us33/n278 ), .B(sa33[1]), .Y(\us33/n204 ) );
  NOR2X1 \us33/U309  ( .A(\us33/n188 ), .B(sa33[1]), .Y(\us33/n179 ) );
  INVX1 \us33/U308  ( .A(\us33/n179 ), .Y(\us33/n330 ) );
  NAND2X1 \us33/U307  ( .A(\us33/n204 ), .B(\us33/n330 ), .Y(\us33/n239 ) );
  NOR2X1 \us33/U306  ( .A(\us33/n136 ), .B(sa33[1]), .Y(\us33/n299 ) );
  NOR2X1 \us33/U305  ( .A(\us33/n299 ), .B(\us33/n210 ), .Y(\us33/n341 ) );
  OAI32X1 \us33/U304  ( .A0(\us33/n27 ), .A1(\us33/n278 ), .A2(\us33/n95 ), 
        .B0(\us33/n341 ), .B1(\us33/n4 ), .Y(\us33/n340 ) );
  INVX1 \us33/U303  ( .A(\us33/n45 ), .Y(\us33/n126 ) );
  NAND2X1 \us33/U302  ( .A(\us33/n126 ), .B(\us33/n101 ), .Y(\us33/n178 ) );
  NOR2X1 \us33/U301  ( .A(\us33/n18 ), .B(\us33/n136 ), .Y(\us33/n280 ) );
  OAI21XL \us33/U300  ( .A0(\us33/n4 ), .A1(\us33/n121 ), .B0(\us33/n339 ), 
        .Y(\us33/n338 ) );
  MXI2X1 \us33/U299  ( .A(\us33/n336 ), .B(\us33/n337 ), .S0(\us33/n252 ), .Y(
        \us33/n335 ) );
  NOR2X1 \us33/U298  ( .A(\us33/n258 ), .B(\us33/n335 ), .Y(\us33/n334 ) );
  MX4X1 \us33/U297  ( .A(\us33/n331 ), .B(\us33/n332 ), .C(\us33/n333 ), .D(
        \us33/n334 ), .S0(sa33[6]), .S1(\us33/n234 ), .Y(sa30_sr[0]) );
  INVX1 \us33/U296  ( .A(\us33/n299 ), .Y(\us33/n80 ) );
  NOR2X1 \us33/U295  ( .A(\us33/n111 ), .B(\us33/n18 ), .Y(\us33/n269 ) );
  INVX1 \us33/U294  ( .A(\us33/n269 ), .Y(\us33/n75 ) );
  OAI221XL \us33/U293  ( .A0(\us33/n18 ), .A1(\us33/n330 ), .B0(\us33/n20 ), 
        .B1(\us33/n80 ), .C0(\us33/n75 ), .Y(\us33/n329 ) );
  AOI221X1 \us33/U292  ( .A0(\us33/n325 ), .A1(\us33/n33 ), .B0(\us33/n24 ), 
        .B1(\us33/n303 ), .C0(\us33/n329 ), .Y(\us33/n319 ) );
  NOR2X1 \us33/U291  ( .A(\us33/n234 ), .B(sa33[5]), .Y(\us33/n14 ) );
  NOR2X1 \us33/U290  ( .A(\us33/n25 ), .B(\us33/n299 ), .Y(\us33/n313 ) );
  NAND2X1 \us33/U289  ( .A(\us33/n44 ), .B(\us33/n226 ), .Y(\us33/n300 ) );
  AND2X1 \us33/U288  ( .A(\us33/n300 ), .B(\us33/n240 ), .Y(\us33/n23 ) );
  OAI32X1 \us33/U287  ( .A0(\us33/n4 ), .A1(\us33/n145 ), .A2(\us33/n210 ), 
        .B0(\us33/n137 ), .B1(\us33/n27 ), .Y(\us33/n328 ) );
  NOR2X1 \us33/U286  ( .A(sa33[0]), .B(sa33[5]), .Y(\us33/n16 ) );
  INVX1 \us33/U285  ( .A(\us33/n16 ), .Y(\us33/n114 ) );
  INVX1 \us33/U284  ( .A(\us33/n145 ), .Y(\us33/n149 ) );
  NOR2X1 \us33/U283  ( .A(\us33/n47 ), .B(sa33[1]), .Y(\us33/n98 ) );
  INVX1 \us33/U282  ( .A(\us33/n98 ), .Y(\us33/n284 ) );
  OAI21XL \us33/U281  ( .A0(\us33/n69 ), .A1(\us33/n284 ), .B0(\us33/n27 ), 
        .Y(\us33/n327 ) );
  AOI31X1 \us33/U280  ( .A0(\us33/n111 ), .A1(\us33/n149 ), .A2(\us33/n327 ), 
        .B0(\us33/n225 ), .Y(\us33/n326 ) );
  OAI21XL \us33/U279  ( .A0(\us33/n325 ), .A1(\us33/n18 ), .B0(\us33/n326 ), 
        .Y(\us33/n322 ) );
  NAND2X1 \us33/U278  ( .A(\us33/n19 ), .B(\us33/n189 ), .Y(\us33/n71 ) );
  NOR2X1 \us33/U277  ( .A(\us33/n71 ), .B(\us33/n18 ), .Y(\us33/n135 ) );
  AOI21X1 \us33/U276  ( .A0(\us33/n40 ), .A1(sa33[4]), .B0(\us33/n135 ), .Y(
        \us33/n324 ) );
  OAI221XL \us33/U275  ( .A0(\us33/n47 ), .A1(\us33/n27 ), .B0(\us33/n65 ), 
        .B1(\us33/n20 ), .C0(\us33/n324 ), .Y(\us33/n323 ) );
  AOI22X1 \us33/U274  ( .A0(\us33/n55 ), .A1(\us33/n322 ), .B0(\us33/n89 ), 
        .B1(\us33/n323 ), .Y(\us33/n321 ) );
  OAI221XL \us33/U273  ( .A0(\us33/n319 ), .A1(\us33/n52 ), .B0(\us33/n320 ), 
        .B1(\us33/n114 ), .C0(\us33/n321 ), .Y(\us33/n304 ) );
  NOR2X1 \us33/U272  ( .A(\us33/n226 ), .B(\us33/n58 ), .Y(\us33/n290 ) );
  INVX1 \us33/U271  ( .A(\us33/n290 ), .Y(\us33/n200 ) );
  NAND2X1 \us33/U270  ( .A(\us33/n34 ), .B(\us33/n200 ), .Y(\us33/n120 ) );
  INVX1 \us33/U269  ( .A(\us33/n210 ), .Y(\us33/n100 ) );
  OAI221XL \us33/U268  ( .A0(\us33/n20 ), .A1(\us33/n100 ), .B0(sa33[3]), .B1(
        \us33/n4 ), .C0(\us33/n262 ), .Y(\us33/n317 ) );
  INVX1 \us33/U267  ( .A(\us33/n258 ), .Y(\us33/n182 ) );
  AOI211X1 \us33/U266  ( .A0(\us33/n33 ), .A1(\us33/n120 ), .B0(\us33/n317 ), 
        .C0(\us33/n318 ), .Y(\us33/n306 ) );
  NAND2X1 \us33/U265  ( .A(\us33/n100 ), .B(\us33/n199 ), .Y(\us33/n151 ) );
  INVX1 \us33/U264  ( .A(\us33/n151 ), .Y(\us33/n314 ) );
  NOR2X1 \us33/U263  ( .A(\us33/n45 ), .B(\us33/n163 ), .Y(\us33/n160 ) );
  INVX1 \us33/U262  ( .A(\us33/n295 ), .Y(\us33/n92 ) );
  AOI21X1 \us33/U261  ( .A0(sa33[1]), .A1(\us33/n58 ), .B0(\us33/n98 ), .Y(
        \us33/n316 ) );
  OAI22X1 \us33/U260  ( .A0(\us33/n92 ), .A1(\us33/n18 ), .B0(\us33/n316 ), 
        .B1(\us33/n27 ), .Y(\us33/n315 ) );
  NOR2X1 \us33/U259  ( .A(\us33/n149 ), .B(\us33/n226 ), .Y(\us33/n41 ) );
  INVX1 \us33/U258  ( .A(\us33/n41 ), .Y(\us33/n105 ) );
  NAND2X1 \us33/U257  ( .A(\us33/n284 ), .B(\us33/n105 ), .Y(\us33/n227 ) );
  AOI21X1 \us33/U256  ( .A0(\us33/n313 ), .A1(\us33/n33 ), .B0(\us33/n269 ), 
        .Y(\us33/n312 ) );
  OAI221XL \us33/U255  ( .A0(\us33/n149 ), .A1(\us33/n20 ), .B0(\us33/n4 ), 
        .B1(\us33/n227 ), .C0(\us33/n312 ), .Y(\us33/n309 ) );
  AOI21X1 \us33/U254  ( .A0(\us33/n226 ), .A1(\us33/n188 ), .B0(\us33/n242 ), 
        .Y(\us33/n185 ) );
  INVX1 \us33/U253  ( .A(\us33/n185 ), .Y(\us33/n48 ) );
  AND2X1 \us33/U252  ( .A(\us33/n223 ), .B(\us33/n240 ), .Y(\us33/n28 ) );
  OAI221XL \us33/U251  ( .A0(\us33/n27 ), .A1(\us33/n44 ), .B0(\us33/n4 ), 
        .B1(\us33/n48 ), .C0(\us33/n311 ), .Y(\us33/n310 ) );
  AOI22X1 \us33/U250  ( .A0(\us33/n89 ), .A1(\us33/n309 ), .B0(\us33/n55 ), 
        .B1(\us33/n310 ), .Y(\us33/n308 ) );
  OAI221XL \us33/U249  ( .A0(\us33/n306 ), .A1(\us33/n52 ), .B0(\us33/n307 ), 
        .B1(\us33/n114 ), .C0(\us33/n308 ), .Y(\us33/n305 ) );
  MX2X1 \us33/U248  ( .A(\us33/n304 ), .B(\us33/n305 ), .S0(sa33[6]), .Y(
        sa30_sr[1]) );
  INVX1 \us33/U247  ( .A(\us33/n187 ), .Y(\us33/n61 ) );
  MXI2X1 \us33/U246  ( .A(\us33/n303 ), .B(\us33/n61 ), .S0(\us33/n69 ), .Y(
        \us33/n301 ) );
  MXI2X1 \us33/U245  ( .A(\us33/n301 ), .B(\us33/n147 ), .S0(\us33/n302 ), .Y(
        \us33/n285 ) );
  NAND2X1 \us33/U244  ( .A(\us33/n200 ), .B(\us33/n300 ), .Y(\us33/n99 ) );
  INVX1 \us33/U243  ( .A(\us33/n99 ), .Y(\us33/n296 ) );
  NOR2X1 \us33/U242  ( .A(\us33/n299 ), .B(\us33/n242 ), .Y(\us33/n298 ) );
  NAND2X1 \us33/U241  ( .A(sa33[1]), .B(\us33/n47 ), .Y(\us33/n122 ) );
  NOR2X1 \us33/U240  ( .A(\us33/n159 ), .B(\us33/n217 ), .Y(\us33/n198 ) );
  OAI221XL \us33/U239  ( .A0(\us33/n298 ), .A1(\us33/n27 ), .B0(\us33/n20 ), 
        .B1(\us33/n122 ), .C0(\us33/n132 ), .Y(\us33/n297 ) );
  AOI221X1 \us33/U238  ( .A0(\us33/n225 ), .A1(\us33/n226 ), .B0(\us33/n296 ), 
        .B1(\us33/n6 ), .C0(\us33/n297 ), .Y(\us33/n291 ) );
  OAI2BB2X1 \us33/U237  ( .B0(\us33/n27 ), .B1(\us33/n295 ), .A0N(\us33/n34 ), 
        .A1N(\us33/n24 ), .Y(\us33/n293 ) );
  AOI21X1 \us33/U236  ( .A0(\us33/n101 ), .A1(\us33/n150 ), .B0(\us33/n20 ), 
        .Y(\us33/n294 ) );
  AOI211X1 \us33/U235  ( .A0(\us33/n5 ), .A1(\us33/n79 ), .B0(\us33/n293 ), 
        .C0(\us33/n294 ), .Y(\us33/n292 ) );
  INVX1 \us33/U234  ( .A(\us33/n89 ), .Y(\us33/n10 ) );
  OAI22X1 \us33/U233  ( .A0(\us33/n291 ), .A1(\us33/n114 ), .B0(\us33/n292 ), 
        .B1(\us33/n10 ), .Y(\us33/n286 ) );
  INVX1 \us33/U232  ( .A(\us33/n225 ), .Y(\us33/n288 ) );
  NAND2X1 \us33/U231  ( .A(\us33/n200 ), .B(\us33/n284 ), .Y(\us33/n102 ) );
  NOR2X1 \us33/U230  ( .A(\us33/n290 ), .B(\us33/n163 ), .Y(\us33/n184 ) );
  AOI22X1 \us33/U229  ( .A0(\us33/n102 ), .A1(\us33/n69 ), .B0(\us33/n184 ), 
        .B1(\us33/n33 ), .Y(\us33/n289 ) );
  AOI31X1 \us33/U228  ( .A0(\us33/n132 ), .A1(\us33/n288 ), .A2(\us33/n289 ), 
        .B0(\us33/n52 ), .Y(\us33/n287 ) );
  AOI211X1 \us33/U227  ( .A0(\us33/n285 ), .A1(\us33/n55 ), .B0(\us33/n286 ), 
        .C0(\us33/n287 ), .Y(\us33/n263 ) );
  NAND2X1 \us33/U226  ( .A(\us33/n284 ), .B(\us33/n122 ), .Y(\us33/n125 ) );
  NOR2X1 \us33/U225  ( .A(\us33/n199 ), .B(\us33/n4 ), .Y(\us33/n50 ) );
  AOI21X1 \us33/U224  ( .A0(\us33/n200 ), .A1(\us33/n223 ), .B0(\us33/n20 ), 
        .Y(\us33/n283 ) );
  AOI211X1 \us33/U223  ( .A0(\us33/n5 ), .A1(\us33/n125 ), .B0(\us33/n50 ), 
        .C0(\us33/n283 ), .Y(\us33/n282 ) );
  OAI221XL \us33/U222  ( .A0(\us33/n281 ), .A1(\us33/n27 ), .B0(\us33/n4 ), 
        .B1(\us33/n111 ), .C0(\us33/n282 ), .Y(\us33/n265 ) );
  INVX1 \us33/U221  ( .A(\us33/n280 ), .Y(\us33/n247 ) );
  NAND2X1 \us33/U220  ( .A(\us33/n41 ), .B(\us33/n33 ), .Y(\us33/n272 ) );
  OAI221XL \us33/U219  ( .A0(sa33[1]), .A1(\us33/n247 ), .B0(\us33/n4 ), .B1(
        \us33/n189 ), .C0(\us33/n272 ), .Y(\us33/n279 ) );
  NAND2X1 \us33/U218  ( .A(sa33[2]), .B(\us33/n149 ), .Y(\us33/n276 ) );
  XNOR2X1 \us33/U217  ( .A(\us33/n129 ), .B(sa33[1]), .Y(\us33/n155 ) );
  MXI2X1 \us33/U216  ( .A(\us33/n276 ), .B(\us33/n277 ), .S0(\us33/n155 ), .Y(
        \us33/n275 ) );
  OAI22X1 \us33/U215  ( .A0(\us33/n273 ), .A1(\us33/n10 ), .B0(\us33/n274 ), 
        .B1(\us33/n52 ), .Y(\us33/n266 ) );
  NOR2X1 \us33/U214  ( .A(\us33/n20 ), .B(\us33/n226 ), .Y(\us33/n176 ) );
  OAI21XL \us33/U213  ( .A0(\us33/n4 ), .A1(\us33/n271 ), .B0(\us33/n272 ), 
        .Y(\us33/n270 ) );
  OAI31X1 \us33/U212  ( .A0(\us33/n176 ), .A1(\us33/n269 ), .A2(\us33/n270 ), 
        .B0(\us33/n16 ), .Y(\us33/n268 ) );
  INVX1 \us33/U211  ( .A(\us33/n268 ), .Y(\us33/n267 ) );
  AOI211X1 \us33/U210  ( .A0(\us33/n55 ), .A1(\us33/n265 ), .B0(\us33/n266 ), 
        .C0(\us33/n267 ), .Y(\us33/n264 ) );
  MXI2X1 \us33/U209  ( .A(\us33/n263 ), .B(\us33/n264 ), .S0(sa33[6]), .Y(
        sa30_sr[2]) );
  NOR2X1 \us33/U208  ( .A(\us33/n94 ), .B(sa33[1]), .Y(\us33/n211 ) );
  INVX1 \us33/U207  ( .A(\us33/n262 ), .Y(\us33/n261 ) );
  AOI211X1 \us33/U206  ( .A0(\us33/n259 ), .A1(\us33/n24 ), .B0(\us33/n260 ), 
        .C0(\us33/n261 ), .Y(\us33/n255 ) );
  OAI22X1 \us33/U205  ( .A0(\us33/n20 ), .A1(\us33/n68 ), .B0(\us33/n27 ), 
        .B1(\us33/n37 ), .Y(\us33/n257 ) );
  NOR3X1 \us33/U204  ( .A(\us33/n257 ), .B(\us33/n258 ), .C(\us33/n50 ), .Y(
        \us33/n256 ) );
  MXI2X1 \us33/U203  ( .A(\us33/n255 ), .B(\us33/n256 ), .S0(\us33/n252 ), .Y(
        \us33/n254 ) );
  AOI221X1 \us33/U202  ( .A0(\us33/n211 ), .A1(\us33/n5 ), .B0(\us33/n40 ), 
        .B1(sa33[4]), .C0(\us33/n254 ), .Y(\us33/n248 ) );
  INVX1 \us33/U201  ( .A(\us33/n211 ), .Y(\us33/n106 ) );
  NAND2X1 \us33/U200  ( .A(\us33/n200 ), .B(\us33/n106 ), .Y(\us33/n83 ) );
  NAND2X1 \us33/U199  ( .A(\us33/n199 ), .B(\us33/n204 ), .Y(\us33/n169 ) );
  AOI2BB2X1 \us33/U198  ( .B0(\us33/n65 ), .B1(\us33/n24 ), .A0N(\us33/n169 ), 
        .A1N(\us33/n20 ), .Y(\us33/n253 ) );
  OAI221XL \us33/U197  ( .A0(\us33/n172 ), .A1(\us33/n18 ), .B0(\us33/n27 ), 
        .B1(\us33/n83 ), .C0(\us33/n253 ), .Y(\us33/n251 ) );
  MXI2X1 \us33/U196  ( .A(\us33/n250 ), .B(\us33/n251 ), .S0(\us33/n252 ), .Y(
        \us33/n249 ) );
  MXI2X1 \us33/U195  ( .A(\us33/n248 ), .B(\us33/n249 ), .S0(\us33/n234 ), .Y(
        \us33/n228 ) );
  OAI21XL \us33/U194  ( .A0(\us33/n58 ), .A1(\us33/n27 ), .B0(\us33/n247 ), 
        .Y(\us33/n245 ) );
  NOR2X1 \us33/U193  ( .A(sa33[7]), .B(\us33/n145 ), .Y(\us33/n246 ) );
  XNOR2X1 \us33/U192  ( .A(\us33/n69 ), .B(sa33[1]), .Y(\us33/n130 ) );
  MXI2X1 \us33/U191  ( .A(\us33/n245 ), .B(\us33/n246 ), .S0(\us33/n130 ), .Y(
        \us33/n243 ) );
  OAI211X1 \us33/U190  ( .A0(\us33/n4 ), .A1(\us33/n149 ), .B0(\us33/n243 ), 
        .C0(\us33/n244 ), .Y(\us33/n230 ) );
  NOR2X1 \us33/U189  ( .A(\us33/n242 ), .B(\us33/n137 ), .Y(\us33/n70 ) );
  OAI221XL \us33/U188  ( .A0(\us33/n159 ), .A1(\us33/n27 ), .B0(\us33/n20 ), 
        .B1(\us33/n34 ), .C0(\us33/n241 ), .Y(\us33/n231 ) );
  NAND2X1 \us33/U187  ( .A(\us33/n101 ), .B(\us33/n240 ), .Y(\us33/n76 ) );
  AOI21X1 \us33/U186  ( .A0(\us33/n122 ), .A1(\us33/n106 ), .B0(\us33/n129 ), 
        .Y(\us33/n237 ) );
  INVX1 \us33/U185  ( .A(\us33/n239 ), .Y(\us33/n238 ) );
  OAI21XL \us33/U184  ( .A0(\us33/n237 ), .A1(\us33/n43 ), .B0(\us33/n238 ), 
        .Y(\us33/n236 ) );
  OAI221XL \us33/U183  ( .A0(\us33/n18 ), .A1(\us33/n76 ), .B0(\us33/n59 ), 
        .B1(\us33/n27 ), .C0(\us33/n236 ), .Y(\us33/n232 ) );
  AOI2BB2X1 \us33/U182  ( .B0(\us33/n24 ), .B1(\us33/n187 ), .A0N(\us33/n227 ), 
        .A1N(\us33/n20 ), .Y(\us33/n235 ) );
  OAI211X1 \us33/U181  ( .A0(\us33/n27 ), .A1(\us33/n122 ), .B0(\us33/n158 ), 
        .C0(\us33/n235 ), .Y(\us33/n233 ) );
  MX4X1 \us33/U180  ( .A(\us33/n230 ), .B(\us33/n231 ), .C(\us33/n232 ), .D(
        \us33/n233 ), .S0(\us33/n234 ), .S1(sa33[5]), .Y(\us33/n229 ) );
  MX2X1 \us33/U179  ( .A(\us33/n228 ), .B(\us33/n229 ), .S0(sa33[6]), .Y(
        sa30_sr[3]) );
  NOR2BX1 \us33/U178  ( .AN(\us33/n204 ), .B(\us33/n137 ), .Y(\us33/n110 ) );
  INVX1 \us33/U177  ( .A(\us33/n110 ), .Y(\us33/n64 ) );
  AOI22X1 \us33/U176  ( .A0(\us33/n225 ), .A1(\us33/n226 ), .B0(\us33/n6 ), 
        .B1(\us33/n227 ), .Y(\us33/n224 ) );
  OAI221XL \us33/U175  ( .A0(\us33/n27 ), .A1(\us33/n64 ), .B0(\us33/n4 ), 
        .B1(\us33/n83 ), .C0(\us33/n224 ), .Y(\us33/n212 ) );
  NAND2X1 \us33/U174  ( .A(\us33/n34 ), .B(\us33/n204 ), .Y(\us33/n221 ) );
  OAI21XL \us33/U173  ( .A0(\us33/n69 ), .A1(\us33/n223 ), .B0(\us33/n27 ), 
        .Y(\us33/n222 ) );
  NOR2X1 \us33/U172  ( .A(\us33/n217 ), .B(\us33/n42 ), .Y(\us33/n208 ) );
  AOI211X1 \us33/U171  ( .A0(\us33/n208 ), .A1(\us33/n5 ), .B0(\us33/n220 ), 
        .C0(\us33/n173 ), .Y(\us33/n219 ) );
  OAI22X1 \us33/U170  ( .A0(\us33/n218 ), .A1(\us33/n10 ), .B0(\us33/n219 ), 
        .B1(\us33/n114 ), .Y(\us33/n213 ) );
  INVX1 \us33/U169  ( .A(\us33/n135 ), .Y(\us33/n215 ) );
  NOR2X1 \us33/U168  ( .A(\us33/n4 ), .B(\us33/n159 ), .Y(\us33/n31 ) );
  INVX1 \us33/U167  ( .A(\us33/n31 ), .Y(\us33/n196 ) );
  AOI31X1 \us33/U166  ( .A0(\us33/n215 ), .A1(\us33/n196 ), .A2(\us33/n216 ), 
        .B0(\us33/n52 ), .Y(\us33/n214 ) );
  AOI211X1 \us33/U165  ( .A0(\us33/n55 ), .A1(\us33/n212 ), .B0(\us33/n213 ), 
        .C0(\us33/n214 ), .Y(\us33/n190 ) );
  INVX1 \us33/U164  ( .A(\us33/n207 ), .Y(\us33/n192 ) );
  NOR2X1 \us33/U163  ( .A(\us33/n25 ), .B(\us33/n98 ), .Y(\us33/n32 ) );
  OAI22X1 \us33/U162  ( .A0(\us33/n28 ), .A1(\us33/n4 ), .B0(\us33/n188 ), 
        .B1(\us33/n27 ), .Y(\us33/n206 ) );
  NAND2X1 \us33/U161  ( .A(\us33/n204 ), .B(\us33/n80 ), .Y(\us33/n118 ) );
  INVX1 \us33/U160  ( .A(\us33/n118 ), .Y(\us33/n123 ) );
  NAND2X1 \us33/U159  ( .A(\us33/n94 ), .B(\us33/n79 ), .Y(\us33/n203 ) );
  OAI2BB1X1 \us33/U158  ( .A0N(\us33/n199 ), .A1N(\us33/n200 ), .B0(\us33/n33 ), .Y(\us33/n195 ) );
  INVX1 \us33/U157  ( .A(\us33/n55 ), .Y(\us33/n12 ) );
  AOI31X1 \us33/U156  ( .A0(\us33/n195 ), .A1(\us33/n196 ), .A2(\us33/n197 ), 
        .B0(\us33/n12 ), .Y(\us33/n194 ) );
  AOI211X1 \us33/U155  ( .A0(\us33/n89 ), .A1(\us33/n192 ), .B0(\us33/n193 ), 
        .C0(\us33/n194 ), .Y(\us33/n191 ) );
  MXI2X1 \us33/U154  ( .A(\us33/n190 ), .B(\us33/n191 ), .S0(sa33[6]), .Y(
        sa30_sr[4]) );
  OAI21XL \us33/U153  ( .A0(\us33/n69 ), .A1(\us33/n189 ), .B0(\us33/n27 ), 
        .Y(\us33/n186 ) );
  INVX1 \us33/U152  ( .A(\us33/n183 ), .Y(\us33/n180 ) );
  NAND2X1 \us33/U151  ( .A(\us33/n74 ), .B(\us33/n182 ), .Y(\us33/n181 ) );
  AOI211X1 \us33/U150  ( .A0(\us33/n179 ), .A1(\us33/n24 ), .B0(\us33/n180 ), 
        .C0(\us33/n181 ), .Y(\us33/n165 ) );
  INVX1 \us33/U149  ( .A(\us33/n178 ), .Y(\us33/n175 ) );
  AOI211X1 \us33/U148  ( .A0(\us33/n175 ), .A1(\us33/n5 ), .B0(\us33/n176 ), 
        .C0(\us33/n177 ), .Y(\us33/n174 ) );
  OAI221XL \us33/U147  ( .A0(\us33/n159 ), .A1(\us33/n27 ), .B0(\us33/n145 ), 
        .B1(\us33/n20 ), .C0(\us33/n174 ), .Y(\us33/n167 ) );
  MXI2X1 \us33/U146  ( .A(\us33/n40 ), .B(\us33/n173 ), .S0(\us33/n96 ), .Y(
        \us33/n170 ) );
  AOI22X1 \us33/U145  ( .A0(\us33/n137 ), .A1(\us33/n24 ), .B0(\us33/n172 ), 
        .B1(\us33/n6 ), .Y(\us33/n171 ) );
  OAI211X1 \us33/U144  ( .A0(\us33/n20 ), .A1(\us33/n169 ), .B0(\us33/n170 ), 
        .C0(\us33/n171 ), .Y(\us33/n168 ) );
  AOI22X1 \us33/U143  ( .A0(\us33/n89 ), .A1(\us33/n167 ), .B0(\us33/n55 ), 
        .B1(\us33/n168 ), .Y(\us33/n166 ) );
  OAI221XL \us33/U142  ( .A0(\us33/n164 ), .A1(\us33/n114 ), .B0(\us33/n165 ), 
        .B1(\us33/n52 ), .C0(\us33/n166 ), .Y(\us33/n138 ) );
  OAI21XL \us33/U141  ( .A0(\us33/n41 ), .A1(\us33/n163 ), .B0(\us33/n69 ), 
        .Y(\us33/n162 ) );
  AOI221X1 \us33/U140  ( .A0(\us33/n159 ), .A1(\us33/n24 ), .B0(\us33/n160 ), 
        .B1(\us33/n33 ), .C0(\us33/n161 ), .Y(\us33/n140 ) );
  OAI21XL \us33/U139  ( .A0(\us33/n157 ), .A1(\us33/n20 ), .B0(\us33/n158 ), 
        .Y(\us33/n156 ) );
  NOR2X1 \us33/U138  ( .A(\us33/n4 ), .B(\us33/n136 ), .Y(\us33/n153 ) );
  NOR2X1 \us33/U137  ( .A(\us33/n145 ), .B(\us33/n69 ), .Y(\us33/n154 ) );
  MXI2X1 \us33/U136  ( .A(\us33/n153 ), .B(\us33/n154 ), .S0(\us33/n155 ), .Y(
        \us33/n152 ) );
  OAI221XL \us33/U135  ( .A0(\us33/n110 ), .A1(\us33/n18 ), .B0(\us33/n20 ), 
        .B1(\us33/n151 ), .C0(\us33/n152 ), .Y(\us33/n143 ) );
  AOI21X1 \us33/U134  ( .A0(\us33/n149 ), .A1(\us33/n150 ), .B0(\us33/n18 ), 
        .Y(\us33/n148 ) );
  AOI2BB1X1 \us33/U133  ( .A0N(\us33/n147 ), .A1N(\us33/n27 ), .B0(\us33/n148 ), .Y(\us33/n146 ) );
  OAI221XL \us33/U132  ( .A0(\us33/n145 ), .A1(\us33/n20 ), .B0(\us33/n4 ), 
        .B1(\us33/n34 ), .C0(\us33/n146 ), .Y(\us33/n144 ) );
  AOI22X1 \us33/U131  ( .A0(\us33/n89 ), .A1(\us33/n143 ), .B0(\us33/n14 ), 
        .B1(\us33/n144 ), .Y(\us33/n142 ) );
  OAI221XL \us33/U130  ( .A0(\us33/n140 ), .A1(\us33/n12 ), .B0(\us33/n141 ), 
        .B1(\us33/n114 ), .C0(\us33/n142 ), .Y(\us33/n139 ) );
  MX2X1 \us33/U129  ( .A(\us33/n138 ), .B(\us33/n139 ), .S0(sa33[6]), .Y(
        sa30_sr[5]) );
  INVX1 \us33/U128  ( .A(\us33/n70 ), .Y(\us33/n133 ) );
  OAI22X1 \us33/U127  ( .A0(\us33/n4 ), .A1(\us33/n136 ), .B0(\us33/n137 ), 
        .B1(\us33/n27 ), .Y(\us33/n134 ) );
  AOI211X1 \us33/U126  ( .A0(\us33/n133 ), .A1(\us33/n69 ), .B0(\us33/n134 ), 
        .C0(\us33/n135 ), .Y(\us33/n112 ) );
  INVX1 \us33/U125  ( .A(\us33/n132 ), .Y(\us33/n131 ) );
  OAI21XL \us33/U124  ( .A0(\us33/n18 ), .A1(\us33/n37 ), .B0(\us33/n128 ), 
        .Y(\us33/n127 ) );
  OAI221XL \us33/U123  ( .A0(\us33/n18 ), .A1(\us33/n105 ), .B0(\us33/n123 ), 
        .B1(\us33/n27 ), .C0(\us33/n124 ), .Y(\us33/n116 ) );
  NAND2X1 \us33/U122  ( .A(\us33/n121 ), .B(\us33/n122 ), .Y(\us33/n30 ) );
  OAI221XL \us33/U121  ( .A0(\us33/n18 ), .A1(\us33/n118 ), .B0(\us33/n27 ), 
        .B1(\us33/n30 ), .C0(\us33/n119 ), .Y(\us33/n117 ) );
  AOI22X1 \us33/U120  ( .A0(\us33/n89 ), .A1(\us33/n116 ), .B0(\us33/n55 ), 
        .B1(\us33/n117 ), .Y(\us33/n115 ) );
  OAI221XL \us33/U119  ( .A0(\us33/n112 ), .A1(\us33/n52 ), .B0(\us33/n113 ), 
        .B1(\us33/n114 ), .C0(\us33/n115 ), .Y(\us33/n84 ) );
  OAI22X1 \us33/U118  ( .A0(\us33/n110 ), .A1(\us33/n4 ), .B0(\us33/n20 ), 
        .B1(\us33/n21 ), .Y(\us33/n108 ) );
  AOI21X1 \us33/U117  ( .A0(sa33[1]), .A1(\us33/n58 ), .B0(\us33/n27 ), .Y(
        \us33/n109 ) );
  AOI211X1 \us33/U116  ( .A0(\us33/n5 ), .A1(\us33/n107 ), .B0(\us33/n108 ), 
        .C0(\us33/n109 ), .Y(\us33/n86 ) );
  OAI22X1 \us33/U115  ( .A0(\us33/n45 ), .A1(\us33/n4 ), .B0(sa33[4]), .B1(
        \us33/n18 ), .Y(\us33/n103 ) );
  AOI21X1 \us33/U114  ( .A0(\us33/n105 ), .A1(\us33/n106 ), .B0(\us33/n20 ), 
        .Y(\us33/n104 ) );
  AOI211X1 \us33/U113  ( .A0(\us33/n33 ), .A1(\us33/n102 ), .B0(\us33/n103 ), 
        .C0(\us33/n104 ), .Y(\us33/n87 ) );
  NAND2X1 \us33/U112  ( .A(\us33/n100 ), .B(\us33/n101 ), .Y(\us33/n62 ) );
  OAI221XL \us33/U111  ( .A0(\us33/n27 ), .A1(\us33/n62 ), .B0(\us33/n4 ), 
        .B1(\us33/n21 ), .C0(\us33/n97 ), .Y(\us33/n90 ) );
  NOR3X1 \us33/U110  ( .A(\us33/n4 ), .B(\us33/n95 ), .C(\us33/n96 ), .Y(
        \us33/n67 ) );
  AOI31X1 \us33/U109  ( .A0(\us33/n79 ), .A1(\us33/n94 ), .A2(\us33/n6 ), .B0(
        \us33/n67 ), .Y(\us33/n93 ) );
  OAI221XL \us33/U108  ( .A0(\us33/n73 ), .A1(\us33/n27 ), .B0(\us33/n92 ), 
        .B1(\us33/n20 ), .C0(\us33/n93 ), .Y(\us33/n91 ) );
  AOI22X1 \us33/U107  ( .A0(\us33/n89 ), .A1(\us33/n90 ), .B0(\us33/n16 ), 
        .B1(\us33/n91 ), .Y(\us33/n88 ) );
  OAI221XL \us33/U106  ( .A0(\us33/n86 ), .A1(\us33/n52 ), .B0(\us33/n87 ), 
        .B1(\us33/n12 ), .C0(\us33/n88 ), .Y(\us33/n85 ) );
  MX2X1 \us33/U105  ( .A(\us33/n84 ), .B(\us33/n85 ), .S0(sa33[6]), .Y(
        sa30_sr[6]) );
  INVX1 \us33/U104  ( .A(\us33/n81 ), .Y(\us33/n77 ) );
  AOI21X1 \us33/U103  ( .A0(\us33/n79 ), .A1(\us33/n80 ), .B0(\us33/n27 ), .Y(
        \us33/n78 ) );
  AOI211X1 \us33/U102  ( .A0(\us33/n5 ), .A1(\us33/n76 ), .B0(\us33/n77 ), 
        .C0(\us33/n78 ), .Y(\us33/n51 ) );
  OAI211X1 \us33/U101  ( .A0(\us33/n73 ), .A1(\us33/n27 ), .B0(\us33/n74 ), 
        .C0(\us33/n75 ), .Y(\us33/n72 ) );
  AOI21X1 \us33/U100  ( .A0(\us33/n68 ), .A1(\us33/n69 ), .B0(\us33/n6 ), .Y(
        \us33/n63 ) );
  INVX1 \us33/U99  ( .A(\us33/n67 ), .Y(\us33/n66 ) );
  OAI221XL \us33/U98  ( .A0(\us33/n63 ), .A1(\us33/n64 ), .B0(\us33/n65 ), 
        .B1(\us33/n27 ), .C0(\us33/n66 ), .Y(\us33/n56 ) );
  AOI2BB2X1 \us33/U97  ( .B0(\us33/n61 ), .B1(\us33/n24 ), .A0N(\us33/n62 ), 
        .A1N(\us33/n20 ), .Y(\us33/n60 ) );
  OAI221XL \us33/U96  ( .A0(\us33/n58 ), .A1(\us33/n18 ), .B0(\us33/n59 ), 
        .B1(\us33/n27 ), .C0(\us33/n60 ), .Y(\us33/n57 ) );
  AOI22X1 \us33/U95  ( .A0(\us33/n55 ), .A1(\us33/n56 ), .B0(\us33/n16 ), .B1(
        \us33/n57 ), .Y(\us33/n54 ) );
  OAI221XL \us33/U94  ( .A0(\us33/n51 ), .A1(\us33/n52 ), .B0(\us33/n53 ), 
        .B1(\us33/n10 ), .C0(\us33/n54 ), .Y(\us33/n7 ) );
  INVX1 \us33/U93  ( .A(\us33/n50 ), .Y(\us33/n49 ) );
  OAI221XL \us33/U92  ( .A0(\us33/n47 ), .A1(\us33/n18 ), .B0(\us33/n27 ), 
        .B1(\us33/n48 ), .C0(\us33/n49 ), .Y(\us33/n46 ) );
  NOR2X1 \us33/U91  ( .A(\us33/n41 ), .B(\us33/n42 ), .Y(\us33/n38 ) );
  INVX1 \us33/U90  ( .A(\us33/n40 ), .Y(\us33/n39 ) );
  INVX1 \us33/U89  ( .A(\us33/n32 ), .Y(\us33/n26 ) );
  AOI21X1 \us33/U88  ( .A0(\us33/n5 ), .A1(\us33/n30 ), .B0(\us33/n31 ), .Y(
        \us33/n29 ) );
  OAI221XL \us33/U87  ( .A0(\us33/n26 ), .A1(\us33/n27 ), .B0(\us33/n28 ), 
        .B1(\us33/n20 ), .C0(\us33/n29 ), .Y(\us33/n15 ) );
  OAI221XL \us33/U86  ( .A0(\us33/n18 ), .A1(\us33/n19 ), .B0(\us33/n20 ), 
        .B1(\us33/n21 ), .C0(\us33/n22 ), .Y(\us33/n17 ) );
  AOI22X1 \us33/U85  ( .A0(\us33/n14 ), .A1(\us33/n15 ), .B0(\us33/n16 ), .B1(
        \us33/n17 ), .Y(\us33/n13 ) );
  OAI221XL \us33/U84  ( .A0(\us33/n9 ), .A1(\us33/n10 ), .B0(\us33/n11 ), .B1(
        \us33/n12 ), .C0(\us33/n13 ), .Y(\us33/n8 ) );
  MX2X1 \us33/U83  ( .A(\us33/n7 ), .B(\us33/n8 ), .S0(sa33[6]), .Y(sa30_sr[7]) );
  NOR2X4 \us33/U82  ( .A(\us33/n129 ), .B(sa33[2]), .Y(\us33/n43 ) );
  CLKINVX3 \us33/U81  ( .A(\us33/n14 ), .Y(\us33/n52 ) );
  OAI22XL \us33/U80  ( .A0(\us33/n201 ), .A1(\us33/n52 ), .B0(\us33/n202 ), 
        .B1(\us33/n114 ), .Y(\us33/n193 ) );
  CLKINVX3 \us33/U79  ( .A(sa33[5]), .Y(\us33/n252 ) );
  NOR2X2 \us33/U78  ( .A(\us33/n252 ), .B(\us33/n234 ), .Y(\us33/n55 ) );
  CLKINVX3 \us33/U77  ( .A(sa33[7]), .Y(\us33/n129 ) );
  NOR2X4 \us33/U76  ( .A(\us33/n129 ), .B(\us33/n69 ), .Y(\us33/n24 ) );
  AOI22XL \us33/U75  ( .A0(\us33/n70 ), .A1(\us33/n24 ), .B0(\us33/n96 ), .B1(
        \us33/n129 ), .Y(\us33/n241 ) );
  NOR2X2 \us33/U74  ( .A(\us33/n252 ), .B(sa33[0]), .Y(\us33/n89 ) );
  CLKINVX3 \us33/U73  ( .A(sa33[0]), .Y(\us33/n234 ) );
  NOR2X4 \us33/U72  ( .A(\us33/n69 ), .B(sa33[7]), .Y(\us33/n33 ) );
  INVX12 \us33/U71  ( .A(\us33/n33 ), .Y(\us33/n27 ) );
  CLKINVX3 \us33/U70  ( .A(\us33/n1 ), .Y(\us33/n6 ) );
  CLKINVX3 \us33/U69  ( .A(\us33/n1 ), .Y(\us33/n5 ) );
  INVXL \us33/U68  ( .A(\us33/n24 ), .Y(\us33/n36 ) );
  INVX4 \us33/U67  ( .A(\us33/n3 ), .Y(\us33/n4 ) );
  INVXL \us33/U66  ( .A(\us33/n36 ), .Y(\us33/n3 ) );
  INVX4 \us33/U65  ( .A(sa33[1]), .Y(\us33/n226 ) );
  INVX4 \us33/U64  ( .A(\us33/n43 ), .Y(\us33/n20 ) );
  AOI221X4 \us33/U63  ( .A0(\us33/n24 ), .A1(\us33/n82 ), .B0(\us33/n43 ), 
        .B1(\us33/n295 ), .C0(\us33/n173 ), .Y(\us33/n346 ) );
  AOI221X4 \us33/U62  ( .A0(\us33/n5 ), .A1(\us33/n96 ), .B0(\us33/n43 ), .B1(
        \us33/n239 ), .C0(\us33/n340 ), .Y(\us33/n336 ) );
  AOI222X4 \us33/U61  ( .A0(\us33/n59 ), .A1(\us33/n43 ), .B0(\us33/n6 ), .B1(
        \us33/n221 ), .C0(\us33/n222 ), .C1(\us33/n187 ), .Y(\us33/n218 ) );
  AOI222X4 \us33/U60  ( .A0(\us33/n123 ), .A1(\us33/n43 ), .B0(sa33[2]), .B1(
        \us33/n203 ), .C0(\us33/n6 ), .C1(\us33/n71 ), .Y(\us33/n202 ) );
  AOI221X4 \us33/U59  ( .A0(\us33/n314 ), .A1(\us33/n43 ), .B0(\us33/n160 ), 
        .B1(\us33/n24 ), .C0(\us33/n315 ), .Y(\us33/n307 ) );
  AOI221X4 \us33/U58  ( .A0(\us33/n43 ), .A1(\us33/n208 ), .B0(\us33/n76 ), 
        .B1(\us33/n24 ), .C0(\us33/n209 ), .Y(\us33/n207 ) );
  AOI221X4 \us33/U57  ( .A0(\us33/n43 ), .A1(\us33/n205 ), .B0(\us33/n32 ), 
        .B1(\us33/n6 ), .C0(\us33/n206 ), .Y(\us33/n201 ) );
  AOI221X4 \us33/U56  ( .A0(\us33/n43 ), .A1(\us33/n44 ), .B0(\us33/n45 ), 
        .B1(\us33/n24 ), .C0(\us33/n46 ), .Y(\us33/n9 ) );
  AOI22XL \us33/U55  ( .A0(\us33/n217 ), .A1(\us33/n43 ), .B0(\us33/n33 ), 
        .B1(\us33/n47 ), .Y(\us33/n216 ) );
  AOI22XL \us33/U54  ( .A0(\us33/n98 ), .A1(\us33/n43 ), .B0(\us33/n6 ), .B1(
        \us33/n99 ), .Y(\us33/n97 ) );
  AOI22XL \us33/U53  ( .A0(\us33/n82 ), .A1(\us33/n43 ), .B0(\us33/n83 ), .B1(
        \us33/n24 ), .Y(\us33/n81 ) );
  AOI2BB2XL \us33/U52  ( .B0(\us33/n43 ), .B1(\us33/n94 ), .A0N(\us33/n120 ), 
        .A1N(\us33/n4 ), .Y(\us33/n119 ) );
  AOI222X4 \us33/U51  ( .A0(\us33/n125 ), .A1(\us33/n33 ), .B0(\us33/n145 ), 
        .B1(\us33/n40 ), .C0(\us33/n43 ), .C1(\us33/n184 ), .Y(\us33/n183 ) );
  AOI22XL \us33/U50  ( .A0(\us33/n43 ), .A1(\us33/n303 ), .B0(\us33/n24 ), 
        .B1(\us33/n96 ), .Y(\us33/n358 ) );
  AOI22XL \us33/U49  ( .A0(\us33/n43 ), .A1(\us33/n100 ), .B0(\us33/n24 ), 
        .B1(\us33/n125 ), .Y(\us33/n124 ) );
  AOI21XL \us33/U48  ( .A0(\us33/n159 ), .A1(\us33/n43 ), .B0(\us33/n40 ), .Y(
        \us33/n262 ) );
  AOI22XL \us33/U47  ( .A0(\us33/n40 ), .A1(\us33/n94 ), .B0(\us33/n43 ), .B1(
        \us33/n187 ), .Y(\us33/n244 ) );
  AOI22XL \us33/U46  ( .A0(\us33/n184 ), .A1(\us33/n5 ), .B0(\us33/n198 ), 
        .B1(\us33/n43 ), .Y(\us33/n197 ) );
  NOR2XL \us33/U45  ( .A(\us33/n33 ), .B(\us33/n2 ), .Y(\us33/n302 ) );
  MXI2XL \us33/U44  ( .A(\us33/n2 ), .B(\us33/n6 ), .S0(\us33/n28 ), .Y(
        \us33/n311 ) );
  INVXL \us33/U43  ( .A(\us33/n20 ), .Y(\us33/n2 ) );
  INVX4 \us33/U42  ( .A(\us33/n6 ), .Y(\us33/n18 ) );
  AOI21XL \us33/U41  ( .A0(\us33/n18 ), .A1(\us33/n162 ), .B0(\us33/n25 ), .Y(
        \us33/n161 ) );
  INVX4 \us33/U40  ( .A(sa33[2]), .Y(\us33/n69 ) );
  NOR2X4 \us33/U39  ( .A(\us33/n226 ), .B(\us33/n4 ), .Y(\us33/n40 ) );
  CLKINVX3 \us33/U38  ( .A(sa33[3]), .Y(\us33/n136 ) );
  NOR2X2 \us33/U37  ( .A(\us33/n136 ), .B(sa33[4]), .Y(\us33/n145 ) );
  CLKINVX3 \us33/U36  ( .A(sa33[4]), .Y(\us33/n58 ) );
  NOR2X2 \us33/U35  ( .A(\us33/n58 ), .B(sa33[3]), .Y(\us33/n159 ) );
  NOR2X2 \us33/U34  ( .A(\us33/n136 ), .B(\us33/n58 ), .Y(\us33/n259 ) );
  NOR2X2 \us33/U33  ( .A(sa33[4]), .B(sa33[3]), .Y(\us33/n278 ) );
  NOR2X2 \us33/U32  ( .A(\us33/n259 ), .B(\us33/n278 ), .Y(\us33/n47 ) );
  CLKINVX3 \us33/U31  ( .A(\us33/n259 ), .Y(\us33/n44 ) );
  NOR2X2 \us33/U30  ( .A(\us33/n44 ), .B(sa33[1]), .Y(\us33/n137 ) );
  AOI21XL \us33/U29  ( .A0(\us33/n44 ), .A1(\us33/n111 ), .B0(\us33/n4 ), .Y(
        \us33/n177 ) );
  AOI22XL \us33/U28  ( .A0(\us33/n23 ), .A1(\us33/n24 ), .B0(\us33/n25 ), .B1(
        sa33[2]), .Y(\us33/n22 ) );
  AOI22XL \us33/U27  ( .A0(\us33/n33 ), .A1(sa33[3]), .B0(\us33/n24 ), .B1(
        \us33/n58 ), .Y(\us33/n277 ) );
  NAND2XL \us33/U26  ( .A(\us33/n198 ), .B(\us33/n24 ), .Y(\us33/n132 ) );
  OAI2BB2XL \us33/U25  ( .B0(\us33/n20 ), .B1(\us33/n111 ), .A0N(\us33/n125 ), 
        .A1N(\us33/n24 ), .Y(\us33/n220 ) );
  NAND2XL \us33/U24  ( .A(\us33/n111 ), .B(\us33/n101 ), .Y(\us33/n21 ) );
  NAND2XL \us33/U23  ( .A(\us33/n111 ), .B(\us33/n300 ), .Y(\us33/n187 ) );
  NAND2XL \us33/U22  ( .A(\us33/n111 ), .B(\us33/n121 ), .Y(\us33/n303 ) );
  AOI221XL \us33/U21  ( .A0(\us33/n43 ), .A1(\us33/n151 ), .B0(\us33/n25 ), 
        .B1(\us33/n69 ), .C0(\us33/n275 ), .Y(\us33/n274 ) );
  NOR2BXL \us33/U20  ( .AN(\us33/n101 ), .B(\us33/n25 ), .Y(\us33/n172 ) );
  NAND2X2 \us33/U19  ( .A(\us33/n58 ), .B(\us33/n226 ), .Y(\us33/n34 ) );
  OAI222X1 \us33/U18  ( .A0(\us33/n27 ), .A1(\us33/n34 ), .B0(\us33/n69 ), 
        .B1(\us33/n205 ), .C0(\us33/n20 ), .C1(\us33/n79 ), .Y(\us33/n260 ) );
  OAI222X1 \us33/U17  ( .A0(\us33/n20 ), .A1(\us33/n99 ), .B0(\us33/n27 ), 
        .B1(\us33/n101 ), .C0(\us33/n184 ), .C1(\us33/n4 ), .Y(\us33/n250 ) );
  OAI222X1 \us33/U16  ( .A0(\us33/n4 ), .A1(\us33/n37 ), .B0(\us33/n38 ), .B1(
        \us33/n20 ), .C0(sa33[4]), .C1(\us33/n39 ), .Y(\us33/n35 ) );
  AOI221X1 \us33/U15  ( .A0(\us33/n5 ), .A1(\us33/n19 ), .B0(\us33/n33 ), .B1(
        \us33/n34 ), .C0(\us33/n35 ), .Y(\us33/n11 ) );
  OR2X2 \us33/U14  ( .A(sa33[2]), .B(sa33[7]), .Y(\us33/n1 ) );
  AOI221XL \us33/U13  ( .A0(\us33/n70 ), .A1(\us33/n43 ), .B0(\us33/n24 ), 
        .B1(\us33/n71 ), .C0(\us33/n72 ), .Y(\us33/n53 ) );
  AOI221XL \us33/U12  ( .A0(\us33/n59 ), .A1(\us33/n33 ), .B0(\us33/n43 ), 
        .B1(\us33/n126 ), .C0(\us33/n127 ), .Y(\us33/n113 ) );
  AOI222XL \us33/U11  ( .A0(\us33/n185 ), .A1(\us33/n43 ), .B0(\us33/n186 ), 
        .B1(\us33/n187 ), .C0(\us33/n6 ), .C1(\us33/n188 ), .Y(\us33/n164 ) );
  AOI221X1 \us33/U10  ( .A0(\us33/n313 ), .A1(\us33/n5 ), .B0(\us33/n23 ), 
        .B1(\us33/n2 ), .C0(\us33/n328 ), .Y(\us33/n320 ) );
  AOI221X1 \us33/U9  ( .A0(\us33/n40 ), .A1(\us33/n136 ), .B0(\us33/n33 ), 
        .B1(\us33/n178 ), .C0(\us33/n338 ), .Y(\us33/n337 ) );
  AOI222XL \us33/U8  ( .A0(\us33/n278 ), .A1(\us33/n24 ), .B0(\us33/n42 ), 
        .B1(\us33/n33 ), .C0(\us33/n43 ), .C1(\us33/n136 ), .Y(\us33/n351 ) );
  AOI31X1 \us33/U7  ( .A0(sa33[2]), .A1(\us33/n58 ), .A2(sa33[1]), .B0(
        \us33/n40 ), .Y(\us33/n350 ) );
  AOI31X1 \us33/U6  ( .A0(\us33/n44 ), .A1(\us33/n129 ), .A2(\us33/n130 ), 
        .B0(\us33/n131 ), .Y(\us33/n128 ) );
  AOI221X1 \us33/U5  ( .A0(\us33/n40 ), .A1(\us33/n136 ), .B0(\us33/n33 ), 
        .B1(\us33/n47 ), .C0(\us33/n156 ), .Y(\us33/n141 ) );
  OAI32X1 \us33/U4  ( .A0(\us33/n18 ), .A1(sa33[1]), .A2(\us33/n159 ), .B0(
        sa33[4]), .B1(\us33/n182 ), .Y(\us33/n318 ) );
  OAI32X1 \us33/U3  ( .A0(\us33/n210 ), .A1(\us33/n145 ), .A2(\us33/n18 ), 
        .B0(\us33/n27 ), .B1(\us33/n211 ), .Y(\us33/n209 ) );
  AOI221X1 \us33/U2  ( .A0(\us33/n278 ), .A1(\us33/n40 ), .B0(\us33/n185 ), 
        .B1(\us33/n2 ), .C0(\us33/n279 ), .Y(\us33/n273 ) );
  AOI31XL \us33/U1  ( .A0(\us33/n79 ), .A1(\us33/n44 ), .A2(\us33/n2 ), .B0(
        \us33/n280 ), .Y(\us33/n339 ) );
endmodule

