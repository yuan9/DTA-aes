library verilog;
use verilog.vl_types.all;
entity PVSS2DGZ is
    port(
        VSSPST          : inout  vl_logic
    );
end PVSS2DGZ;
