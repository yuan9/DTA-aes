library verilog;
use verilog.vl_types.all;
entity PVSS3DGZ is
    port(
        VSS             : inout  vl_logic
    );
end PVSS3DGZ;
