library verilog;
use verilog.vl_types.all;
entity PVDD1DGZ is
    port(
        VDD             : inout  vl_logic
    );
end PVDD1DGZ;
