library verilog;
use verilog.vl_types.all;
entity and3_lib is
    port(
        in0             : in     vl_logic;
        in1             : in     vl_logic;
        in2             : in     vl_logic;
        \out\           : out    vl_logic
    );
end and3_lib;
