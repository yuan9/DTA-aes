library verilog;
use verilog.vl_types.all;
entity PVDD1ANA is
    port(
        AVDD            : inout  vl_logic
    );
end PVDD1ANA;
