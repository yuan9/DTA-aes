library verilog;
use verilog.vl_types.all;
entity PDISDGZ is
    port(
        PAD             : in     vl_logic;
        C               : out    vl_logic
    );
end PDISDGZ;
