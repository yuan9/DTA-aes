library verilog;
use verilog.vl_types.all;
entity BUFXL is
    port(
        Y               : out    vl_logic;
        A               : in     vl_logic
    );
end BUFXL;
