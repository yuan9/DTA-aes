library verilog;
use verilog.vl_types.all;
entity ANTENNA is
    port(
        A               : in     vl_logic
    );
end ANTENNA;
