library verilog;
use verilog.vl_types.all;
entity PRO24CDG is
    port(
        I               : in     vl_logic;
        PAD             : out    vl_logic
    );
end PRO24CDG;
