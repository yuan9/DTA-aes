module PDB1A (
	inout AIO
);

	assign AIO = 1'b1; // dummy logic for as a place-holder

endmodule
