library verilog;
use verilog.vl_types.all;
entity PRCUT is
end PRCUT;
