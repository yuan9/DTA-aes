library verilog;
use verilog.vl_types.all;
entity PVSS1ANA is
    port(
        AVSS            : inout  vl_logic
    );
end PVSS1ANA;
