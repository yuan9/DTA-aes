************************************************************************************
* TSMC Library/IP Product
* Filename: tcb018gbwp7t_270a.spi
* Technology: CL018
* Product Type: Standard Cell
* Product Name: tcb018gbwp7t
* Version: 270a
*************************************************************************************
**
*  STATEMENT OF USE
*
*  This information contains confidential and proprietary information of TSMC.
*  No part of this information may be reproduced, transmitted, transcribed,
*  stored in a retrieval system, or translated into any human or computer
*  language, in any form or by any means, electronic, mechanical, magnetic,
*  optical, chemical, manual, or otherwise, without the prior written permission
*  of TSMC.  This information was prepared for informational purpose and is for
*  use by TSMC's customers only.  TSMC reserves the right to make changes in the
*  information at any time and without notice.
*
**************************************************************************************
.global VDD VSS
.subckt AN2D0BWP7T A1 A2 Z VDD VSS 
M_u3-M_u2 Z net6 VSS VSS n w=0.5u l=0.18u
M_u2-M_u4 X_u2-net6 A2 VSS VSS n w=0.5u l=0.18u
M_u2-M_u3 net6 A1 X_u2-net6 VSS n w=0.5u l=0.18u
M_u3-M_u3 Z net6 VDD VDD p w=0.685u l=0.18u
M_u2-M_u2 net6 A2 VDD VDD p w=0.685u l=0.18u
M_u2-M_u1 net6 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt AN2D1BWP7T A1 A2 Z VDD VSS 
M_u3-M_u2 Z net6 VSS VSS n w=1u l=0.18u
M_u2-M_u4 X_u2-net6 A2 VSS VSS n w=0.5u l=0.18u
M_u2-M_u3 net6 A1 X_u2-net6 VSS n w=0.5u l=0.18u
M_u3-M_u3 Z net6 VDD VDD p w=1.37u l=0.18u
M_u2-M_u2 net6 A2 VDD VDD p w=0.685u l=0.18u
M_u2-M_u1 net6 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt AN2D2BWP7T A1 A2 Z VDD VSS 
M_u3-M_u2 Z net10 VSS VSS n w=2u l=0.18u
M_u2-M_u4 X_u2-net6 A2 VSS VSS n w=1u l=0.18u
M_u2-M_u3 net10 A1 X_u2-net6 VSS n w=1u l=0.18u
M_u3-M_u3 Z net10 VDD VDD p w=2.74u l=0.18u
M_u2-M_u2 net10 A2 VDD VDD p w=1.37u l=0.18u
M_u2-M_u1 net10 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AN2D4BWP7T A1 A2 Z VDD VSS 
M_u3_0-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_2-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_3-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u2_0-M_u4 X_u2_0-net6 A2 VSS VSS n w=1u l=0.18u
M_u2_0-M_u3 p0 A1 X_u2_0-net6 VSS n w=1u l=0.18u
M_u2_1-M_u4 X_u2_1-net6 A2 VSS VSS n w=1u l=0.18u
M_u2_1-M_u3 p0 A1 X_u2_1-net6 VSS n w=1u l=0.18u
M_u3_0-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_2-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_3-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u2_0-M_u2 p0 A2 VDD VDD p w=1.37u l=0.18u
M_u2_0-M_u1 p0 A1 VDD VDD p w=1.37u l=0.18u
M_u2_1-M_u2 p0 A2 VDD VDD p w=1.37u l=0.18u
M_u2_1-M_u1 p0 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AN2XD1BWP7T A1 A2 Z VDD VSS 
M_u3-M_u2 Z net6 VSS VSS n w=1u l=0.18u
M_u2-M_u4 X_u2-net6 A2 VSS VSS n w=1u l=0.18u
M_u2-M_u3 net6 A1 X_u2-net6 VSS n w=1u l=0.18u
M_u3-M_u3 Z net6 VDD VDD p w=1.37u l=0.18u
M_u2-M_u2 net6 A2 VDD VDD p w=1.37u l=0.18u
M_u2-M_u1 net6 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AN3D0BWP7T A1 A2 A3 Z VDD VSS 
M_u4-M_u4 net7 A1 X_u4-net10 VSS n w=0.5u l=0.18u
M_u4-M_u5 X_u4-net10 A2 X_u4-net13 VSS n w=0.5u l=0.18u
M_u4-M_u6 X_u4-net13 A3 VSS VSS n w=0.5u l=0.18u
M_u3-M_u2 Z net7 VSS VSS n w=0.5u l=0.18u
M_u4-M_u3 net7 A3 VDD VDD p w=0.685u l=0.18u
M_u4-M_u1 net7 A1 VDD VDD p w=0.685u l=0.18u
M_u4-M_u2 net7 A2 VDD VDD p w=0.685u l=0.18u
M_u3-M_u3 Z net7 VDD VDD p w=0.685u l=0.18u
.ends
.subckt AN3D1BWP7T A1 A2 A3 Z VDD VSS 
M_u4-M_u4 net7 A1 X_u4-net10 VSS n w=0.5u l=0.18u
M_u4-M_u5 X_u4-net10 A2 X_u4-net13 VSS n w=0.5u l=0.18u
M_u4-M_u6 X_u4-net13 A3 VSS VSS n w=0.5u l=0.18u
M_u3-M_u2 Z net7 VSS VSS n w=1u l=0.18u
M_u4-M_u3 net7 A3 VDD VDD p w=0.685u l=0.18u
M_u4-M_u1 net7 A1 VDD VDD p w=0.685u l=0.18u
M_u4-M_u2 net7 A2 VDD VDD p w=0.685u l=0.18u
M_u3-M_u3 Z net7 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AN3D2BWP7T A1 A2 A3 Z VDD VSS 
M_u4-M_u4 net15 A1 X_u4-net10 VSS n w=1u l=0.18u
M_u4-M_u5 X_u4-net10 A2 X_u4-net13 VSS n w=1u l=0.18u
M_u4-M_u6 X_u4-net13 A3 VSS VSS n w=1u l=0.18u
M_u3_0-M_u2 Z net15 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z net15 VSS VSS n w=1u l=0.18u
M_u4-M_u3 net15 A3 VDD VDD p w=1.37u l=0.18u
M_u4-M_u1 net15 A1 VDD VDD p w=1.37u l=0.18u
M_u4-M_u2 net15 A2 VDD VDD p w=1.37u l=0.18u
M_u3_0-M_u3 Z net15 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z net15 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AN3D4BWP7T A1 A2 A3 Z VDD VSS 
M_u4_0-M_u4 p0 A1 X_u4_0-net10 VSS n w=1u l=0.18u
M_u4_0-M_u5 X_u4_0-net10 A2 X_u4_0-net13 VSS n w=1u l=0.18u
M_u4_0-M_u6 X_u4_0-net13 A3 VSS VSS n w=1u l=0.18u
M_u4_1-M_u4 p0 A1 X_u4_1-net10 VSS n w=1u l=0.18u
M_u4_1-M_u5 X_u4_1-net10 A2 X_u4_1-net13 VSS n w=1u l=0.18u
M_u4_1-M_u6 X_u4_1-net13 A3 VSS VSS n w=1u l=0.18u
M_u3_0-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_2-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_3-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u4_0-M_u3 p0 A3 VDD VDD p w=1.37u l=0.18u
M_u4_0-M_u1 p0 A1 VDD VDD p w=1.37u l=0.18u
M_u4_0-M_u2 p0 A2 VDD VDD p w=1.37u l=0.18u
M_u4_1-M_u3 p0 A3 VDD VDD p w=1.37u l=0.18u
M_u4_1-M_u1 p0 A1 VDD VDD p w=1.37u l=0.18u
M_u4_1-M_u2 p0 A2 VDD VDD p w=1.37u l=0.18u
M_u3_0-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_2-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_3-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AN3XD1BWP7T A1 A2 A3 Z VDD VSS 
M_u4-M_u4 net7 A1 X_u4-net10 VSS n w=1u l=0.18u
M_u4-M_u5 X_u4-net10 A2 X_u4-net13 VSS n w=1u l=0.18u
M_u4-M_u6 X_u4-net13 A3 VSS VSS n w=1u l=0.18u
M_u3-M_u2 Z net7 VSS VSS n w=1u l=0.18u
M_u4-M_u3 net7 A3 VDD VDD p w=1.37u l=0.18u
M_u4-M_u1 net7 A1 VDD VDD p w=1.37u l=0.18u
M_u4-M_u2 net7 A2 VDD VDD p w=1.37u l=0.18u
M_u3-M_u3 Z net7 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AN4D0BWP7T A1 A2 A3 A4 Z VDD VSS 
M_u3-M_u2 Z net6 VSS VSS n w=0.5u l=0.18u
MU30-M_u5 net6 A1 XU30-net23 VSS n w=0.5u l=0.18u
MU30-M_u6 XU30-net23 A2 XU30-net26 VSS n w=0.5u l=0.18u
MU30-M_u7 XU30-net26 A3 XU30-net29 VSS n w=0.5u l=0.18u
MU30-M_u8 XU30-net29 A4 VSS VSS n w=0.5u l=0.18u
M_u3-M_u3 Z net6 VDD VDD p w=0.685u l=0.18u
MU30-M_u4 net6 A4 VDD VDD p w=0.685u l=0.18u
MU30-M_u3 net6 A3 VDD VDD p w=0.685u l=0.18u
MU30-M_u2 net6 A2 VDD VDD p w=0.685u l=0.18u
MU30-M_u1 net6 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt AN4D1BWP7T A1 A2 A3 A4 Z VDD VSS 
M_u3-M_u2 Z net6 VSS VSS n w=1u l=0.18u
MU30-M_u5 net6 A1 XU30-net23 VSS n w=0.5u l=0.18u
MU30-M_u6 XU30-net23 A2 XU30-net26 VSS n w=0.5u l=0.18u
MU30-M_u7 XU30-net26 A3 XU30-net29 VSS n w=0.5u l=0.18u
MU30-M_u8 XU30-net29 A4 VSS VSS n w=0.5u l=0.18u
M_u3-M_u3 Z net6 VDD VDD p w=1.37u l=0.18u
MU30-M_u4 net6 A4 VDD VDD p w=0.685u l=0.18u
MU30-M_u3 net6 A3 VDD VDD p w=0.685u l=0.18u
MU30-M_u2 net6 A2 VDD VDD p w=0.685u l=0.18u
MU30-M_u1 net6 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt AN4D2BWP7T A1 A2 A3 A4 Z VDD VSS 
MU18_0-M_u2 Z net19 VSS VSS n w=1u l=0.18u
MU18_1-M_u2 Z net19 VSS VSS n w=1u l=0.18u
MU20-M_u5 net19 A1 XU20-net23 VSS n w=1u l=0.18u
MU20-M_u6 XU20-net23 A2 XU20-net26 VSS n w=1u l=0.18u
MU20-M_u7 XU20-net26 A3 XU20-net29 VSS n w=1u l=0.18u
MU20-M_u8 XU20-net29 A4 VSS VSS n w=1u l=0.18u
MU18_0-M_u3 Z net19 VDD VDD p w=1.37u l=0.18u
MU18_1-M_u3 Z net19 VDD VDD p w=1.37u l=0.18u
MU20-M_u4 net19 A4 VDD VDD p w=1.37u l=0.18u
MU20-M_u3 net19 A3 VDD VDD p w=1.37u l=0.18u
MU20-M_u2 net19 A2 VDD VDD p w=1.37u l=0.18u
MU20-M_u1 net19 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AN4D4BWP7T A1 A2 A3 A4 Z VDD VSS 
MU18_0-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU18_1-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU18_2-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU18_3-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MI4-M_u5 n0 A1 XI4-net23 VSS n w=1u l=0.18u
MI4-M_u6 XI4-net23 A2 XI4-net26 VSS n w=1u l=0.18u
MI4-M_u7 XI4-net26 A3 XI4-net29 VSS n w=1u l=0.18u
MI4-M_u8 XI4-net29 A4 VSS VSS n w=1u l=0.18u
MU30-M_u5 n0 A1 XU30-net23 VSS n w=1u l=0.18u
MU30-M_u6 XU30-net23 A2 XU30-net26 VSS n w=1u l=0.18u
MU30-M_u7 XU30-net26 A3 XU30-net29 VSS n w=1u l=0.18u
MU30-M_u8 XU30-net29 A4 VSS VSS n w=1u l=0.18u
MU18_0-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU18_1-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU18_2-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU18_3-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MI4-M_u4 n0 A4 VDD VDD p w=1.37u l=0.18u
MI4-M_u3 n0 A3 VDD VDD p w=1.37u l=0.18u
MI4-M_u2 n0 A2 VDD VDD p w=1.305u l=0.18u
MI4-M_u1 n0 A1 VDD VDD p w=1.305u l=0.18u
MU30-M_u4 n0 A4 VDD VDD p w=1.37u l=0.18u
MU30-M_u3 n0 A3 VDD VDD p w=1.37u l=0.18u
MU30-M_u2 n0 A2 VDD VDD p w=1.305u l=0.18u
MU30-M_u1 n0 A1 VDD VDD p w=1.305u l=0.18u
.ends
.subckt AN4XD1BWP7T A1 A2 A3 A4 Z VDD VSS 
M_u3-M_u2 Z net6 VSS VSS n w=1u l=0.18u
MU30-M_u5 net6 A1 XU30-net23 VSS n w=1u l=0.18u
MU30-M_u6 XU30-net23 A2 XU30-net26 VSS n w=1u l=0.18u
MU30-M_u7 XU30-net26 A3 XU30-net29 VSS n w=1u l=0.18u
MU30-M_u8 XU30-net29 A4 VSS VSS n w=1u l=0.18u
M_u3-M_u3 Z net6 VDD VDD p w=1.37u l=0.18u
MU30-M_u4 net6 A4 VDD VDD p w=1.37u l=0.18u
MU30-M_u3 net6 A3 VDD VDD p w=1.37u l=0.18u
MU30-M_u2 net6 A2 VDD VDD p w=1.37u l=0.18u
MU30-M_u1 net6 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ANTENNABWP7T I VDD VSS 
DI3 VSS I dn 0.2037p
.ends
.subckt AO211D0BWP7T A1 A2 B C Z VDD VSS 
M_u12 net27 C VSS VSS n w=0.5u l=0.18u
M_u13 net27 B VSS VSS n w=0.5u l=0.18u
MI12-M_u10 net27 A1 XI12-net17 VSS n w=0.5u l=0.18u
MI12-M_u11 XI12-net17 A2 VSS VSS n w=0.5u l=0.18u
MI8-M_u2 Z net27 VSS VSS n w=0.5u l=0.18u
MI8-M_u3 Z net27 VDD VDD p w=0.685u l=0.18u
M_u3 net11 A1 net27 VDD p w=0.685u l=0.18u
MI0 net11 A2 net27 VDD p w=0.685u l=0.18u
MI16-MI12 net11 B XI16-net11 VDD p w=0.685u l=0.18u
MI16-MI13 XI16-net11 C VDD VDD p w=0.685u l=0.18u
.ends
.subckt AO211D1BWP7T A1 A2 B C Z VDD VSS 
M_u12 net27 C VSS VSS n w=1u l=0.18u
M_u13 net27 B VSS VSS n w=1u l=0.18u
MI12-M_u10 net27 A1 XI12-net17 VSS n w=1u l=0.18u
MI12-M_u11 XI12-net17 A2 VSS VSS n w=1u l=0.18u
MI8-M_u2 Z net27 VSS VSS n w=1u l=0.18u
MI8-M_u3 Z net27 VDD VDD p w=1.37u l=0.18u
M_u3 net11 A1 net27 VDD p w=1.37u l=0.18u
MI0 net11 A2 net27 VDD p w=1.37u l=0.18u
MI16-MI12 net11 B XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 C VDD VDD p w=1.37u l=0.18u
.ends
.subckt AO211D2BWP7T A1 A2 B C Z VDD VSS 
M_u12 net27 C VSS VSS n w=1u l=0.18u
M_u13 net27 B VSS VSS n w=1u l=0.18u
MI12-M_u10 net27 A1 XI12-net17 VSS n w=1u l=0.18u
MI12-M_u11 XI12-net17 A2 VSS VSS n w=1u l=0.18u
MI8_0-M_u2 Z net27 VSS VSS n w=1u l=0.18u
MI8_1-M_u2 Z net27 VSS VSS n w=1u l=0.18u
MI8_0-M_u3 Z net27 VDD VDD p w=1.37u l=0.18u
MI8_1-M_u3 Z net27 VDD VDD p w=1.37u l=0.18u
M_u3 net11 A1 net27 VDD p w=1.37u l=0.18u
MI0 net11 A2 net27 VDD p w=1.37u l=0.18u
MI16-MI12 net11 B XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 C VDD VDD p w=1.37u l=0.18u
.ends
.subckt AO21D0BWP7T A1 A2 B Z VDD VSS 
MI7 net32 A2 VSS VSS n w=0.5u l=0.18u
M_u7 net59 A1 net32 VSS n w=0.5u l=0.18u
MI6 net59 B VSS VSS n w=0.5u l=0.18u
MI8-M_u2 Z net59 VSS VSS n w=0.5u l=0.18u
MI8-M_u3 Z net59 VDD VDD p w=0.685u l=0.18u
M_u3 net22 A1 net59 VDD p w=0.685u l=0.18u
M_u4 net22 A2 net59 VDD p w=0.685u l=0.18u
M_u2 net22 B VDD VDD p w=0.685u l=0.18u
.ends
.subckt AO21D1BWP7T A1 A2 B Z VDD VSS 
MI7 net32 A2 VSS VSS n w=1u l=0.18u
M_u7 net59 A1 net32 VSS n w=1u l=0.18u
MI6 net59 B VSS VSS n w=1u l=0.18u
MI8-M_u2 Z net59 VSS VSS n w=1u l=0.18u
MI8-M_u3 Z net59 VDD VDD p w=1.37u l=0.18u
M_u3 net22 A1 net59 VDD p w=1.37u l=0.18u
M_u4 net22 A2 net59 VDD p w=1.37u l=0.18u
M_u2 net22 B VDD VDD p w=1.37u l=0.18u
.ends
.subckt AO21D2BWP7T A1 A2 B Z VDD VSS 
MI7 net32 A2 VSS VSS n w=1u l=0.18u
M_u7 net59 A1 net32 VSS n w=1u l=0.18u
MI6 net59 B VSS VSS n w=1u l=0.18u
MI8_0-M_u2 Z net59 VSS VSS n w=1u l=0.18u
MI8_1-M_u2 Z net59 VSS VSS n w=1u l=0.18u
MI8_0-M_u3 Z net59 VDD VDD p w=1.37u l=0.18u
MI8_1-M_u3 Z net59 VDD VDD p w=1.37u l=0.18u
M_u3 net22 A1 net59 VDD p w=1.37u l=0.18u
M_u4 net22 A2 net59 VDD p w=1.37u l=0.18u
M_u2 net22 B VDD VDD p w=1.37u l=0.18u
.ends
.subckt AO221D0BWP7T A1 A2 B1 B2 C Z VDD VSS 
MU20 net31 C VSS VSS n w=0.5u l=0.18u
MI17-M_u10 net31 B1 XI17-net17 VSS n w=0.5u l=0.18u
MI17-M_u11 XI17-net17 B2 VSS VSS n w=0.5u l=0.18u
MI1-M_u10 net31 A1 XI1-net17 VSS n w=0.5u l=0.18u
MI1-M_u11 XI1-net17 A2 VSS VSS n w=0.5u l=0.18u
MI8-M_u2 Z net31 VSS VSS n w=0.5u l=0.18u
MI8-M_u3 Z net31 VDD VDD p w=0.685u l=0.18u
MI5 net30 A1 net31 VDD p w=0.685u l=0.18u
MI4 net30 A2 net31 VDD p w=0.685u l=0.18u
MU22 VDD C net36 VDD p w=0.685u l=0.18u
MI2 net36 B2 net30 VDD p w=0.685u l=0.18u
MI3 net36 B1 net30 VDD p w=0.685u l=0.18u
.ends
.subckt AO221D1BWP7T A1 A2 B1 B2 C Z VDD VSS 
MU20 net31 C VSS VSS n w=1u l=0.18u
MI17-M_u10 net31 B1 XI17-net17 VSS n w=1u l=0.18u
MI17-M_u11 XI17-net17 B2 VSS VSS n w=1u l=0.18u
MI1-M_u10 net31 A1 XI1-net17 VSS n w=1u l=0.18u
MI1-M_u11 XI1-net17 A2 VSS VSS n w=1u l=0.18u
MI8-M_u2 Z net31 VSS VSS n w=1u l=0.18u
MI8-M_u3 Z net31 VDD VDD p w=1.37u l=0.18u
MI5 net30 A1 net31 VDD p w=1.37u l=0.18u
MI4 net30 A2 net31 VDD p w=1.37u l=0.18u
MU22 VDD C net36 VDD p w=1.37u l=0.18u
MI2 net36 B2 net30 VDD p w=1.37u l=0.18u
MI3 net36 B1 net30 VDD p w=1.37u l=0.18u
.ends
.subckt AO221D2BWP7T A1 A2 B1 B2 C Z VDD VSS 
MU20 net31 C VSS VSS n w=1u l=0.18u
MI17-M_u10 net31 B1 XI17-net17 VSS n w=1u l=0.18u
MI17-M_u11 XI17-net17 B2 VSS VSS n w=1u l=0.18u
MI1-M_u10 net31 A1 XI1-net17 VSS n w=1u l=0.18u
MI1-M_u11 XI1-net17 A2 VSS VSS n w=1u l=0.18u
MI8_0-M_u2 Z net31 VSS VSS n w=1u l=0.18u
MI8_1-M_u2 Z net31 VSS VSS n w=1u l=0.18u
MI8_0-M_u3 Z net31 VDD VDD p w=1.37u l=0.18u
MI8_1-M_u3 Z net31 VDD VDD p w=1.37u l=0.18u
MI5 net30 A1 net31 VDD p w=1.37u l=0.18u
MI4 net30 A2 net31 VDD p w=1.37u l=0.18u
MU22 VDD C net36 VDD p w=1.37u l=0.18u
MI2 net36 B2 net30 VDD p w=1.37u l=0.18u
MI3 net36 B1 net30 VDD p w=1.37u l=0.18u
.ends
.subckt AO222D0BWP7T A1 A2 B1 B2 C1 C2 Z VDD VSS 
MI14-M_u10 net39 C1 XI14-net17 VSS n w=0.5u l=0.18u
MI14-M_u11 XI14-net17 C2 VSS VSS n w=0.5u l=0.18u
MI6-M_u10 net39 A1 XI6-net17 VSS n w=0.5u l=0.18u
MI6-M_u11 XI6-net17 A2 VSS VSS n w=0.5u l=0.18u
MI13-M_u10 net39 B1 XI13-net17 VSS n w=0.5u l=0.18u
MI13-M_u11 XI13-net17 B2 VSS VSS n w=0.5u l=0.18u
MI15-M_u2 Z net39 VSS VSS n w=0.5u l=0.18u
MI15-M_u3 Z net39 VDD VDD p w=0.685u l=0.18u
MI8 VDD C1 net22 VDD p w=0.685u l=0.18u
MU27 VDD C2 net22 VDD p w=0.685u l=0.18u
MI12 net16 A1 net39 VDD p w=0.685u l=0.18u
MI11 net16 A2 net39 VDD p w=0.685u l=0.18u
MI10 net22 B1 net16 VDD p w=0.685u l=0.18u
MI9 net22 B2 net16 VDD p w=0.685u l=0.18u
.ends
.subckt AO222D1BWP7T A1 A2 B1 B2 C1 C2 Z VDD VSS 
MI14-M_u10 net39 C1 XI14-net17 VSS n w=1u l=0.18u
MI14-M_u11 XI14-net17 C2 VSS VSS n w=1u l=0.18u
MI6-M_u10 net39 A1 XI6-net17 VSS n w=1u l=0.18u
MI6-M_u11 XI6-net17 A2 VSS VSS n w=1u l=0.18u
MI13-M_u10 net39 B1 XI13-net17 VSS n w=1u l=0.18u
MI13-M_u11 XI13-net17 B2 VSS VSS n w=1u l=0.18u
MI15-M_u2 Z net39 VSS VSS n w=1u l=0.18u
MI15-M_u3 Z net39 VDD VDD p w=1.37u l=0.18u
MI8 VDD C1 net22 VDD p w=1.37u l=0.18u
MU27 VDD C2 net22 VDD p w=1.37u l=0.18u
MI12 net16 A1 net39 VDD p w=1.37u l=0.18u
MI11 net16 A2 net39 VDD p w=1.37u l=0.18u
MI10 net22 B1 net16 VDD p w=1.37u l=0.18u
MI9 net22 B2 net16 VDD p w=1.37u l=0.18u
.ends
.subckt AO222D2BWP7T A1 A2 B1 B2 C1 C2 Z VDD VSS 
MI14-M_u10 net39 C1 XI14-net17 VSS n w=1u l=0.18u
MI14-M_u11 XI14-net17 C2 VSS VSS n w=1u l=0.18u
MI6-M_u10 net39 A1 XI6-net17 VSS n w=1u l=0.18u
MI6-M_u11 XI6-net17 A2 VSS VSS n w=1u l=0.18u
MI13-M_u10 net39 B1 XI13-net17 VSS n w=1u l=0.18u
MI13-M_u11 XI13-net17 B2 VSS VSS n w=1u l=0.18u
MI15_0-M_u2 Z net39 VSS VSS n w=1u l=0.18u
MI15_1-M_u2 Z net39 VSS VSS n w=1u l=0.18u
MI15_0-M_u3 Z net39 VDD VDD p w=1.37u l=0.18u
MI15_1-M_u3 Z net39 VDD VDD p w=1.37u l=0.18u
MI8 VDD C1 net22 VDD p w=1.37u l=0.18u
MU27 VDD C2 net22 VDD p w=1.37u l=0.18u
MI12 net16 A1 net39 VDD p w=1.37u l=0.18u
MI11 net16 A2 net39 VDD p w=1.37u l=0.18u
MI10 net22 B1 net16 VDD p w=1.37u l=0.18u
MI9 net22 B2 net16 VDD p w=1.37u l=0.18u
.ends
.subckt AO22D0BWP7T A1 A2 B1 B2 Z VDD VSS 
MI18 net29 A2 VSS VSS n w=0.5u l=0.18u
MI16 net26 B1 net20 VSS n w=0.5u l=0.18u
M_u7 net26 A1 net29 VSS n w=0.5u l=0.18u
MI17 net20 B2 VSS VSS n w=0.5u l=0.18u
MI8-M_u2 Z net26 VSS VSS n w=0.5u l=0.18u
MI8-M_u3 Z net26 VDD VDD p w=0.685u l=0.18u
MI14 net26 A1 net40 VDD p w=0.685u l=0.18u
MI15 net26 A2 net40 VDD p w=0.685u l=0.18u
M_u2 net40 B2 VDD VDD p w=0.685u l=0.18u
MI13 net40 B1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt AO22D1BWP7T A1 A2 B1 B2 Z VDD VSS 
MI28 net52 A1 net37 VSS n w=1u l=0.18u
MI21 net52 B1 net31 VSS n w=1u l=0.18u
MI22 net31 B2 VSS VSS n w=1u l=0.18u
MI29 net37 A2 VSS VSS n w=1u l=0.18u
MI20-M_u2 Z net52 VSS VSS n w=1u l=0.18u
MI20-M_u3 Z net52 VDD VDD p w=1.37u l=0.18u
MI15 net54 B2 VDD VDD p w=1.37u l=0.18u
MI18 net52 A2 net54 VDD p w=1.37u l=0.18u
MI17 net54 B1 VDD VDD p w=1.37u l=0.18u
MI19 net52 A1 net54 VDD p w=1.37u l=0.18u
.ends
.subckt AO22D2BWP7T A1 A2 B1 B2 Z VDD VSS 
MI28 net52 A1 net37 VSS n w=1u l=0.18u
MI21 net52 B1 net31 VSS n w=1u l=0.18u
MI22 net31 B2 VSS VSS n w=1u l=0.18u
MI29 net37 A2 VSS VSS n w=1u l=0.18u
MI20_0-M_u2 Z net52 VSS VSS n w=1u l=0.18u
MI20_1-M_u2 Z net52 VSS VSS n w=1u l=0.18u
MI20_0-M_u3 Z net52 VDD VDD p w=1.37u l=0.18u
MI20_1-M_u3 Z net52 VDD VDD p w=1.37u l=0.18u
MI15 net54 B2 VDD VDD p w=1.37u l=0.18u
MI18 net52 A2 net54 VDD p w=1.37u l=0.18u
MI17 net54 B1 VDD VDD p w=1.37u l=0.18u
MI19 net52 A1 net54 VDD p w=1.37u l=0.18u
.ends
.subckt AO31D0BWP7T A1 A2 A3 B Z VDD VSS 
MU14 net26 B VSS VSS n w=0.5u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=0.5u l=0.18u
MI20-M_u10 net26 A1 XI20-net17 VSS n w=0.5u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=0.5u l=0.18u
MI8-M_u2 Z net26 VSS VSS n w=0.5u l=0.18u
MI8-M_u3 Z net26 VDD VDD p w=0.685u l=0.18u
MU17 net26 A1 net19 VDD p w=0.685u l=0.18u
MU18 net26 A3 net19 VDD p w=0.685u l=0.18u
MU16 net26 A2 net19 VDD p w=0.685u l=0.18u
MU20 net19 B VDD VDD p w=0.685u l=0.18u
.ends
.subckt AO31D1BWP7T A1 A2 A3 B Z VDD VSS 
MU14 net26 B VSS VSS n w=1u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=1u l=0.18u
MI20-M_u10 net26 A1 XI20-net17 VSS n w=1u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=1u l=0.18u
MI8-M_u2 Z net26 VSS VSS n w=1u l=0.18u
MI8-M_u3 Z net26 VDD VDD p w=1.37u l=0.18u
MU17 net26 A1 net19 VDD p w=1.37u l=0.18u
MU18 net26 A3 net19 VDD p w=1.37u l=0.18u
MU16 net26 A2 net19 VDD p w=1.37u l=0.18u
MU20 net19 B VDD VDD p w=1.37u l=0.18u
.ends
.subckt AO31D2BWP7T A1 A2 A3 B Z VDD VSS 
MU14 net26 B VSS VSS n w=1u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=1u l=0.18u
MI20-M_u10 net26 A1 XI20-net17 VSS n w=1u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=1u l=0.18u
MI8_0-M_u2 Z net26 VSS VSS n w=1u l=0.18u
MI8_1-M_u2 Z net26 VSS VSS n w=1u l=0.18u
MI8_0-M_u3 Z net26 VDD VDD p w=1.37u l=0.18u
MI8_1-M_u3 Z net26 VDD VDD p w=1.37u l=0.18u
MU17 net26 A1 net19 VDD p w=1.37u l=0.18u
MU18 net26 A3 net19 VDD p w=1.37u l=0.18u
MU16 net26 A2 net19 VDD p w=1.37u l=0.18u
MU20 net19 B VDD VDD p w=1.37u l=0.18u
.ends
.subckt AO32D0BWP7T A1 A2 A3 B1 B2 Z VDD VSS 
MI17-M_u10 net27 B1 XI17-net17 VSS n w=0.5u l=0.18u
MI17-M_u11 XI17-net17 B2 VSS VSS n w=0.5u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=0.5u l=0.18u
MI20-M_u10 net27 A1 XI20-net17 VSS n w=0.5u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=0.5u l=0.18u
MI8-M_u2 Z net27 VSS VSS n w=0.5u l=0.18u
MI8-M_u3 Z net27 VDD VDD p w=0.685u l=0.18u
MU17 net27 A1 net23 VDD p w=0.685u l=0.18u
MU18 net27 A3 net23 VDD p w=0.685u l=0.18u
MU16 net27 A2 net23 VDD p w=0.685u l=0.18u
MU20 net23 B1 VDD VDD p w=0.685u l=0.18u
MU19 net23 B2 VDD VDD p w=0.685u l=0.18u
.ends
.subckt AO32D1BWP7T A1 A2 A3 B1 B2 Z VDD VSS 
MI17-M_u10 net27 B1 XI17-net17 VSS n w=1u l=0.18u
MI17-M_u11 XI17-net17 B2 VSS VSS n w=1u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=1u l=0.18u
MI20-M_u10 net27 A1 XI20-net17 VSS n w=1u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=1u l=0.18u
MI8-M_u2 Z net27 VSS VSS n w=1u l=0.18u
MI8-M_u3 Z net27 VDD VDD p w=1.37u l=0.18u
MU17 net27 A1 net23 VDD p w=1.37u l=0.18u
MU18 net27 A3 net23 VDD p w=1.37u l=0.18u
MU16 net27 A2 net23 VDD p w=1.37u l=0.18u
MU20 net23 B1 VDD VDD p w=1.37u l=0.18u
MU19 net23 B2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AO32D2BWP7T A1 A2 A3 B1 B2 Z VDD VSS 
MI17-M_u10 net27 B1 XI17-net17 VSS n w=1u l=0.18u
MI17-M_u11 XI17-net17 B2 VSS VSS n w=1u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=1u l=0.18u
MI20-M_u10 net27 A1 XI20-net17 VSS n w=1u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=1u l=0.18u
MI8_0-M_u2 Z net27 VSS VSS n w=1u l=0.18u
MI8_1-M_u2 Z net27 VSS VSS n w=1u l=0.18u
MI8_0-M_u3 Z net27 VDD VDD p w=1.37u l=0.18u
MI8_1-M_u3 Z net27 VDD VDD p w=1.37u l=0.18u
MU17 net27 A1 net23 VDD p w=1.37u l=0.18u
MU18 net27 A3 net23 VDD p w=1.37u l=0.18u
MU16 net27 A2 net23 VDD p w=1.37u l=0.18u
MU20 net23 B1 VDD VDD p w=1.37u l=0.18u
MU19 net23 B2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AO33D0BWP7T A1 A2 A3 B1 B2 B3 Z VDD VSS 
MI14-MI12 XI14-net13 A3 VSS VSS n w=0.5u l=0.18u
MI14-M_u10 net30 A1 XI14-net17 VSS n w=0.5u l=0.18u
MI14-M_u11 XI14-net17 A2 XI14-net13 VSS n w=0.5u l=0.18u
MI7-MI12 XI7-net13 B3 VSS VSS n w=0.5u l=0.18u
MI7-M_u10 net30 B1 XI7-net17 VSS n w=0.5u l=0.18u
MI7-M_u11 XI7-net17 B2 XI7-net13 VSS n w=0.5u l=0.18u
MI8-M_u2 Z net30 VSS VSS n w=0.5u l=0.18u
MI8-M_u3 Z net30 VDD VDD p w=0.685u l=0.18u
MI6 net40 A1 net30 VDD p w=0.685u l=0.18u
M_u16 VDD B3 net40 VDD p w=0.685u l=0.18u
MI3 VDD B1 net40 VDD p w=0.685u l=0.18u
MI4 net40 A3 net30 VDD p w=0.685u l=0.18u
MI5 net40 A2 net30 VDD p w=0.685u l=0.18u
MI2 VDD B2 net40 VDD p w=0.685u l=0.18u
.ends
.subckt AO33D1BWP7T A1 A2 A3 B1 B2 B3 Z VDD VSS 
MI14-MI12 XI14-net13 A3 VSS VSS n w=1u l=0.18u
MI14-M_u10 net30 A1 XI14-net17 VSS n w=1u l=0.18u
MI14-M_u11 XI14-net17 A2 XI14-net13 VSS n w=1u l=0.18u
MI15-MI12 XI15-net13 B3 VSS VSS n w=1u l=0.18u
MI15-M_u10 net30 B1 XI15-net17 VSS n w=1u l=0.18u
MI15-M_u11 XI15-net17 B2 XI15-net13 VSS n w=1u l=0.18u
MI8-M_u2 Z net30 VSS VSS n w=1u l=0.18u
MI8-M_u3 Z net30 VDD VDD p w=1.37u l=0.18u
MI6 net40 A1 net30 VDD p w=1.37u l=0.18u
MI13 VDD B3 net40 VDD p w=1.37u l=0.18u
MI11 VDD B1 net40 VDD p w=1.37u l=0.18u
MI10 net40 A3 net30 VDD p w=1.37u l=0.18u
MI9 net40 A2 net30 VDD p w=1.37u l=0.18u
MI12 VDD B2 net40 VDD p w=1.37u l=0.18u
.ends
.subckt AO33D2BWP7T A1 A2 A3 B1 B2 B3 Z VDD VSS 
MI14-MI12 XI14-net13 A3 VSS VSS n w=1u l=0.18u
MI14-M_u10 net30 A1 XI14-net17 VSS n w=1u l=0.18u
MI14-M_u11 XI14-net17 A2 XI14-net13 VSS n w=1u l=0.18u
MI15-MI12 XI15-net13 B3 VSS VSS n w=1u l=0.18u
MI15-M_u10 net30 B1 XI15-net17 VSS n w=1u l=0.18u
MI15-M_u11 XI15-net17 B2 XI15-net13 VSS n w=1u l=0.18u
MI8_0-M_u2 Z net30 VSS VSS n w=1u l=0.18u
MI8_1-M_u2 Z net30 VSS VSS n w=1u l=0.18u
MI8_0-M_u3 Z net30 VDD VDD p w=1.37u l=0.18u
MI8_1-M_u3 Z net30 VDD VDD p w=1.37u l=0.18u
MI6 net40 A1 net30 VDD p w=1.37u l=0.18u
MI13 VDD B3 net40 VDD p w=1.37u l=0.18u
MI11 VDD B1 net40 VDD p w=1.37u l=0.18u
MI10 net40 A3 net30 VDD p w=1.37u l=0.18u
MI9 net40 A2 net30 VDD p w=1.37u l=0.18u
MI12 VDD B2 net40 VDD p w=1.37u l=0.18u
.ends
.subckt AOI211D0BWP7T A1 A2 B C ZN VDD VSS 
M_u12 ZN C VSS VSS n w=0.5u l=0.18u
M_u13 ZN B VSS VSS n w=0.5u l=0.18u
MI12-M_u10 ZN A1 XI12-net17 VSS n w=0.5u l=0.18u
MI12-M_u11 XI12-net17 A2 VSS VSS n w=0.5u l=0.18u
M_u3 net11 A1 ZN VDD p w=0.685u l=0.18u
MI0 net11 A2 ZN VDD p w=0.685u l=0.18u
MI16-MI12 net11 B XI16-net11 VDD p w=0.685u l=0.18u
MI16-MI13 XI16-net11 C VDD VDD p w=0.685u l=0.18u
.ends
.subckt AOI211D1BWP7T A1 A2 B C ZN VDD VSS 
M_u12 ZN C VSS VSS n w=1u l=0.18u
M_u13 ZN B VSS VSS n w=1u l=0.18u
MI17-M_u10 ZN A1 XI17-net17 VSS n w=1u l=0.18u
MI17-M_u11 XI17-net17 A2 VSS VSS n w=1u l=0.18u
M_u3 net71 A1 ZN VDD p w=1.37u l=0.18u
M_u2 net71 A2 ZN VDD p w=1.37u l=0.18u
MI19-MI12 net71 B XI19-net11 VDD p w=1.37u l=0.18u
MI19-MI13 XI19-net11 C VDD VDD p w=1.37u l=0.18u
.ends
.subckt AOI211D2BWP7T A1 A2 B C ZN VDD VSS 
M_u12_0 ZN C VSS VSS n w=1u l=0.18u
M_u12_1 ZN C VSS VSS n w=1u l=0.18u
M_u13_0 ZN B VSS VSS n w=1u l=0.18u
M_u13_1 ZN B VSS VSS n w=1u l=0.18u
MI17_0-M_u10 ZN A1 XI17_0-net17 VSS n w=1u l=0.18u
MI17_0-M_u11 XI17_0-net17 A2 VSS VSS n w=1u l=0.18u
MI17_1-M_u10 ZN A1 XI17_1-net17 VSS n w=1u l=0.18u
MI17_1-M_u11 XI17_1-net17 A2 VSS VSS n w=1u l=0.18u
M_u3_0 net34 A1 ZN VDD p w=1.37u l=0.18u
M_u3_1 net34 A1 ZN VDD p w=1.37u l=0.18u
M_u2_0 net34 A2 ZN VDD p w=1.37u l=0.18u
M_u2_1 net34 A2 ZN VDD p w=1.37u l=0.18u
MI19-MI12 net34 B XI19-net11 VDD p w=1.37u l=0.18u
MI19-MI13 XI19-net11 C VDD VDD p w=1.37u l=0.18u
MI2-MI12 net34 B XI2-net11 VDD p w=1.37u l=0.18u
MI2-MI13 XI2-net11 C VDD VDD p w=1.37u l=0.18u
.ends
.subckt AOI211XD0BWP7T A1 A2 B C ZN VDD VSS 
M_u12 ZN C VSS VSS n w=0.5u l=0.18u
M_u13 ZN B VSS VSS n w=0.5u l=0.18u
MI12-M_u10 ZN A1 XI12-net17 VSS n w=0.5u l=0.18u
MI12-M_u11 XI12-net17 A2 VSS VSS n w=0.5u l=0.18u
M_u3 net11 A1 ZN VDD p w=1.37u l=0.18u
MI0 net11 A2 ZN VDD p w=1.37u l=0.18u
MI16-MI12 net11 B XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 C VDD VDD p w=1.37u l=0.18u
.ends
.subckt AOI211XD1BWP7T A1 A2 B C ZN VDD VSS 
M_u12 ZN C VSS VSS n w=1u l=0.18u
M_u13 ZN B VSS VSS n w=1u l=0.18u
MI17-M_u10 ZN A1 XI17-net17 VSS n w=1u l=0.18u
MI17-M_u11 XI17-net17 A2 VSS VSS n w=1u l=0.18u
MI1 net034 B net030 VDD p w=1.37u l=0.18u
MI0 VDD C net034 VDD p w=1.37u l=0.18u
MI2 net034 B net030 VDD p w=1.37u l=0.18u
MI3 VDD C net034 VDD p w=1.37u l=0.18u
M_u3 net030 A1 ZN VDD p w=2.74u l=0.18u
M_u2 net030 A2 ZN VDD p w=2.74u l=0.18u
.ends
.subckt AOI211XD2BWP7T A1 A2 B C ZN VDD VSS 
M_u12_0 ZN C VSS VSS n w=1u l=0.18u
M_u12_1 ZN C VSS VSS n w=1u l=0.18u
M_u13_0 ZN B VSS VSS n w=1u l=0.18u
M_u13_1 ZN B VSS VSS n w=1u l=0.18u
MI17-M_u10 ZN A1 XI17-net17 VSS n w=2u l=0.18u
MI17-M_u11 XI17-net17 A2 VSS VSS n w=2u l=0.18u
M_u3 net034 A1 ZN VDD p w=5.48u l=0.18u
M_u2 net034 A2 ZN VDD p w=5.48u l=0.18u
MI19-MI12 net034 B XI19-net11 VDD p w=5.48u l=0.18u
MI19-MI13 XI19-net11 C VDD VDD p w=5.48u l=0.18u
.ends
.subckt AOI21D0BWP7T A1 A2 B ZN VDD VSS 
MI2 ZN A1 net27 VSS n w=0.5u l=0.18u
MI7 net27 A2 VSS VSS n w=0.5u l=0.18u
MI6 ZN B VSS VSS n w=0.5u l=0.18u
MI5 ZN A2 net13 VDD p w=0.685u l=0.18u
M_u2 net13 B VDD VDD p w=0.685u l=0.18u
MI4 ZN A1 net13 VDD p w=0.685u l=0.18u
.ends
.subckt AOI21D1BWP7T A1 A2 B ZN VDD VSS 
MI2 ZN A1 net27 VSS n w=1u l=0.18u
MI3 net27 A2 VSS VSS n w=1u l=0.18u
M_u7 ZN B VSS VSS n w=1u l=0.18u
M_u4 net13 A2 ZN VDD p w=1.37u l=0.18u
M_u2 net13 B VDD VDD p w=1.37u l=0.18u
M_u3 net13 A1 ZN VDD p w=1.37u l=0.18u
.ends
.subckt AOI21D2BWP7T A1 A2 B ZN VDD VSS 
MI2 ZN A1 p0 VSS n w=1u l=0.18u
MI12 p0 A2 VSS VSS n w=1u l=0.18u
MI13 ZN A1 net23 VSS n w=1u l=0.18u
MI14 net23 A2 VSS VSS n w=1u l=0.18u
MI11_0 ZN B VSS VSS n w=1u l=0.18u
MI11_1 ZN B VSS VSS n w=1u l=0.18u
MI8 ZN A2 net74 VDD p w=2.74u l=0.18u
M_u2 net74 B VDD VDD p w=2.74u l=0.18u
MI9 ZN A1 net74 VDD p w=2.74u l=0.18u
.ends
.subckt AOI221D0BWP7T A1 A2 B1 B2 C ZN VDD VSS 
MU20 ZN C VSS VSS n w=0.5u l=0.18u
MI17-M_u10 ZN B1 XI17-net17 VSS n w=0.5u l=0.18u
MI17-M_u11 XI17-net17 B2 VSS VSS n w=0.5u l=0.18u
MI1-M_u10 ZN A1 XI1-net17 VSS n w=0.5u l=0.18u
MI1-M_u11 XI1-net17 A2 VSS VSS n w=0.5u l=0.18u
MI5 net30 A1 ZN VDD p w=0.685u l=0.18u
MI4 net30 A2 ZN VDD p w=0.685u l=0.18u
MU22 VDD C net36 VDD p w=0.685u l=0.18u
MI2 net36 B2 net30 VDD p w=0.685u l=0.18u
MI3 net36 B1 net30 VDD p w=0.685u l=0.18u
.ends
.subckt AOI221D1BWP7T A1 A2 B1 B2 C ZN VDD VSS 
MU20 ZN C VSS VSS n w=1u l=0.18u
MI17-M_u10 ZN B1 XI17-net17 VSS n w=1u l=0.18u
MI17-M_u11 XI17-net17 B2 VSS VSS n w=1u l=0.18u
MI1-M_u10 ZN A1 XI1-net17 VSS n w=1u l=0.18u
MI1-M_u11 XI1-net17 A2 VSS VSS n w=1u l=0.18u
M_u5 net36 B2 net30 VDD p w=1.37u l=0.18u
MU22 VDD C net36 VDD p w=1.37u l=0.18u
M_u2 net30 A1 ZN VDD p w=1.37u l=0.18u
M_u3 net30 A2 ZN VDD p w=1.37u l=0.18u
M_u4 net36 B1 net30 VDD p w=1.37u l=0.18u
.ends
.subckt AOI221D2BWP7T A1 A2 B1 B2 C ZN VDD VSS 
MU20 ZN C VSS VSS n w=2u l=0.18u
MI17_0-M_u10 ZN B1 XI17_0-net17 VSS n w=1u l=0.18u
MI17_0-M_u11 XI17_0-net17 B2 VSS VSS n w=1u l=0.18u
MI17_1-M_u10 ZN B1 XI17_1-net17 VSS n w=1u l=0.18u
MI17_1-M_u11 XI17_1-net17 B2 VSS VSS n w=1u l=0.18u
MI8_0-M_u10 ZN A1 XI8_0-net17 VSS n w=1u l=0.18u
MI8_0-M_u11 XI8_0-net17 A2 VSS VSS n w=1u l=0.18u
MI8_1-M_u10 ZN A1 XI8_1-net17 VSS n w=1u l=0.18u
MI8_1-M_u11 XI8_1-net17 A2 VSS VSS n w=1u l=0.18u
MI7 net27 A1 ZN VDD p w=2.74u l=0.18u
MI4 net33 B2 net27 VDD p w=2.74u l=0.18u
MU22 VDD C net33 VDD p w=2.74u l=0.18u
MI6 net27 A2 ZN VDD p w=2.74u l=0.18u
MI5 net33 B1 net27 VDD p w=2.74u l=0.18u
.ends
.subckt AOI222D0BWP7T A1 A2 B1 B2 C1 C2 ZN VDD VSS 
MI14-M_u10 ZN C1 XI14-net17 VSS n w=0.5u l=0.18u
MI14-M_u11 XI14-net17 C2 VSS VSS n w=0.5u l=0.18u
MI6-M_u10 ZN A1 XI6-net17 VSS n w=0.5u l=0.18u
MI6-M_u11 XI6-net17 A2 VSS VSS n w=0.5u l=0.18u
MI13-M_u10 ZN B1 XI13-net17 VSS n w=0.5u l=0.18u
MI13-M_u11 XI13-net17 B2 VSS VSS n w=0.5u l=0.18u
MI8 VDD C1 net22 VDD p w=0.685u l=0.18u
MU27 VDD C2 net22 VDD p w=0.685u l=0.18u
MI12 net16 A1 ZN VDD p w=0.685u l=0.18u
MI11 net16 A2 ZN VDD p w=0.685u l=0.18u
MI10 net22 B1 net16 VDD p w=0.685u l=0.18u
MI9 net22 B2 net16 VDD p w=0.685u l=0.18u
.ends
.subckt AOI222D1BWP7T A1 A2 B1 B2 C1 C2 ZN VDD VSS 
MI17-M_u10 ZN C1 XI17-net17 VSS n w=1u l=0.18u
MI17-M_u11 XI17-net17 C2 VSS VSS n w=1u l=0.18u
MI6-M_u10 ZN A1 XI6-net17 VSS n w=1u l=0.18u
MI6-M_u11 XI6-net17 A2 VSS VSS n w=1u l=0.18u
MI7-M_u10 ZN B1 XI7-net17 VSS n w=1u l=0.18u
MI7-M_u11 XI7-net17 B2 VSS VSS n w=1u l=0.18u
MU22 VDD C1 net22 VDD p w=1.37u l=0.18u
MU27 VDD C2 net22 VDD p w=1.37u l=0.18u
M_u2 net16 A1 ZN VDD p w=1.37u l=0.18u
M_u3 net16 A2 ZN VDD p w=1.37u l=0.18u
M_u4 net22 B1 net16 VDD p w=1.37u l=0.18u
M_u5 net22 B2 net16 VDD p w=1.37u l=0.18u
.ends
.subckt AOI222D2BWP7T A1 A2 B1 B2 C1 C2 ZN VDD VSS 
MI21_0-M_u10 ZN C1 XI21_0-net17 VSS n w=1u l=0.18u
MI21_0-M_u11 XI21_0-net17 C2 VSS VSS n w=1u l=0.18u
MI21_1-M_u10 ZN C1 XI21_1-net17 VSS n w=1u l=0.18u
MI21_1-M_u11 XI21_1-net17 C2 VSS VSS n w=1u l=0.18u
MI6_0-M_u10 ZN A1 XI6_0-net17 VSS n w=1u l=0.18u
MI6_0-M_u11 XI6_0-net17 A2 VSS VSS n w=1u l=0.18u
MI6_1-M_u10 ZN A1 XI6_1-net17 VSS n w=1u l=0.18u
MI6_1-M_u11 XI6_1-net17 A2 VSS VSS n w=1u l=0.18u
MI20_0-M_u10 ZN B1 XI20_0-net17 VSS n w=1u l=0.18u
MI20_0-M_u11 XI20_0-net17 B2 VSS VSS n w=1u l=0.18u
MI20_1-M_u10 ZN B1 XI20_1-net17 VSS n w=1u l=0.18u
MI20_1-M_u11 XI20_1-net17 B2 VSS VSS n w=1u l=0.18u
MI15 VDD C1 net35 VDD p w=2.74u l=0.18u
MU27 VDD C2 net35 VDD p w=2.74u l=0.18u
MI25 net29 A1 ZN VDD p w=2.74u l=0.18u
MI24 net29 A2 ZN VDD p w=2.74u l=0.18u
MI23 net35 B1 net29 VDD p w=2.74u l=0.18u
MI22 net35 B2 net29 VDD p w=2.74u l=0.18u
.ends
.subckt AOI22D0BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI16 ZN B1 net29 VSS n w=0.5u l=0.18u
MI15 net29 B2 VSS VSS n w=0.5u l=0.18u
MI9 ZN A1 net23 VSS n w=0.5u l=0.18u
MI14 net23 A2 VSS VSS n w=0.5u l=0.18u
MI13 net20 A1 ZN VDD p w=0.685u l=0.18u
MI12 net20 A2 ZN VDD p w=0.685u l=0.18u
MI11 VDD B1 net20 VDD p w=0.685u l=0.18u
M_u5 VDD B2 net20 VDD p w=0.685u l=0.18u
.ends
.subckt AOI22D1BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI3 ZN B1 net29 VSS n w=1u l=0.18u
MI8 net29 B2 VSS VSS n w=1u l=0.18u
MI9 ZN A1 net23 VSS n w=1u l=0.18u
MI10 net23 A2 VSS VSS n w=1u l=0.18u
M_u2 net20 A1 ZN VDD p w=1.37u l=0.18u
M_u4 VDD B1 net20 VDD p w=1.37u l=0.18u
M_u3 net20 A2 ZN VDD p w=1.37u l=0.18u
M_u5 VDD B2 net20 VDD p w=1.37u l=0.18u
.ends
.subckt AOI22D2BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI16 ZN B1 net29 VSS n w=1u l=0.18u
MI15 net29 B2 VSS VSS n w=1u l=0.18u
MI17 ZN B1 net39 VSS n w=1u l=0.18u
MI18 net39 B2 VSS VSS n w=1u l=0.18u
MI20 net23 A2 VSS VSS n w=1u l=0.18u
MI22 net27 A2 VSS VSS n w=1u l=0.18u
MI21 ZN A1 net27 VSS n w=1u l=0.18u
MI19 ZN A1 net23 VSS n w=1u l=0.18u
MI13 net20 A1 ZN VDD p w=2.74u l=0.18u
M_u4 VDD B1 net20 VDD p w=2.74u l=0.18u
MI12 net20 A2 ZN VDD p w=2.74u l=0.18u
MI11 VDD B2 net20 VDD p w=2.74u l=0.18u
.ends
.subckt AOI31D0BWP7T A1 A2 A3 B ZN VDD VSS 
MU14 ZN B VSS VSS n w=0.5u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=0.5u l=0.18u
MI20-M_u10 ZN A1 XI20-net17 VSS n w=0.5u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=0.5u l=0.18u
MI3 ZN A1 net19 VDD p w=0.685u l=0.18u
MI1 ZN A3 net19 VDD p w=0.685u l=0.18u
MI2 ZN A2 net19 VDD p w=0.685u l=0.18u
MU20 net19 B VDD VDD p w=0.685u l=0.18u
.ends
.subckt AOI31D1BWP7T A1 A2 A3 B ZN VDD VSS 
MU14 ZN B VSS VSS n w=1u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=1u l=0.18u
MI20-M_u10 ZN A1 XI20-net17 VSS n w=1u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=1u l=0.18u
MU17 ZN A1 net19 VDD p w=1.37u l=0.18u
MU18 ZN A3 net19 VDD p w=1.37u l=0.18u
MU16 ZN A2 net19 VDD p w=1.37u l=0.18u
MU20 net19 B VDD VDD p w=1.37u l=0.18u
.ends
.subckt AOI31D2BWP7T A1 A2 A3 B ZN VDD VSS 
MU14 ZN B VSS VSS n w=2u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=1u l=0.18u
MI20-M_u10 ZN A1 XI20-net17 VSS n w=0.845u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=0.845u l=0.18u
MI7-MI12 XI7-net13 A3 VSS VSS n w=0.88u l=0.18u
MI7-M_u10 ZN A1 XI7-net17 VSS n w=0.88u l=0.18u
MI7-M_u11 XI7-net17 A2 XI7-net13 VSS n w=0.88u l=0.18u
MI6 ZN A1 net19 VDD p w=2.6u l=0.18u
MI4 ZN A3 net19 VDD p w=2.6u l=0.18u
MI5 ZN A2 net19 VDD p w=2.6u l=0.18u
MU20 net19 B VDD VDD p w=2.6u l=0.18u
.ends
.subckt AOI32D0BWP7T A1 A2 A3 B1 B2 ZN VDD VSS 
MI17-M_u10 ZN B1 XI17-net17 VSS n w=0.5u l=0.18u
MI17-M_u11 XI17-net17 B2 VSS VSS n w=0.5u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=0.5u l=0.18u
MI20-M_u10 ZN A1 XI20-net17 VSS n w=0.5u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=0.5u l=0.18u
MI4 ZN A1 net23 VDD p w=0.685u l=0.18u
MI2 ZN A3 net23 VDD p w=0.685u l=0.18u
MI3 ZN A2 net23 VDD p w=0.685u l=0.18u
MU20 net23 B1 VDD VDD p w=0.685u l=0.18u
MI1 net23 B2 VDD VDD p w=0.685u l=0.18u
.ends
.subckt AOI32D1BWP7T A1 A2 A3 B1 B2 ZN VDD VSS 
MI17-M_u10 ZN B1 XI17-net17 VSS n w=1u l=0.18u
MI17-M_u11 XI17-net17 B2 VSS VSS n w=1u l=0.18u
MI20-MI12 XI20-net13 A3 VSS VSS n w=1u l=0.18u
MI20-M_u10 ZN A1 XI20-net17 VSS n w=1u l=0.18u
MI20-M_u11 XI20-net17 A2 XI20-net13 VSS n w=1u l=0.18u
MU17 ZN A1 net23 VDD p w=1.37u l=0.18u
MU18 ZN A3 net23 VDD p w=1.37u l=0.18u
MU16 ZN A2 net23 VDD p w=1.37u l=0.18u
MU20 net23 B1 VDD VDD p w=1.37u l=0.18u
MU19 net23 B2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt AOI32D2BWP7T A1 A2 A3 B1 B2 ZN VDD VSS 
MI17_0-M_u10 ZN B1 XI17_0-net17 VSS n w=1u l=0.18u
MI17_0-M_u11 XI17_0-net17 B2 VSS VSS n w=1u l=0.18u
MI17_1-M_u10 ZN B1 XI17_1-net17 VSS n w=1u l=0.18u
MI17_1-M_u11 XI17_1-net17 B2 VSS VSS n w=1u l=0.18u
MI20_0-MI12 XI20_0-net13 A3 VSS VSS n w=0.905u l=0.18u
MI20_0-M_u10 ZN A1 XI20_0-net17 VSS n w=0.905u l=0.18u
MI20_0-M_u11 XI20_0-net17 A2 XI20_0-net13 VSS n w=0.905u l=0.18u
MI20_1-MI12 XI20_1-net13 A3 VSS VSS n w=0.905u l=0.18u
MI20_1-M_u10 ZN A1 XI20_1-net17 VSS n w=0.905u l=0.18u
MI20_1-M_u11 XI20_1-net17 A2 XI20_1-net13 VSS n w=0.905u l=0.18u
MI8 ZN A1 net23 VDD p w=2.55u l=0.18u
MI6 ZN A3 net23 VDD p w=2.55u l=0.18u
MI7 ZN A2 net23 VDD p w=2.55u l=0.18u
MU20 net23 B1 VDD VDD p w=2.74u l=0.18u
MI5 net23 B2 VDD VDD p w=2.74u l=0.18u
.ends
.subckt AOI33D0BWP7T A1 A2 A3 B1 B2 B3 ZN VDD VSS 
MI14-MI12 XI14-net13 A3 VSS VSS n w=0.5u l=0.18u
MI14-M_u10 ZN A1 XI14-net17 VSS n w=0.5u l=0.18u
MI14-M_u11 XI14-net17 A2 XI14-net13 VSS n w=0.5u l=0.18u
MI7-MI12 XI7-net13 B3 VSS VSS n w=0.5u l=0.18u
MI7-M_u10 ZN B1 XI7-net17 VSS n w=0.5u l=0.18u
MI7-M_u11 XI7-net17 B2 XI7-net13 VSS n w=0.5u l=0.18u
MI6 net40 A1 ZN VDD p w=0.685u l=0.18u
M_u16 VDD B3 net40 VDD p w=0.685u l=0.18u
MI3 VDD B1 net40 VDD p w=0.685u l=0.18u
MI4 net40 A3 ZN VDD p w=0.685u l=0.18u
MI5 net40 A2 ZN VDD p w=0.685u l=0.18u
MI2 VDD B2 net40 VDD p w=0.685u l=0.18u
.ends
.subckt AOI33D1BWP7T A1 A2 A3 B1 B2 B3 ZN VDD VSS 
MI14-MI12 XI14-net13 A3 VSS VSS n w=1u l=0.18u
MI14-M_u10 ZN A1 XI14-net17 VSS n w=1u l=0.18u
MI14-M_u11 XI14-net17 A2 XI14-net13 VSS n w=1u l=0.18u
MI2-MI12 XI2-net13 B3 VSS VSS n w=1u l=0.18u
MI2-M_u10 ZN B1 XI2-net17 VSS n w=1u l=0.18u
MI2-M_u11 XI2-net17 B2 XI2-net13 VSS n w=1u l=0.18u
M_u16 VDD B3 net40 VDD p w=1.37u l=0.18u
M_u15 VDD B2 net40 VDD p w=1.37u l=0.18u
M_u13 net40 A3 ZN VDD p w=1.37u l=0.18u
M_u12 net40 A2 ZN VDD p w=1.37u l=0.18u
M_u11 net40 A1 ZN VDD p w=1.37u l=0.18u
M_u14 VDD B1 net40 VDD p w=1.37u l=0.18u
.ends
.subckt AOI33D2BWP7T A1 A2 A3 B1 B2 B3 ZN VDD VSS 
MI9_0-MI12 XI9_0-net13 A3 VSS VSS n w=0.95u l=0.18u
MI9_0-M_u10 ZN A1 XI9_0-net17 VSS n w=0.95u l=0.18u
MI9_0-M_u11 XI9_0-net17 A2 XI9_0-net13 VSS n w=0.95u l=0.18u
MI9_1-MI12 XI9_1-net13 A3 VSS VSS n w=0.95u l=0.18u
MI9_1-M_u10 ZN A1 XI9_1-net17 VSS n w=0.95u l=0.18u
MI9_1-M_u11 XI9_1-net17 A2 XI9_1-net13 VSS n w=0.95u l=0.18u
MI2_0-MI12 XI2_0-net13 B3 VSS VSS n w=0.95u l=0.18u
MI2_0-M_u10 ZN B1 XI2_0-net17 VSS n w=0.95u l=0.18u
MI2_0-M_u11 XI2_0-net17 B2 XI2_0-net13 VSS n w=0.95u l=0.18u
MI2_1-MI12 XI2_1-net13 B3 VSS VSS n w=0.95u l=0.18u
MI2_1-M_u10 ZN B1 XI2_1-net17 VSS n w=0.95u l=0.18u
MI2_1-M_u11 XI2_1-net17 B2 XI2_1-net13 VSS n w=0.95u l=0.18u
MI7 net40 A1 ZN VDD p w=2.46u l=0.18u
M_u16 VDD B3 net40 VDD p w=2.46u l=0.18u
MI4 VDD B1 net40 VDD p w=2.46u l=0.18u
MI5 net40 A3 ZN VDD p w=2.46u l=0.18u
MI6 net40 A2 ZN VDD p w=2.46u l=0.18u
MI3 VDD B2 net40 VDD p w=2.46u l=0.18u
.ends
.subckt BHDBWP7T Z VDD VSS 
MU11 Z net8 VSS VSS n w=0.42u l=0.68u
M_u3 net8 Z VSS VSS n w=0.5u l=0.18u
MU12 Z net8 VDD VDD p w=0.42u l=0.68u
M_u7 net8 Z VDD VDD p w=0.685u l=0.18u
.ends
.subckt BUFFD0BWP7T I Z VDD VSS 
MI1-M_u2 Z net6 VSS VSS n w=0.5u l=0.18u
MI2-M_u2 net6 I VSS VSS n w=0.5u l=0.18u
MI1-M_u3 Z net6 VDD VDD p w=0.685u l=0.18u
MI2-M_u3 net6 I VDD VDD p w=0.685u l=0.18u
.ends
.subckt BUFFD10BWP7T I Z VDD VSS 
MI6-M_u2 n0 I VSS VSS n w=0.465u l=0.18u
MU8_0-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_1-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_2-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_3-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_4-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_5-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_6-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_7-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_8-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_9-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u2_0-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u2_1-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u2_2-M_u2 n0 I VSS VSS n w=1u l=0.18u
MI6-M_u3 n0 I VDD VDD p w=0.835u l=0.18u
MU8_0-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_1-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_2-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_3-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_4-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_5-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_6-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_7-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_8-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_9-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u2_0-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u2_1-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u2_2-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
.ends
.subckt BUFFD12BWP7T I Z VDD VSS 
MU8_0-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_1-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_2-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_3-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_4-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_5-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_6-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_7-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_8-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_9-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_10-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_11-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u2_0-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u2_1-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u2_2-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u2_3-M_u2 n0 I VSS VSS n w=1u l=0.18u
MU8_0-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_1-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_2-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_3-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_4-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_5-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_6-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_7-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_8-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_9-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_10-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_11-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u2_0-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u2_1-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u2_2-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u2_3-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
.ends
.subckt BUFFD1BWP7T I Z VDD VSS 
MI1-M_u2 Z net6 VSS VSS n w=1u l=0.18u
MI2-M_u2 net6 I VSS VSS n w=0.5u l=0.18u
MI1-M_u3 Z net6 VDD VDD p w=1.37u l=0.18u
MI2-M_u3 net6 I VDD VDD p w=0.685u l=0.18u
.ends
.subckt BUFFD1P5BWP7T I Z VDD VSS 
M_u3-M_u2 Z net8 VSS VSS n w=1.465u l=0.18u
M_u2-M_u2 net8 I VSS VSS n w=1u l=0.18u
M_u3-M_u3 Z net8 VDD VDD p w=2.055u l=0.18u
M_u2-M_u3 net8 I VDD VDD p w=1.37u l=0.18u
.ends
.subckt BUFFD2BWP7T I Z VDD VSS 
M_u2-M_u2 net8 I VSS VSS n w=1u l=0.18u
M_u3_0-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u2-M_u3 net8 I VDD VDD p w=1.37u l=0.18u
M_u3_0-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
.ends
.subckt BUFFD2P5BWP7T I Z VDD VSS 
M_u2-M_u2 net8 I VSS VSS n w=1u l=0.18u
M_u3-M_u2 Z net8 VSS VSS n w=2.5u l=0.18u
M_u2-M_u3 net8 I VDD VDD p w=1.37u l=0.18u
M_u3-M_u3 Z net8 VDD VDD p w=3.425u l=0.18u
.ends
.subckt BUFFD3BWP7T I Z VDD VSS 
M_u3_0-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_2-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u2-M_u2 net8 I VSS VSS n w=1u l=0.18u
M_u3_0-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_2-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u2-M_u3 net8 I VDD VDD p w=1.37u l=0.18u
.ends
.subckt BUFFD4BWP7T I Z VDD VSS 
M_u3_0-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_2-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_3-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u2_0-M_u2 p0 I VSS VSS n w=1u l=0.18u
M_u2_1-M_u2 p0 I VSS VSS n w=1u l=0.18u
M_u3_0-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_2-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_3-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u2_0-M_u3 p0 I VDD VDD p w=1.37u l=0.18u
M_u2_1-M_u3 p0 I VDD VDD p w=1.37u l=0.18u
.ends
.subckt BUFFD5BWP7T I Z VDD VSS 
MU8_0-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_1-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_2-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_3-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU8_4-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u2-M_u2 n0 I VSS VSS n w=2u l=0.18u
MU8_0-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_1-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_2-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_3-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU8_4-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u2-M_u3 n0 I VDD VDD p w=2.74u l=0.18u
.ends
.subckt BUFFD6BWP7T I Z VDD VSS 
M_u3_0-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_2-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_3-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_4-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_5-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u2-M_u2 net8 I VSS VSS n w=2u l=0.18u
M_u3_0-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_2-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_3-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_4-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_5-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u2-M_u3 net8 I VDD VDD p w=2.74u l=0.18u
.ends
.subckt BUFFD8BWP7T I Z VDD VSS 
M_u2_0-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u2_1-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u2_2-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u7_0-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_1-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_2-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_3-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_4-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_5-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_6-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_7-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u2_0-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u2_1-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u2_2-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u7_0-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_1-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_2-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_3-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_4-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_5-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_6-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_7-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
.ends
.subckt BUFTD0BWP7T I OE Z VDD VSS 
M_u17-M_u2 net31 OE VSS VSS n w=0.5u l=0.18u
M_u7 Z INEN VSS VSS n w=0.5u l=0.18u
MU19-M_u4 INEN I VSS VSS n w=0.5u l=0.18u
MU19-M_u3 INEN net31 VSS VSS n w=0.5u l=0.18u
MU18-M_u4 XU18-net6 I VSS VSS n w=0.5u l=0.18u
MU18-M_u3 INEP OE XU18-net6 VSS n w=0.5u l=0.18u
M_u17-M_u3 net31 OE VDD VDD p w=0.685u l=0.18u
MU19-M_u1 XU19-net8 net31 VDD VDD p w=0.685u l=0.18u
MU19-M_u2 INEN I XU19-net8 VDD p w=0.685u l=0.18u
MU18-M_u2 INEP I VDD VDD p w=0.685u l=0.18u
MU18-M_u1 INEP OE VDD VDD p w=0.685u l=0.18u
M_u6 Z INEP VDD VDD p w=0.685u l=0.18u
.ends
.subckt BUFTD1BWP7T I OE Z VDD VSS 
M_u17-M_u2 net31 OE VSS VSS n w=0.5u l=0.18u
M_u7 Z INEN VSS VSS n w=0.7u l=0.18u
MU19-M_u4 INEN I VSS VSS n w=0.5u l=0.18u
MU19-M_u3 INEN net31 VSS VSS n w=0.5u l=0.18u
MU18-M_u4 XU18-net6 I VSS VSS n w=0.685u l=0.18u
MU18-M_u3 INEP OE XU18-net6 VSS n w=0.685u l=0.18u
M_u17-M_u3 net31 OE VDD VDD p w=0.685u l=0.18u
MU19-M_u1 XU19-net8 net31 VDD VDD p w=1.315u l=0.18u
MU19-M_u2 INEN I XU19-net8 VDD p w=1.315u l=0.18u
MU18-M_u2 INEP I VDD VDD p w=0.70u l=0.18u
MU18-M_u1 INEP OE VDD VDD p w=0.70u l=0.18u
M_u6 Z INEP VDD VDD p w=1.37u l=0.18u
.ends
.subckt BUFTD2BWP7T I OE Z VDD VSS 
M_u17-M_u2 net31 OE VSS VSS n w=0.5u l=0.18u
M_u7 Z INEN VSS VSS n w=1.63u l=0.18u
MU19-M_u4 INEN I VSS VSS n w=0.5u l=0.18u
MU19-M_u3 INEN net31 VSS VSS n w=0.5u l=0.18u
MU18-M_u4 XU18-net6 I VSS VSS n w=0.685u l=0.18u
MU18-M_u3 INEP OE XU18-net6 VSS n w=0.685u l=0.18u
M_u17-M_u3 net31 OE VDD VDD p w=0.685u l=0.18u
MU19-M_u1 XU19-net8 net31 VDD VDD p w=1.23u l=0.18u
MU19-M_u2 INEN I XU19-net8 VDD p w=1.23u l=0.18u
MU18-M_u2 INEP I VDD VDD p w=0.65u l=0.18u
MU18-M_u1 INEP OE VDD VDD p w=0.65u l=0.18u
M_u6 Z INEP VDD VDD p w=2.37u l=0.18u
.ends
.subckt BUFTD3BWP7T I OE Z VDD VSS 
M_u17-M_u2 net31 OE VSS VSS n w=0.5u l=0.18u
M_u7 Z INEN VSS VSS n w=2.43u l=0.18u
MU19-M_u4 INEN I VSS VSS n w=0.5u l=0.18u
MU19-M_u3 INEN net31 VSS VSS n w=0.5u l=0.18u
MU18-M_u4 XU18-net6 I VSS VSS n w=0.685u l=0.18u
MU18-M_u3 INEP OE XU18-net6 VSS n w=0.685u l=0.18u
M_u17-M_u3 net31 OE VDD VDD p w=0.685u l=0.18u
MU19-M_u1 XU19-net8 net31 VDD VDD p w=1.23u l=0.18u
MU19-M_u2 INEN I XU19-net8 VDD p w=1.23u l=0.18u
MU18-M_u2 INEP I VDD VDD p w=0.685u l=0.18u
MU18-M_u1 INEP OE VDD VDD p w=0.685u l=0.18u
M_u6 Z INEP VDD VDD p w=3.585u l=0.18u
.ends
.subckt BUFTD4BWP7T I OE Z VDD VSS 
M_u17-M_u2 net31 OE VSS VSS n w=0.5u l=0.18u
M_u7 Z INEN VSS VSS n w=3.26u l=0.18u
MU19-M_u4 INEN I VSS VSS n w=0.5u l=0.18u
MU19-M_u3 INEN net31 VSS VSS n w=0.5u l=0.18u
MU18-M_u4 XU18-net6 I VSS VSS n w=0.685u l=0.18u
MU18-M_u3 INEP OE XU18-net6 VSS n w=0.685u l=0.18u
M_u17-M_u3 net31 OE VDD VDD p w=0.685u l=0.18u
MU19-M_u1 XU19-net8 net31 VDD VDD p w=1.23u l=0.18u
MU19-M_u2 INEN I XU19-net8 VDD p w=1.23u l=0.18u
MU18-M_u2 INEP I VDD VDD p w=0.685u l=0.18u
MU18-M_u1 INEP OE VDD VDD p w=0.685u l=0.18u
M_u6 Z INEP VDD VDD p w=4.78u l=0.18u
.ends
.subckt BUFTD6BWP7T I OE Z VDD VSS 
MI5_0-M_u4 INEN net13 VSS VSS n w=0.73u l=0.18u
MI5_0-M_u3 INEN I VSS VSS n w=0.73u l=0.18u
MI5_1-M_u4 INEN net13 VSS VSS n w=0.73u l=0.18u
MI5_1-M_u3 INEN I VSS VSS n w=0.73u l=0.18u
M_u17-M_u2 net13 OE VSS VSS n w=0.5u l=0.18u
M_u7 Z INEN VSS VSS n w=5.01u l=0.18u
MI7_0-M_u4 XI7_0-net6 I VSS VSS n w=0.57u l=0.18u
MI7_0-M_u3 INEP OE XI7_0-net6 VSS n w=0.57u l=0.18u
MI7_1-M_u4 XI7_1-net6 I VSS VSS n w=0.57u l=0.18u
MI7_1-M_u3 INEP OE XI7_1-net6 VSS n w=0.57u l=0.18u
MI5_0-M_u1 XI5_0-net8 I VDD VDD p w=1.035u l=0.18u
MI5_0-M_u2 INEN net13 XI5_0-net8 VDD p w=1.035u l=0.18u
MI5_1-M_u1 XI5_1-net8 I VDD VDD p w=1.035u l=0.18u
MI5_1-M_u2 INEN net13 XI5_1-net8 VDD p w=1.035u l=0.18u
M_u17-M_u3 net13 OE VDD VDD p w=0.685u l=0.18u
MI7_0-M_u2 INEP I VDD VDD p w=0.88u l=0.18u
MI7_0-M_u1 INEP OE VDD VDD p w=0.88u l=0.18u
MI7_1-M_u2 INEP I VDD VDD p w=0.88u l=0.18u
MI7_1-M_u1 INEP OE VDD VDD p w=0.88u l=0.18u
M_u6 Z INEP VDD VDD p w=7.59u l=0.18u
.ends
.subckt BUFTD8BWP7T I OE Z VDD VSS 
MI5_0-M_u4 INEN net31 VSS VSS n w=0.73u l=0.18u
MI5_0-M_u3 INEN I VSS VSS n w=0.73u l=0.18u
MI5_1-M_u4 INEN net31 VSS VSS n w=0.73u l=0.18u
MI5_1-M_u3 INEN I VSS VSS n w=0.73u l=0.18u
M_u17-M_u2 net31 OE VSS VSS n w=0.5u l=0.18u
M_u7 Z INEN VSS VSS n w=6.68u l=0.18u
MI7_0-M_u4 XI7_0-net6 I VSS VSS n w=0.57u l=0.18u
MI7_0-M_u3 INEP OE XI7_0-net6 VSS n w=0.57u l=0.18u
MI7_1-M_u4 XI7_1-net6 I VSS VSS n w=0.57u l=0.18u
MI7_1-M_u3 INEP OE XI7_1-net6 VSS n w=0.57u l=0.18u
MI5_0-M_u1 XI5_0-net8 I VDD VDD p w=1.035u l=0.18u
MI5_0-M_u2 INEN net31 XI5_0-net8 VDD p w=1.035u l=0.18u
MI5_1-M_u1 XI5_1-net8 I VDD VDD p w=1.035u l=0.18u
MI5_1-M_u2 INEN net31 XI5_1-net8 VDD p w=1.035u l=0.18u
M_u17-M_u3 net31 OE VDD VDD p w=0.685u l=0.18u
MI7_0-M_u2 INEP I VDD VDD p w=0.88u l=0.18u
MI7_0-M_u1 INEP OE VDD VDD p w=0.88u l=0.18u
MI7_1-M_u2 INEP I VDD VDD p w=0.88u l=0.18u
MI7_1-M_u1 INEP OE VDD VDD p w=0.88u l=0.18u
M_u6 Z INEP VDD VDD p w=10.12u l=0.18u
.ends
.subckt CKAN2D0BWP7T A1 A2 Z VDD VSS 
MI10 net015 A2 VSS VSS n w=0.42u l=0.18u
MI11 net6 A1 net015 VSS n w=0.42u l=0.18u
M_u3-M_u2 Z net6 VSS VSS n w=0.42u l=0.18u
M_u3-M_u3 Z net6 VDD VDD p w=1.13u l=0.18u
MI2 net6 A2 VDD VDD p w=0.755u l=0.18u
MI1 VDD A1 net6 VDD p w=0.71u l=0.18u
.ends
.subckt CKAN2D1BWP7T A1 A2 Z VDD VSS 
M_u7 net6 A1 net012 VSS n w=0.5u l=0.18u
MI7 net012 A2 VSS VSS n w=0.5u l=0.18u
M_u3-M_u2 Z net6 VSS VSS n w=0.525u l=0.18u
M_u3-M_u3 Z net6 VDD VDD p w=1.37u l=0.18u
MI1 VDD A1 net6 VDD p w=0.85u l=0.18u
MI2 net6 A2 VDD VDD p w=0.9u l=0.18u
.ends
.subckt CKAN2D2BWP7T A1 A2 Z VDD VSS 
M_u7 net017 A1 net015 VSS n w=0.74u l=0.18u
MI7 net015 A2 VSS VSS n w=0.74u l=0.18u
M_u3_0-M_u2 Z net017 VSS VSS n w=0.525u l=0.18u
M_u3_1-M_u2 Z net017 VSS VSS n w=0.525u l=0.18u
M_u3_0-M_u3 Z net017 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z net017 VDD VDD p w=1.37u l=0.18u
MI1 VDD A1 net017 VDD p w=1.23u l=0.18u
MI2 net017 A2 VDD VDD p w=1.29u l=0.18u
.ends
.subckt CKAN2D4BWP7T A1 A2 Z VDD VSS 
MI7 net16 A2 VSS VSS n w=1.08u l=0.18u
M_u7 net28 A1 net16 VSS n w=1.08u l=0.18u
M_u3_0-M_u2 Z net28 VSS VSS n w=0.525u l=0.18u
M_u3_1-M_u2 Z net28 VSS VSS n w=0.525u l=0.18u
M_u3_2-M_u2 Z net28 VSS VSS n w=0.525u l=0.18u
M_u3_3-M_u2 Z net28 VSS VSS n w=0.525u l=0.18u
M_u3_0-M_u3 Z net28 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z net28 VDD VDD p w=1.37u l=0.18u
M_u3_2-M_u3 Z net28 VDD VDD p w=1.37u l=0.18u
M_u3_3-M_u3 Z net28 VDD VDD p w=1.37u l=0.18u
MI2 net28 A2 VDD VDD p w=2.19u l=0.18u
MI1 VDD A1 net28 VDD p w=2.19u l=0.18u
.ends
.subckt CKAN2D8BWP7T A1 A2 Z VDD VSS 
MI7_0 n1 A2 VSS VSS n w=0.67u l=0.18u
MI7_1 n1 A2 VSS VSS n w=0.67u l=0.18u
MI7_2 n1 A2 VSS VSS n w=0.67u l=0.18u
M_u7_0 n0 A1 n1 VSS n w=0.67u l=0.18u
M_u7_1 n0 A1 n1 VSS n w=0.67u l=0.18u
M_u7_2 n0 A1 n1 VSS n w=0.67u l=0.18u
M_u3-M_u2 Z n0 VSS VSS n w=4.2u l=0.18u
M_u3-M_u3 Z n0 VDD VDD p w=10.94u l=0.18u
MI2_0 n0 A2 VDD VDD p w=1.37u l=0.18u
MI2_1 n0 A2 VDD VDD p w=1.37u l=0.18u
MI2_2 n0 A2 VDD VDD p w=1.37u l=0.18u
MI1_0 VDD A1 n0 VDD p w=1.32u l=0.18u
MI1_1 VDD A1 n0 VDD p w=1.32u l=0.18u
MI1_2 VDD A1 n0 VDD p w=1.32u l=0.18u
.ends
.subckt CKBD0BWP7T I Z VDD VSS 
MU23 Z net21 VSS VSS n w=0.42u l=0.18u
M_u15 net21 I VSS VSS n w=0.42u l=0.18u
MU21 Z net21 VDD VDD p w=1.13u l=0.18u
M_u3 net21 I VDD VDD p w=1.27u l=0.18u
.ends
.subckt CKBD10BWP7T I Z VDD VSS 
DI3 VSS I dn 0.2037p
MU23 Z net25 VSS VSS n w=5.49u l=0.18u
M_u15 net25 I VSS VSS n w=2.35u l=0.18u
MU21 Z net25 VDD VDD p w=13.69u l=0.18u
M_u3 net25 I VDD VDD p w=7.05u l=0.18u
.ends
.subckt CKBD12BWP7T I Z VDD VSS 
DI3 VSS I dn 0.2037p
MU23 Z N1 VSS VSS n w=6.595u l=0.18u
M_u15_0 N1 I VSS VSS n w=0.59u l=0.18u
M_u15_1 N1 I VSS VSS n w=0.59u l=0.18u
M_u15_2 N1 I VSS VSS n w=0.59u l=0.18u
M_u15_3 N1 I VSS VSS n w=0.59u l=0.18u
M_u15_4 N1 I VSS VSS n w=0.59u l=0.18u
MU21 Z N1 VDD VDD p w=15.06u l=0.18u
M_u3 N1 I VDD VDD p w=8.1u l=0.18u
.ends
.subckt CKBD1BWP7T I Z VDD VSS 
MU23 Z net21 VSS VSS n w=0.52u l=0.18u
M_u15 net21 I VSS VSS n w=0.455u l=0.18u
MU21 Z net21 VDD VDD p w=1.37u l=0.18u
M_u3 net21 I VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKBD2BWP7T I Z VDD VSS 
MU23_0 Z net025 VSS VSS n w=0.525u l=0.18u
MU23_1 Z net025 VSS VSS n w=0.525u l=0.18u
M_u15 net025 I VSS VSS n w=0.525u l=0.18u
MU21_0 Z net025 VDD VDD p w=1.37u l=0.18u
MU21_1 Z net025 VDD VDD p w=1.37u l=0.18u
M_u3 net025 I VDD VDD p w=1.54u l=0.18u
.ends
.subckt CKBD3BWP7T I Z VDD VSS 
DI3 VSS I dn 0.2037p
MU23_0 Z net28 VSS VSS n w=0.83u l=0.18u
MU23_1 Z net28 VSS VSS n w=0.83u l=0.18u
M_u15 net28 I VSS VSS n w=0.8u l=0.18u
MU21 Z net28 VDD VDD p w=4.11u l=0.18u
M_u3_0 net28 I VDD VDD p w=1.14u l=0.18u
M_u3_1 net28 I VDD VDD p w=1.14u l=0.18u
.ends
.subckt CKBD4BWP7T I Z VDD VSS 
DI3 VSS I dn 0.2037p
MU23 Z net23 VSS VSS n w=2.19u l=0.18u
M_u15_0 net23 I VSS VSS n w=0.455u l=0.18u
M_u15_1 net23 I VSS VSS n w=0.455u l=0.18u
MU21_0 Z net23 VDD VDD p w=1.37u l=0.18u
MU21_1 Z net23 VDD VDD p w=1.37u l=0.18u
MU21_2 Z net23 VDD VDD p w=1.37u l=0.18u
MU21_3 Z net23 VDD VDD p w=1.37u l=0.18u
M_u3_0 net23 I VDD VDD p w=1.37u l=0.18u
M_u3_1 net23 I VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKBD6BWP7T I Z VDD VSS 
DI3 VSS I dn 0.2037p
MU23 Z net25 VSS VSS n w=3.225u l=0.18u
M_u15_0 net25 I VSS VSS n w=0.72u l=0.18u
M_u15_1 net25 I VSS VSS n w=0.72u l=0.18u
MU21_0 Z net25 VDD VDD p w=1.37u l=0.18u
MU21_1 Z net25 VDD VDD p w=1.37u l=0.18u
MU21_2 Z net25 VDD VDD p w=1.37u l=0.18u
MU21_3 Z net25 VDD VDD p w=1.37u l=0.18u
MU21_4 Z net25 VDD VDD p w=1.37u l=0.18u
MU21_5 Z net25 VDD VDD p w=1.37u l=0.18u
M_u3_0 net25 I VDD VDD p w=1.37u l=0.18u
M_u3_1 net25 I VDD VDD p w=1.37u l=0.18u
M_u3_2 net25 I VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKBD8BWP7T I Z VDD VSS 
DI3 VSS I dn 0.2037p
MU23_0 Z net28 VSS VSS n w=0.62u l=0.18u
MU23_1 Z net28 VSS VSS n w=0.62u l=0.18u
MU23_2 Z net28 VSS VSS n w=0.62u l=0.18u
MU23_3 Z net28 VSS VSS n w=0.62u l=0.18u
MU23_4 Z net28 VSS VSS n w=0.62u l=0.18u
MU23_5 Z net28 VSS VSS n w=0.62u l=0.18u
M_u15 net28 I VSS VSS n w=1.66u l=0.18u
MU21 Z net28 VDD VDD p w=9.59u l=0.18u
M_u3 net28 I VDD VDD p w=5.11u l=0.18u
.ends
.subckt CKLHQD1BWP7T  Q TE CPN E VDD VSS 
MU19 net50 E VSS VSS n w=0.42u l=0.18u
MU20 net50 TE VSS VSS n w=0.42u l=0.18u
MI82 net53 INCP net50 VSS n w=0.42u l=0.18u
MI89-M_u2 net36 QD VSS VSS n w=0.505u l=0.18u
MI80-M_u2 QD net53 VSS VSS n w=0.5u l=0.18u
MU75-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MU82-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MU81-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI1-M_u4 d3 CPN VSS VSS n w=0.42u l=0.18u
MI1-M_u3 d3 net36 VSS VSS n w=0.42u l=0.18u
MI79-MU3 net53 INCPB XI79-net16 VSS n w=0.42u l=0.18u
MI79-MU4 XI79-net16 QD VSS VSS n w=0.42u l=0.18u
MI89-M_u3 net36 QD VDD VDD p w=0.685u l=0.18u
MI80-M_u3 QD net53 VDD VDD p w=0.62u l=0.18u
MU75-M_u3 Q d3 VDD VDD p w=1.27u l=0.18u
MU82-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MU81-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI1-M_u1 XI1-net8 net36 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 d3 CPN XI1-net8 VDD p w=1.37u l=0.18u
MU16 net53 INCPB net61 VDD p w=0.52u l=0.18u
MU17 net61 E net58 VDD p w=1.37u l=0.18u
MI81 net58 TE VDD VDD p w=1.37u l=0.18u
MI79-MU2 net53 INCP XI79-net6 VDD p w=0.42u l=0.18u
MI79-MU1 XI79-net6 QD VDD VDD p w=0.42u l=0.18u
.ends
.subckt CKLHQD2BWP7T  Q TE CPN E VDD VSS 
MU19 net50 E VSS VSS n w=0.42u l=0.18u
MU20 net50 TE VSS VSS n w=0.42u l=0.18u
MI82 net53 INCP net50 VSS n w=0.42u l=0.18u
MI1-M_u4 net38 CPN VSS VSS n w=0.42u l=0.18u
MI1-M_u3 net38 net36 VSS VSS n w=0.42u l=0.18u
MI89-M_u2 net36 QD VSS VSS n w=0.505u l=0.18u
MI88-M_u2 Q net38 VSS VSS n w=2u l=0.18u
MI80-M_u2 QD net53 VSS VSS n w=0.5u l=0.18u
MU82-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MU81-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI79-MU3 net53 INCPB XI79-net16 VSS n w=0.42u l=0.18u
MI79-MU4 XI79-net16 QD VSS VSS n w=0.42u l=0.18u
MI1-M_u1 XI1-net8 net36 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 net38 CPN XI1-net8 VDD p w=1.37u l=0.18u
MI89-M_u3 net36 QD VDD VDD p w=0.685u l=0.18u
MI88-M_u3 Q net38 VDD VDD p w=2.2u l=0.18u
MI80-M_u3 QD net53 VDD VDD p w=0.62u l=0.18u
MU82-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MU81-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MU16 net53 INCPB net61 VDD p w=0.52u l=0.18u
MU17 net61 E net58 VDD p w=1.37u l=0.18u
MI81 net58 TE VDD VDD p w=1.37u l=0.18u
MI79-MU2 net53 INCP XI79-net6 VDD p w=0.42u l=0.18u
MI79-MU1 XI79-net6 QD VDD VDD p w=0.42u l=0.18u
.ends
.subckt CKLHQD4BWP7T  Q TE CPN E VDD VSS 
MU19 net50 E VSS VSS n w=0.42u l=0.18u
MU20 net50 TE VSS VSS n w=0.42u l=0.18u
MI82 net53 INCP net50 VSS n w=0.42u l=0.18u
MI89-M_u2 net85 QD VSS VSS n w=0.94u l=0.18u
MI80-M_u2 QD net53 VSS VSS n w=0.5u l=0.18u
MU75_0-M_u2 Q net52 VSS VSS n w=1u l=0.18u
MU75_1-M_u2 Q net52 VSS VSS n w=1u l=0.18u
MU75_2-M_u2 Q net52 VSS VSS n w=1u l=0.18u
MU75_3-M_u2 Q net52 VSS VSS n w=1u l=0.18u
MU82-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MU81-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI1-M_u4 net52 CPN VSS VSS n w=0.49u l=0.18u
MI1-M_u3 net52 net85 VSS VSS n w=0.49u l=0.18u
MI90-M_u4 net52 CPN VSS VSS n w=0.49u l=0.18u
MI90-M_u3 net52 net85 VSS VSS n w=0.49u l=0.18u
MI79-MU3 net53 INCPB XI79-net16 VSS n w=0.42u l=0.18u
MI79-MU4 XI79-net16 QD VSS VSS n w=0.42u l=0.18u
MU16 net53 INCPB net61 VDD p w=0.52u l=0.18u
MU17 net61 E net58 VDD p w=1.37u l=0.18u
MI81 net58 TE VDD VDD p w=1.37u l=0.18u
MI89-M_u3 net85 QD VDD VDD p w=1.33u l=0.18u
MI80-M_u3 QD net53 VDD VDD p w=0.62u l=0.18u
MU75_0-M_u3 Q net52 VDD VDD p w=0.98u l=0.18u
MU75_1-M_u3 Q net52 VDD VDD p w=0.98u l=0.18u
MU75_2-M_u3 Q net52 VDD VDD p w=0.98u l=0.18u
MU75_3-M_u3 Q net52 VDD VDD p w=0.98u l=0.18u
MU82-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MU81-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI1-M_u1 XI1-net8 net85 VDD VDD p w=1.33u l=0.18u
MI1-M_u2 net52 CPN XI1-net8 VDD p w=1.33u l=0.18u
MI90-M_u1 XI90-net8 net85 VDD VDD p w=1.33u l=0.18u
MI90-M_u2 net52 CPN XI90-net8 VDD p w=1.33u l=0.18u
MI79-MU2 net53 INCP XI79-net6 VDD p w=0.42u l=0.18u
MI79-MU1 XI79-net6 QD VDD VDD p w=0.42u l=0.18u
.ends
.subckt CKLHQD6BWP7T  Q TE CPN E VDD VSS 
MU19 net50 E VSS VSS n w=0.42u l=0.18u
MU20 net50 TE VSS VSS n w=0.42u l=0.18u
MI82 net53 INCP net50 VSS n w=0.42u l=0.18u
MI89-M_u2 net85 QD VSS VSS n w=0.94u l=0.18u
MI80-M_u2 QD net53 VSS VSS n w=0.5u l=0.18u
MU75_0-M_u2 Q net52 VSS VSS n w=1u l=0.18u
MU75_1-M_u2 Q net52 VSS VSS n w=1u l=0.18u
MU75_2-M_u2 Q net52 VSS VSS n w=1u l=0.18u
MU75_3-M_u2 Q net52 VSS VSS n w=1u l=0.18u
MU75_4-M_u2 Q net52 VSS VSS n w=1u l=0.18u
MU75_5-M_u2 Q net52 VSS VSS n w=1u l=0.18u
MU82-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MU81-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI1-M_u4 net52 CPN VSS VSS n w=0.49u l=0.18u
MI1-M_u3 net52 net85 VSS VSS n w=0.49u l=0.18u
MI90-M_u4 net52 CPN VSS VSS n w=0.49u l=0.18u
MI90-M_u3 net52 net85 VSS VSS n w=0.49u l=0.18u
MI79-MU3 net53 INCPB XI79-net16 VSS n w=0.42u l=0.18u
MI79-MU4 XI79-net16 QD VSS VSS n w=0.42u l=0.18u
MI89-M_u3 net85 QD VDD VDD p w=1.37u l=0.18u
MI80-M_u3 QD net53 VDD VDD p w=0.62u l=0.18u
MU75_0-M_u3 Q net52 VDD VDD p w=0.9u l=0.18u
MU75_1-M_u3 Q net52 VDD VDD p w=0.9u l=0.18u
MU75_2-M_u3 Q net52 VDD VDD p w=0.9u l=0.18u
MU75_3-M_u3 Q net52 VDD VDD p w=0.9u l=0.18u
MU75_4-M_u3 Q net52 VDD VDD p w=0.9u l=0.18u
MU75_5-M_u3 Q net52 VDD VDD p w=0.9u l=0.18u
MU82-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MU81-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI1-M_u1 XI1-net8 net85 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 net52 CPN XI1-net8 VDD p w=1.37u l=0.18u
MI90-M_u1 XI90-net8 net85 VDD VDD p w=1.37u l=0.18u
MI90-M_u2 net52 CPN XI90-net8 VDD p w=1.37u l=0.18u
MU16 net53 INCPB net61 VDD p w=0.52u l=0.18u
MU17 net61 E net58 VDD p w=1.37u l=0.18u
MI81 net58 TE VDD VDD p w=1.37u l=0.18u
MI79-MU2 net53 INCP XI79-net6 VDD p w=0.42u l=0.18u
MI79-MU1 XI79-net6 QD VDD VDD p w=0.42u l=0.18u
.ends
.subckt CKLHQD8BWP7T  Q TE CPN E VDD VSS 
MU19 net50 E VSS VSS n w=0.42u l=0.18u
MU20 net50 TE VSS VSS n w=0.42u l=0.18u
MI82 net53 INCP net50 VSS n w=0.42u l=0.18u
MI89-M_u2 net061 QD VSS VSS n w=0.94u l=0.18u
MI80-M_u2 QD net53 VSS VSS n w=0.5u l=0.18u
MU75_0-M_u2 Q net111 VSS VSS n w=1u l=0.18u
MU75_1-M_u2 Q net111 VSS VSS n w=1u l=0.18u
MU75_2-M_u2 Q net111 VSS VSS n w=1u l=0.18u
MU75_3-M_u2 Q net111 VSS VSS n w=1u l=0.18u
MU75_4-M_u2 Q net111 VSS VSS n w=1u l=0.18u
MU75_5-M_u2 Q net111 VSS VSS n w=1u l=0.18u
MU75_6-M_u2 Q net111 VSS VSS n w=1u l=0.18u
MU75_7-M_u2 Q net111 VSS VSS n w=1u l=0.18u
MU82-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MU81-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI1-M_u4 net111 CPN VSS VSS n w=0.49u l=0.18u
MI1-M_u3 net111 net061 VSS VSS n w=0.49u l=0.18u
MI95-M_u4 net111 CPN VSS VSS n w=0.49u l=0.18u
MI95-M_u3 net111 net061 VSS VSS n w=0.49u l=0.18u
MI79-MU3 net53 INCPB XI79-net16 VSS n w=0.42u l=0.18u
MI79-MU4 XI79-net16 QD VSS VSS n w=0.42u l=0.18u
MI89-M_u3 net061 QD VDD VDD p w=1.37u l=0.18u
MI80-M_u3 QD net53 VDD VDD p w=0.62u l=0.18u
MU75_0-M_u3 Q net111 VDD VDD p w=0.92u l=0.18u
MU75_1-M_u3 Q net111 VDD VDD p w=0.92u l=0.18u
MU75_2-M_u3 Q net111 VDD VDD p w=0.92u l=0.18u
MU75_3-M_u3 Q net111 VDD VDD p w=0.92u l=0.18u
MU75_4-M_u3 Q net111 VDD VDD p w=0.92u l=0.18u
MU75_5-M_u3 Q net111 VDD VDD p w=0.92u l=0.18u
MU75_6-M_u3 Q net111 VDD VDD p w=0.92u l=0.18u
MU75_7-M_u3 Q net111 VDD VDD p w=0.92u l=0.18u
MU82-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MU81-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI1-M_u1 XI1-net8 net061 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 net111 CPN XI1-net8 VDD p w=1.37u l=0.18u
MI95-M_u1 XI95-net8 net061 VDD VDD p w=1.37u l=0.18u
MI95-M_u2 net111 CPN XI95-net8 VDD p w=1.37u l=0.18u
MU16 net53 INCPB net61 VDD p w=0.52u l=0.18u
MU17 net61 E net58 VDD p w=1.37u l=0.18u
MI81 net58 TE VDD VDD p w=1.37u l=0.18u
MI79-MU2 net53 INCP XI79-net6 VDD p w=0.42u l=0.18u
MI79-MU1 XI79-net6 QD VDD VDD p w=0.42u l=0.18u
.ends
.subckt CKLNQD1BWP7T TE E CP Q VDD VSS 
MU19 net50 E VSS VSS n w=0.5u l=0.18u
MU20 net50 TE VSS VSS n w=0.5u l=0.18u
MI82 net53 INCPB net50 VSS n w=0.5u l=0.18u
MI80-M_u2 QD net53 VSS VSS n w=0.5u l=0.18u
MU75-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU82-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MU81-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI85-M_u4 XI85-net6 QD VSS VSS n w=0.5u l=0.18u
MI85-M_u3 d3 CP XI85-net6 VSS n w=0.5u l=0.18u
MI79-MU3 net53 INCP XI79-net16 VSS n w=0.42u l=0.18u
MI79-MU4 XI79-net16 QD VSS VSS n w=0.42u l=0.18u
MI80-M_u3 QD net53 VDD VDD p w=0.685u l=0.18u
MU75-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU82-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MU81-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI85-M_u2 d3 QD VDD VDD p w=0.85u l=0.18u
MI85-M_u1 d3 CP VDD VDD p w=0.9u l=0.18u
MU16 net53 INCP net61 VDD p w=0.52u l=0.18u
MU17 net61 E net58 VDD p w=1.37u l=0.18u
MI81 net58 TE VDD VDD p w=1.37u l=0.18u
MI79-MU2 net53 INCPB XI79-net6 VDD p w=0.42u l=0.18u
MI79-MU1 XI79-net6 QD VDD VDD p w=0.42u l=0.18u
.ends
.subckt CKLNQD2BWP7T TE E CP Q VDD VSS 
MU19 net50 E VSS VSS n w=0.5u l=0.18u
MU20 net50 TE VSS VSS n w=0.5u l=0.18u
MI82 net53 INCPB net50 VSS n w=0.5u l=0.18u
MI80-M_u2 QD net53 VSS VSS n w=0.5u l=0.18u
MU75_0-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU75_1-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU82-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MU81-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI85-M_u4 XI85-net6 QD VSS VSS n w=0.7u l=0.18u
MI85-M_u3 d3 CP XI85-net6 VSS n w=0.7u l=0.18u
MI79-MU3 net53 INCP XI79-net16 VSS n w=0.42u l=0.18u
MI79-MU4 XI79-net16 QD VSS VSS n w=0.42u l=0.18u
MI80-M_u3 QD net53 VDD VDD p w=0.685u l=0.18u
MU75_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU75_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU82-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MU81-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI85-M_u2 d3 QD VDD VDD p w=1.37u l=0.18u
MI85-M_u1 d3 CP VDD VDD p w=1.37u l=0.18u
MU16 net53 INCP net61 VDD p w=0.52u l=0.18u
MU17 net61 E net58 VDD p w=1.37u l=0.18u
MI81 net58 TE VDD VDD p w=1.37u l=0.18u
MI79-MU2 net53 INCPB XI79-net6 VDD p w=0.42u l=0.18u
MI79-MU1 XI79-net6 QD VDD VDD p w=0.42u l=0.18u
.ends
.subckt CKLNQD4BWP7T TE E CP Q VDD VSS 
MU19 net50 E VSS VSS n w=0.5u l=0.18u
MU20 net50 TE VSS VSS n w=0.5u l=0.18u
MI82 net53 INCPB net50 VSS n w=0.5u l=0.18u
MI80-M_u2 QD net53 VSS VSS n w=0.5u l=0.18u
MU75_0-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU75_1-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU75_2-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU75_3-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU82-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MU81-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI87-M_u4 XI87-net6 CP VSS VSS n w=1.08u l=0.18u
MI87-M_u3 d3 QD XI87-net6 VSS n w=1.08u l=0.18u
MI79-MU3 net53 INCP XI79-net16 VSS n w=0.42u l=0.18u
MI79-MU4 XI79-net16 QD VSS VSS n w=0.42u l=0.18u
MI80-M_u3 QD net53 VDD VDD p w=0.685u l=0.18u
MU75_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU75_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU75_2-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU75_3-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU82-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MU81-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI87-M_u2 d3 CP VDD VDD p w=2.19u l=0.18u
MI87-M_u1 d3 QD VDD VDD p w=2.19u l=0.18u
MU16 net53 INCP net61 VDD p w=0.52u l=0.18u
MU17 net61 E net58 VDD p w=1.37u l=0.18u
MI81 net58 TE VDD VDD p w=1.37u l=0.18u
MI79-MU2 net53 INCPB XI79-net6 VDD p w=0.42u l=0.18u
MI79-MU1 XI79-net6 QD VDD VDD p w=0.42u l=0.18u
.ends
.subckt CKLNQD6BWP7T TE E CP Q VDD VSS 
MU19 net50 E VSS VSS n w=0.5u l=0.18u
MU20 net50 TE VSS VSS n w=0.5u l=0.18u
MI82 net53 INCPB net50 VSS n w=0.5u l=0.18u
MI87-M_u4 XI87-net6 QD VSS VSS n w=1.62u l=0.18u
MI87-M_u3 d3 CP XI87-net6 VSS n w=1.62u l=0.18u
MI80-M_u2 QD net53 VSS VSS n w=0.5u l=0.18u
MU75_0-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU75_1-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU75_2-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU75_3-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU75_4-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU75_5-M_u2 Q d3 VSS VSS n w=0.525u l=0.18u
MU82-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MU81-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI79-MU3 net53 INCP XI79-net16 VSS n w=0.42u l=0.18u
MI79-MU4 XI79-net16 QD VSS VSS n w=0.42u l=0.18u
MI87-M_u2 d3 QD VDD VDD p w=3.3u l=0.18u
MI87-M_u1 d3 CP VDD VDD p w=3.3u l=0.18u
MI80-M_u3 QD net53 VDD VDD p w=0.685u l=0.18u
MU75_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU75_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU75_2-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU75_3-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU75_4-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU75_5-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU82-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MU81-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU16 net53 INCP net61 VDD p w=0.52u l=0.18u
MU17 net61 E net58 VDD p w=1.37u l=0.18u
MI81 net58 TE VDD VDD p w=1.37u l=0.18u
MI79-MU2 net53 INCPB XI79-net6 VDD p w=0.42u l=0.18u
MI79-MU1 XI79-net6 QD VDD VDD p w=0.42u l=0.18u
.ends
.subckt CKLNQD8BWP7T TE E CP Q VDD VSS 
MU19 net50 E VSS VSS n w=0.5u l=0.18u
MU20 net50 TE VSS VSS n w=0.5u l=0.18u
MI82 net53 INCPB net50 VSS n w=0.5u l=0.18u
MI87-M_u4 XI87-net6 QD VSS VSS n w=1.68u l=0.18u
MI87-M_u3 d3 CP XI87-net6 VSS n w=1.68u l=0.18u
MI80-M_u2 QD net53 VSS VSS n w=0.5u l=0.18u
MU75-M_u2 Q d3 VSS VSS n w=4.305u l=0.18u
MU82-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MU81-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI79-MU3 net53 INCP XI79-net16 VSS n w=0.42u l=0.18u
MI79-MU4 XI79-net16 QD VSS VSS n w=0.42u l=0.18u
MI87-M_u2 d3 QD VDD VDD p w=3.3u l=0.18u
MI87-M_u1 d3 CP VDD VDD p w=3.3u l=0.18u
MI80-M_u3 QD net53 VDD VDD p w=0.685u l=0.18u
MU75-M_u3 Q d3 VDD VDD p w=10.96u l=0.18u
MU82-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MU81-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU16 net53 INCP net61 VDD p w=0.52u l=0.18u
MU17 net61 E net58 VDD p w=1.37u l=0.18u
MI81 net58 TE VDD VDD p w=1.37u l=0.18u
MI79-MU2 net53 INCPB XI79-net6 VDD p w=0.42u l=0.18u
MI79-MU1 XI79-net6 QD VDD VDD p w=0.42u l=0.18u
.ends
.subckt CKMUX2D0BWP7T I0 I1 S Z VDD VSS 
MU29-M_u2 Z net28 VSS VSS n w=0.42u l=0.18u
MI111 net47 I0 VSS VSS n w=0.42u l=0.18u
MI5 net28 net6 net47 VSS n w=0.42u l=0.18u
MI14 net044 I1 VSS VSS n w=0.42u l=0.18u
MI13 net28 S net044 VSS n w=0.42u l=0.18u
MU24 net6 S VSS VSS n w=0.42u l=0.18u
MU29-M_u3 Z net28 VDD VDD p w=0.92u l=0.18u
MI2 VDD I0 net055 VDD p w=1.225u l=0.18u
MI4 net055 S net28 VDD p w=1.225u l=0.18u
MI12 net44 net6 net28 VDD p w=1.225u l=0.18u
MI10 VDD I1 net44 VDD p w=1.225u l=0.18u
MU25 VDD S net6 VDD p w=1.13u l=0.18u
.ends
.subckt CKMUX2D1BWP7T I0 I1 S Z VDD VSS 
MU29-M_u2 Z net28 VSS VSS n w=0.7u l=0.18u
MI111 net47 I0 VSS VSS n w=0.465u l=0.18u
MI5 net28 net6 net47 VSS n w=0.465u l=0.18u
MI7 net28 S net047 VSS n w=0.465u l=0.18u
MI8 net047 I1 VSS VSS n w=0.465u l=0.18u
MU24 net6 S VSS VSS n w=0.525u l=0.18u
MU29-M_u3 Z net28 VDD VDD p w=1.37u l=0.18u
MI2 VDD I0 net055 VDD p w=1.37u l=0.18u
MI4 net055 S net28 VDD p w=1.37u l=0.18u
MI9 net44 net6 net28 VDD p w=1.37u l=0.18u
MI10 VDD I1 net44 VDD p w=1.37u l=0.18u
MU25 VDD S net6 VDD p w=1.37u l=0.18u
.ends
.subckt CKMUX2D2BWP7T I0 I1 S Z VDD VSS 
MU29_0-M_u2 Z net28 VSS VSS n w=0.71u l=0.18u
MU29_1-M_u2 Z net28 VSS VSS n w=0.71u l=0.18u
MI111 net47 I0 VSS VSS n w=0.62u l=0.18u
MI5 net28 net6 net47 VSS n w=0.62u l=0.18u
MI7 net28 S net046 VSS n w=0.62u l=0.18u
MI8 net046 I1 VSS VSS n w=0.62u l=0.18u
MU24 net6 S VSS VSS n w=0.525u l=0.18u
MU29_0-M_u3 Z net28 VDD VDD p w=1.37u l=0.18u
MU29_1-M_u3 Z net28 VDD VDD p w=1.37u l=0.18u
MI2 VDD I0 net054 VDD p w=1.71u l=0.18u
MI4 net054 S net28 VDD p w=1.71u l=0.18u
MI9 net44 net6 net28 VDD p w=1.71u l=0.18u
MI10 VDD I1 net44 VDD p w=1.71u l=0.18u
MU25 VDD S net6 VDD p w=1.37u l=0.18u
.ends
.subckt CKND0BWP7T I ZN VDD VSS 
M_u2 ZN I VSS VSS n w=0.42u l=0.18u
M_u1 ZN I VDD VDD p w=1.13u l=0.18u
.ends
.subckt CKND10BWP7T I ZN VDD VSS 
DI3 VSS I dn 0.2037p
M_u2 ZN I VSS VSS n w=5.24u l=0.18u
M_u1 ZN I VDD VDD p w=13.695u l=0.18u
.ends
.subckt CKND12BWP7T I ZN VDD VSS 
DI3 VSS I dn 0.2037p
M_u2_0 ZN I VSS VSS n w=0.9u l=0.18u
M_u2_1 ZN I VSS VSS n w=0.9u l=0.18u
M_u2_2 ZN I VSS VSS n w=0.9u l=0.18u
M_u2_3 ZN I VSS VSS n w=0.9u l=0.18u
M_u2_4 ZN I VSS VSS n w=0.9u l=0.18u
M_u2_5 ZN I VSS VSS n w=0.9u l=0.18u
M_u2_6 ZN I VSS VSS n w=0.9u l=0.18u
M_u1_0 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_1 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_2 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_3 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_4 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_5 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_6 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_7 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_8 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_9 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_10 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_11 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKND1BWP7T I ZN VDD VSS 
M_u2 ZN I VSS VSS n w=0.525u l=0.18u
M_u1 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKND2BWP7T I ZN VDD VSS 
M_u2_0 ZN I VSS VSS n w=0.525u l=0.18u
M_u2_1 ZN I VSS VSS n w=0.525u l=0.18u
M_u1_0 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_1 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKND2D0BWP7T A1 A2 ZN VDD VSS 
MU1-M_u4 XU1-net6 A2 VSS VSS n w=0.42u l=0.18u
MU1-M_u3 ZN A1 XU1-net6 VSS n w=0.48u l=0.18u
MU1-M_u2 ZN A2 VDD VDD p w=0.8u l=0.18u
MU1-M_u1 ZN A1 VDD VDD p w=0.8u l=0.18u
.ends
.subckt CKND2D1BWP7T A1 A2 ZN VDD VSS 
MI0-M_u4 XI0-net6 A2 VSS VSS n w=0.685u l=0.18u
MI0-M_u3 ZN A1 XI0-net6 VSS n w=1u l=0.18u
MI0-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
MI0-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKND2D2BWP7T A1 A2 ZN VDD VSS 
MI0-M_u4 XI0-net6 A2 VSS VSS n w=1.2u l=0.18u
MI0-M_u3 ZN A1 XI0-net6 VSS n w=1.6u l=0.18u
MI0-M_u2 ZN A2 VDD VDD p w=2.74u l=0.18u
MI0-M_u1 ZN A1 VDD VDD p w=2.74u l=0.18u
.ends
.subckt CKND2D3BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 XI1-net6 A2 VSS VSS n w=1.8u l=0.18u
MI1-M_u3 ZN A1 XI1-net6 VSS n w=2.4u l=0.18u
MI1-M_u2 ZN A2 VDD VDD p w=4.11u l=0.18u
MI1-M_u1 ZN A1 VDD VDD p w=4.11u l=0.18u
.ends
.subckt CKND2D4BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 XI1-net6 A2 VSS VSS n w=2.4u l=0.18u
MI1-M_u3 ZN A1 XI1-net6 VSS n w=3.2u l=0.18u
MI1-M_u2 ZN A2 VDD VDD p w=5.48u l=0.18u
MI1-M_u1 ZN A1 VDD VDD p w=5.48u l=0.18u
.ends
.subckt CKND2D8BWP7T A1 A2 ZN VDD VSS 
MI21_0 ZN A1 N1 VSS n w=1u l=0.18u
MI21_1 ZN A1 N1 VSS n w=1u l=0.18u
MI21_2 ZN A1 N1 VSS n w=1u l=0.18u
MI21_3 ZN A1 N1 VSS n w=1u l=0.18u
MI21_4 ZN A1 N1 VSS n w=1u l=0.18u
MI21_5 ZN A1 N1 VSS n w=1u l=0.18u
MI21_6 ZN A1 N1 VSS n w=1u l=0.18u
MI21_7 ZN A1 N1 VSS n w=1u l=0.18u
MI20_0 N1 A2 VSS VSS n w=0.68u l=0.18u
MI20_1 N1 A2 VSS VSS n w=0.68u l=0.18u
MI20_2 N1 A2 VSS VSS n w=0.68u l=0.18u
MI20_3 N1 A2 VSS VSS n w=0.68u l=0.18u
MI20_4 N1 A2 VSS VSS n w=0.68u l=0.18u
MI20_5 N1 A2 VSS VSS n w=0.68u l=0.18u
MI20_6 N1 A2 VSS VSS n w=0.68u l=0.18u
MI20_7 N1 A2 VSS VSS n w=0.68u l=0.18u
M_u2_0 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_1 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_2 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_3 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_4 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_5 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_6 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_7 ZN A2 VDD VDD p w=1.37u l=0.18u
MI6_0 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_2 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_3 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_4 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_5 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_6 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_7 ZN A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKND3BWP7T I ZN VDD VSS 
DI3 VSS I dn 0.2037p
M_u2_0 ZN I VSS VSS n w=0.525u l=0.18u
M_u2_1 ZN I VSS VSS n w=0.525u l=0.18u
M_u2_2 ZN I VSS VSS n w=0.525u l=0.18u
M_u1_0 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_1 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_2 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKND4BWP7T I ZN VDD VSS 
DI3 VSS I dn 0.2037p
M_u2_0 ZN I VSS VSS n w=0.7u l=0.18u
M_u2_1 ZN I VSS VSS n w=0.7u l=0.18u
M_u2_2 ZN I VSS VSS n w=0.7u l=0.18u
M_u1_0 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_1 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_2 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_3 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKND6BWP7T I ZN VDD VSS 
DI3 VSS I dn 0.2037p
M_u2_0 ZN I VSS VSS n w=0.79u l=0.18u
M_u2_1 ZN I VSS VSS n w=0.79u l=0.18u
M_u2_2 ZN I VSS VSS n w=0.79u l=0.18u
M_u2_3 ZN I VSS VSS n w=0.79u l=0.18u
M_u1_0 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_1 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_2 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_3 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_4 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_5 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKND8BWP7T I ZN VDD VSS 
DI3 VSS I dn 0.2037p
M_u2_0 ZN I VSS VSS n w=0.84u l=0.18u
M_u2_1 ZN I VSS VSS n w=0.84u l=0.18u
M_u2_2 ZN I VSS VSS n w=0.84u l=0.18u
M_u2_3 ZN I VSS VSS n w=0.84u l=0.18u
M_u2_4 ZN I VSS VSS n w=0.84u l=0.18u
M_u1_0 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_1 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_2 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_3 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_4 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_5 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_6 ZN I VDD VDD p w=1.37u l=0.18u
M_u1_7 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt CKXOR2D0BWP7T A1 A2 Z VDD VSS 
MI5 net14 A1 net016 VSS n w=0.42u l=0.18u
MI111 net016 net4 VSS VSS n w=0.42u l=0.18u
M_u6-M_u2 net4 net10 net14 VSS n w=0.42u l=0.18u
MI1-M_u2 net4 A2 VSS VSS n w=0.42u l=0.18u
M_u4-M_u2 Z net14 VSS VSS n w=0.42u l=0.18u
MI2-M_u2 net10 A1 VSS VSS n w=0.94u l=0.18u
MI6 VDD net4 net024 VDD p w=0.94u l=0.18u
MI4 net024 net10 net14 VDD p w=0.94u l=0.18u
M_u6-M_u3 net4 A1 net14 VDD p w=1.185u l=0.18u
MI1-M_u3 net4 A2 VDD VDD p w=0.94u l=0.18u
M_u4-M_u3 Z net14 VDD VDD p w=0.88u l=0.18u
MI2-M_u3 net10 A1 VDD VDD p w=0.6u l=0.18u
.ends
.subckt CKXOR2D1BWP7T A1 A2 Z VDD VSS 
MI5 net14 A1 net016 VSS n w=0.42u l=0.18u
MI111 net016 net4 VSS VSS n w=0.42u l=0.18u
M_u6-M_u2 net4 net10 net14 VSS n w=0.42u l=0.18u
MI1-M_u2 net4 A2 VSS VSS n w=0.42u l=0.18u
M_u4-M_u2 Z net14 VSS VSS n w=0.8u l=0.18u
MI2-M_u2 net10 A1 VSS VSS n w=0.94u l=0.18u
MI6 VDD net4 net024 VDD p w=0.94u l=0.18u
MI4 net024 net10 net14 VDD p w=0.94u l=0.18u
M_u6-M_u3 net4 A1 net14 VDD p w=1.185u l=0.18u
MI1-M_u3 net4 A2 VDD VDD p w=1u l=0.18u
M_u4-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
MI2-M_u3 net10 A1 VDD VDD p w=0.6u l=0.18u
.ends
.subckt CKXOR2D2BWP7T A1 A2 Z VDD VSS 
MI5 net14 A1 net016 VSS n w=0.6u l=0.18u
MI111 net016 net4 VSS VSS n w=0.42u l=0.18u
M_u6-M_u2 net4 net10 net14 VSS n w=0.8u l=0.18u
MI1-M_u2 net4 A2 VSS VSS n w=0.6u l=0.18u
M_u4_0-M_u2 Z net14 VSS VSS n w=1u l=0.18u
M_u4_1-M_u2 Z net14 VSS VSS n w=1u l=0.18u
MI2-M_u2 net10 A1 VSS VSS n w=0.94u l=0.18u
MI6 VDD net4 net024 VDD p w=1.2u l=0.18u
MI4 net024 net10 net14 VDD p w=1.2u l=0.18u
M_u6-M_u3 net4 A1 net14 VDD p w=1.185u l=0.18u
MI1-M_u3 net4 A2 VDD VDD p w=1.2u l=0.18u
M_u4_0-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
M_u4_1-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
MI2-M_u3 net10 A1 VDD VDD p w=0.6u l=0.18u
.ends
.subckt CKXOR2D4BWP7T A1 A2 Z VDD VSS 
MI5 net14 A1 net016 VSS n w=0.84u l=0.18u
MI111 net016 net4 VSS VSS n w=1u l=0.18u
M_u6_0-M_u2 net4 net10 net14 VSS n w=0.42u l=0.18u
M_u6_1-M_u2 net4 net10 net14 VSS n w=0.42u l=0.18u
MI1-M_u2 net4 A2 VSS VSS n w=1.5u l=0.18u
M_u4_0-M_u2 Z net14 VSS VSS n w=1.2u l=0.18u
M_u4_1-M_u2 Z net14 VSS VSS n w=1.2u l=0.18u
MI2-M_u2 net10 A1 VSS VSS n w=0.525u l=0.18u
MI6 VDD net4 net016 VDD p w=3.015u l=0.18u
MI4 net016 net10 net14 VDD p w=2.07u l=0.18u
M_u6_0-M_u3 net4 A1 net14 VDD p w=1.13u l=0.18u
M_u6_1-M_u3 net4 A1 net14 VDD p w=1.13u l=0.18u
MI1-M_u3 net4 A2 VDD VDD p w=4.11u l=0.18u
M_u4_0-M_u3 Z net14 VDD VDD p w=2.74u l=0.18u
M_u4_1-M_u3 Z net14 VDD VDD p w=2.74u l=0.18u
MI2-M_u3 net10 A1 VDD VDD p w=1.31u l=0.18u
.ends
.subckt DCAP16BWP7T VDD VSS 
MI7 VSS net6 VSS VSS n w=4.7u l=0.965u
M_u2 net8 net6 VSS VSS n w=0.94u l=0.18u
MI5 VDD net8 VDD VDD p w=6.335u l=0.965u
M_u1 net6 net8 VDD VDD p w=1.095u l=0.18u
.ends
.subckt DCAP32BWP7T VDD VSS 
M_u2 net20 net12 VSS VSS n w=1.88u l=0.18u
MI7 VSS net12 VSS VSS n w=9.4u l=1.035u
MI5 VDD net20 VDD VDD p w=12.67u l=1.035u
M_u1 net12 net20 VDD VDD p w=2.19u l=0.18u
.ends
.subckt DCAP4BWP7T VDD VSS 
MI4 VSS net6 VSS VSS n w=1u l=0.28u
M_u2 net8 net6 VSS VSS n w=1u l=0.18u
MI3 VDD net8 VDD VDD p w=1.17u l=0.28u
M_u1 net6 net8 VDD VDD p w=1.17u l=0.18u
.ends
.subckt DCAP64BWP7T VDD VSS 
M_u2 net81 net55 VSS VSS n w=1.88u l=0.18u
MI7 VSS net55 VSS VSS n w=20.68u l=0.99u
M_u1 net55 net81 VDD VDD p w=2.19u l=0.18u
MI5 VDD net81 VDD VDD p w=28.39u l=0.99u
.ends
.subckt DCAP8BWP7T VDD VSS 
MI4 VSS net6 VSS VSS n w=1.89u l=0.99u
M_u2 net8 net6 VSS VSS n w=0.945u l=0.18u
MI3 VDD net8 VDD VDD p w=2.605u l=0.99u
M_u1 net6 net8 VDD VDD p w=1.235u l=0.18u
.ends
.subckt DCAPBWP7T VDD VSS 
M_u2 net8 net6 VSS VSS n w=1u l=0.18u
M_u1 net6 net8 VDD VDD p w=1.37u l=0.18u
.ends
.subckt DEL015BWP7T I Z VDD VSS 
MI15-M_u2 net3 I VSS VSS n w=1u l=0.18u
MI2-M_u2 Z net3 VSS VSS n w=0.52u l=0.18u
MI15-M_u3 net3 I VDD VDD p w=1.37u l=0.18u
MI2-M_u3 Z net3 VDD VDD p w=1.06u l=0.18u
.ends
.subckt DEL01BWP7T I Z VDD VSS 
MI15-M_u2 net3 I VSS VSS n w=1u l=0.18u
MI2-M_u2 Z net3 VSS VSS n w=1u l=0.18u
MI15-M_u3 net3 I VDD VDD p w=1.37u l=0.18u
MI2-M_u3 Z net3 VDD VDD p w=1.37u l=0.18u
.ends
.subckt DEL02BWP7T I Z VDD VSS 
MI15-M_u2 net3 I VSS VSS n w=0.76u l=0.18u
MI2-M_u2 Z net3 VSS VSS n w=0.42u l=0.18u
MI15-M_u3 net3 I VDD VDD p w=0.42u l=0.18u
MI2-M_u3 Z net3 VDD VDD p w=0.66u l=0.18u
.ends
.subckt DEL0BWP7T I Z VDD VSS 
MI2-M_u2 Z net3 VSS VSS n w=1u l=0.18u
MU7-M_u2 net3 net5 VSS VSS n w=0.7u l=0.28u
MU5-M_u2 net5 net9 VSS VSS n w=0.67u l=0.28u
MI1-M_u2 net9 I VSS VSS n w=0.5u l=0.18u
MI2-M_u3 Z net3 VDD VDD p w=1.37u l=0.18u
MU7-M_u3 net3 net5 VDD VDD p w=0.9u l=0.28u
MU5-M_u3 net5 net9 VDD VDD p w=0.79u l=0.28u
MI1-M_u3 net9 I VDD VDD p w=0.685u l=0.18u
.ends
.subckt DEL1BWP7T I Z VDD VSS 
MI2-M_u2 Z net3 VSS VSS n w=1u l=0.18u
MU7-M_u2 net3 net5 VSS VSS n w=0.6u l=0.7u
MU5-M_u2 net5 net9 VSS VSS n w=0.83u l=0.7u
MI1-M_u2 net9 I VSS VSS n w=0.5u l=0.18u
MI2-M_u3 Z net3 VDD VDD p w=1.37u l=0.18u
MU7-M_u3 net3 net5 VDD VDD p w=0.9u l=0.7u
MU5-M_u3 net5 net9 VDD VDD p w=1.2u l=0.7u
MI1-M_u3 net9 I VDD VDD p w=0.685u l=0.18u
.ends
.subckt DEL2BWP7T I Z VDD VSS 
MI2-M_u2 Z net3 VSS VSS n w=1u l=0.18u
MU7-M_u2 net3 net5 VSS VSS n w=0.45u l=1.25u
MU5-M_u2 net5 net9 VSS VSS n w=0.6u l=1.25u
MI1-M_u2 net9 I VSS VSS n w=0.5u l=0.18u
MI2-M_u3 Z net3 VDD VDD p w=1.37u l=0.18u
MU7-M_u3 net3 net5 VDD VDD p w=0.58u l=1.25u
MU5-M_u3 net5 net9 VDD VDD p w=0.95u l=1.25u
MI1-M_u3 net9 I VDD VDD p w=0.685u l=0.18u
.ends
.subckt DEL3BWP7T I Z VDD VSS 
MI8-M_u2 net010 net08 VSS VSS n w=0.55u l=0.95u
MI9-M_u2 net08 net9 VSS VSS n w=0.58u l=0.95u
MI6-M_u2 net9 net012 VSS VSS n w=0.58u l=0.95u
MI2-M_u2 Z net010 VSS VSS n w=1u l=0.18u
MI5-M_u2 net012 net014 VSS VSS n w=0.5u l=0.95u
MI1-M_u2 net014 I VSS VSS n w=0.5u l=0.18u
MI8-M_u3 net010 net08 VDD VDD p w=0.48u l=0.95u
MI9-M_u3 net08 net9 VDD VDD p w=0.96u l=0.95u
MI6-M_u3 net9 net012 VDD VDD p w=0.96u l=0.95u
MI2-M_u3 Z net010 VDD VDD p w=1.37u l=0.18u
MI5-M_u3 net012 net014 VDD VDD p w=0.67u l=0.95u
MI1-M_u3 net014 I VDD VDD p w=0.685u l=0.18u
.ends
.subckt DEL4BWP7T I Z VDD VSS 
MI4-M_u2 net08 net9 VSS VSS n w=0.7u l=1.2u
MI6-M_u2 net9 net012 VSS VSS n w=0.7u l=1.2u
MI3-M_u2 net010 net08 VSS VSS n w=0.49u l=1.2u
MI2-M_u2 Z net010 VSS VSS n w=1u l=0.18u
MI5-M_u2 net012 net014 VSS VSS n w=0.55u l=1.2u
MI1-M_u2 net014 I VSS VSS n w=0.5u l=0.18u
MI4-M_u3 net08 net9 VDD VDD p w=0.93u l=1.2u
MI6-M_u3 net9 net012 VDD VDD p w=0.93u l=1.2u
MI3-M_u3 net010 net08 VDD VDD p w=0.5u l=1.2u
MI2-M_u3 Z net010 VDD VDD p w=1.37u l=0.18u
MI5-M_u3 net012 net014 VDD VDD p w=0.8u l=1.2u
MI1-M_u3 net014 I VDD VDD p w=0.685u l=0.18u
.ends
.subckt DFCND0BWP7T D CP CDN Q QN VDD VSS 
MI4 net52 INCPB VSS VSS n w=0.94u l=0.18u
MI15 d1 INCP d2 VSS n w=0.91u l=0.18u
MI5 d0 D net52 VSS n w=0.94u l=0.18u
MI18 net101 INCPB d2 VSS n w=0.42u l=0.18u
MI47 d0 INCP net59 VSS n w=0.42u l=0.18u
MI48 net59 CDN net62 VSS n w=0.42u l=0.18u
MI49 net62 d1 VSS VSS n w=0.42u l=0.18u
MI21-M_u4 XI21-net6 CDN VSS VSS n w=0.97u l=0.18u
MI21-M_u3 d3 d2 XI21-net6 VSS n w=0.97u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net101 VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net101 d3 VSS VSS n w=0.42u l=0.18u
MI21-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI21-M_u1 d3 d2 VDD VDD p w=1.31u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net101 VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI14-M_u3 net101 d3 VDD VDD p w=0.6u l=0.18u
MI6 d0 D net85 VDD p w=1.37u l=0.18u
MI7 net85 INCP VDD VDD p w=1.37u l=0.18u
MI16 d1 INCPB d2 VDD p w=0.62u l=0.18u
MI17 net101 INCP d2 VDD p w=0.42u l=0.18u
MI45 d0 INCPB net98 VDD p w=0.42u l=0.18u
MI43 net98 d1 VDD VDD p w=0.42u l=0.18u
MI44 net98 CDN VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFCND1BWP7T D CP CDN Q QN VDD VSS 
MI4 net52 INCPB VSS VSS n w=0.94u l=0.18u
MI15 d1 INCP d2 VSS n w=0.91u l=0.18u
MI5 d0 D net52 VSS n w=0.94u l=0.18u
MI18 net101 INCPB d2 VSS n w=0.42u l=0.18u
MI47 d0 INCP net59 VSS n w=0.42u l=0.18u
MI48 net59 CDN net62 VSS n w=0.42u l=0.18u
MI49 net62 d1 VSS VSS n w=0.42u l=0.18u
MI21-M_u4 XI21-net6 CDN VSS VSS n w=0.97u l=0.18u
MI21-M_u3 d3 d2 XI21-net6 VSS n w=0.97u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net101 VSS VSS n w=0.94u l=0.18u
MI27-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net101 d3 VSS VSS n w=0.42u l=0.18u
MI21-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI21-M_u1 d3 d2 VDD VDD p w=1.37u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net101 VDD VDD p w=0.835u l=0.18u
MI27-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI14-M_u3 net101 d3 VDD VDD p w=0.6u l=0.18u
MI6 d0 D net85 VDD p w=1.37u l=0.18u
MI7 net85 INCP VDD VDD p w=1.37u l=0.18u
MI16 d1 INCPB d2 VDD p w=0.62u l=0.18u
MI17 net101 INCP d2 VDD p w=0.42u l=0.18u
MI45 d0 INCPB net98 VDD p w=0.42u l=0.18u
MI43 net98 d1 VDD VDD p w=0.42u l=0.18u
MI44 net98 CDN VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFCND2BWP7T D CP CDN Q QN VDD VSS 
MI4 net52 INCPB VSS VSS n w=0.94u l=0.18u
MI15 d1 INCP d2 VSS n w=0.91u l=0.18u
MI5 d0 D net52 VSS n w=0.94u l=0.18u
MI18 net059 INCPB d2 VSS n w=0.42u l=0.18u
MI47 d0 INCP net59 VSS n w=0.42u l=0.18u
MI48 net59 CDN net62 VSS n w=0.42u l=0.18u
MI49 net62 d1 VSS VSS n w=0.42u l=0.18u
MI21-M_u4 XI21-net6 CDN VSS VSS n w=0.97u l=0.18u
MI21-M_u3 d3 d2 XI21-net6 VSS n w=0.97u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29_0-M_u2 QN net059 VSS VSS n w=1u l=0.18u
MI29_1-M_u2 QN net059 VSS VSS n w=1u l=0.18u
MI27_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net059 d3 VSS VSS n w=0.97u l=0.18u
MI21-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI21-M_u1 d3 d2 VDD VDD p w=1.23u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29_0-M_u3 QN net059 VDD VDD p w=1.3u l=0.18u
MI29_1-M_u3 QN net059 VDD VDD p w=1.3u l=0.18u
MI27_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI14-M_u3 net059 d3 VDD VDD p w=0.97u l=0.18u
MI6 d0 D net85 VDD p w=1.37u l=0.18u
MI7 net85 INCP VDD VDD p w=1.37u l=0.18u
MI16 d1 INCPB d2 VDD p w=0.62u l=0.18u
MI17 net059 INCP d2 VDD p w=0.42u l=0.18u
MI45 d0 INCPB net98 VDD p w=0.42u l=0.18u
MI43 net98 d1 VDD VDD p w=0.42u l=0.18u
MI44 net98 CDN VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFCNQD1BWP7T D CP CDN Q VDD VSS 
MI4 net52 INCPB VSS VSS n w=0.94u l=0.18u
MI15 d1 INCP d2 VSS n w=0.91u l=0.18u
MI5 d0 D net52 VSS n w=0.94u l=0.18u
MI18 net101 INCPB d2 VSS n w=0.42u l=0.18u
MI47 d0 INCP net59 VSS n w=0.42u l=0.18u
MI48 net59 CDN net62 VSS n w=0.42u l=0.18u
MI49 net62 d1 VSS VSS n w=0.42u l=0.18u
MI21-M_u4 XI21-net6 CDN VSS VSS n w=0.97u l=0.18u
MI21-M_u3 d3 d2 XI21-net6 VSS n w=0.97u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net101 d3 VSS VSS n w=0.42u l=0.18u
MI21-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI21-M_u1 d3 d2 VDD VDD p w=1.37u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI14-M_u3 net101 d3 VDD VDD p w=0.42u l=0.18u
MI6 d0 D net85 VDD p w=1.37u l=0.18u
MI7 net85 INCP VDD VDD p w=1.37u l=0.18u
MI16 d1 INCPB d2 VDD p w=0.62u l=0.18u
MI17 net101 INCP d2 VDD p w=0.42u l=0.18u
MI45 d0 INCPB net98 VDD p w=0.42u l=0.18u
MI43 net98 d1 VDD VDD p w=0.42u l=0.18u
MI44 net98 CDN VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFCNQD2BWP7T D CP CDN Q VDD VSS 
MI4 net52 INCPB VSS VSS n w=0.94u l=0.18u
MI15 d1 INCP d2 VSS n w=0.91u l=0.18u
MI5 d0 D net52 VSS n w=0.94u l=0.18u
MI18 net101 INCPB d2 VSS n w=0.42u l=0.18u
MI47 d0 INCP net59 VSS n w=0.42u l=0.18u
MI48 net59 CDN net62 VSS n w=0.42u l=0.18u
MI49 net62 d1 VSS VSS n w=0.42u l=0.18u
MI21-M_u4 XI21-net6 CDN VSS VSS n w=0.97u l=0.18u
MI21-M_u3 d3 d2 XI21-net6 VSS n w=0.97u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net101 d3 VSS VSS n w=0.42u l=0.18u
MI21-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI21-M_u1 d3 d2 VDD VDD p w=1.37u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI14-M_u3 net101 d3 VDD VDD p w=0.42u l=0.18u
MI6 d0 D net85 VDD p w=1.37u l=0.18u
MI7 net85 INCP VDD VDD p w=1.37u l=0.18u
MI16 d1 INCPB d2 VDD p w=0.62u l=0.18u
MI17 net101 INCP d2 VDD p w=0.42u l=0.18u
MI45 d0 INCPB net98 VDD p w=0.42u l=0.18u
MI43 net98 d1 VDD VDD p w=0.42u l=0.18u
MI44 net98 CDN VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFD0BWP7T D CP Q QN VDD VSS 
MI4 net43 INCPB VSS VSS n w=0.94u l=0.18u
MI5 P000 D net43 VSS n w=0.94u l=0.18u
MI47 P000 INCP net50 VSS n w=0.42u l=0.18u
MI48 net50 P0001 VSS VSS n w=0.42u l=0.18u
MI55 P0002 INCPB N0028 VSS n w=0.42u l=0.18u
MI50 P0001 INCP N0028 VSS n w=0.91u l=0.18u
MI56-M_u2 P0002 P0003 VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN P0002 VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q P0003 VSS VSS n w=0.5u l=0.18u
MI53-M_u2 P0003 N0028 VSS VSS n w=0.5u l=0.18u
MI13-M_u2 P0001 P000 VSS VSS n w=0.54u l=0.18u
MI56-M_u3 P0002 P0003 VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN P0002 VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q P0003 VDD VDD p w=0.685u l=0.18u
MI53-M_u3 P0003 N0028 VDD VDD p w=0.685u l=0.18u
MI13-M_u3 P0001 P000 VDD VDD p w=0.96u l=0.18u
MI6 P000 D net74 VDD p w=0.92u l=0.18u
MI7 net74 INCP VDD VDD p w=0.92u l=0.18u
MI52 P0001 INCPB N0028 VDD p w=1.34u l=0.18u
MI54 P0002 INCP N0028 VDD p w=0.42u l=0.18u
MI45 P000 INCPB net86 VDD p w=0.42u l=0.18u
MI43 net86 P0001 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFD1BWP7T D CP Q QN VDD VSS 
MI4 net43 INCPB VSS VSS n w=0.94u l=0.18u
MI5 P000 D net43 VSS n w=0.94u l=0.18u
MI47 P000 INCP net50 VSS n w=0.42u l=0.18u
MI48 net50 P0001 VSS VSS n w=0.42u l=0.18u
MI55 P0002 INCPB N0028 VSS n w=0.42u l=0.18u
MI50 P0001 INCP N0028 VSS n w=0.91u l=0.18u
MI56-M_u2 P0002 P0003 VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN P0002 VSS VSS n w=0.94u l=0.18u
MI27-M_u2 Q P0003 VSS VSS n w=1u l=0.18u
MI53-M_u2 P0003 N0028 VSS VSS n w=1u l=0.18u
MI13-M_u2 P0001 P000 VSS VSS n w=0.54u l=0.18u
MI56-M_u3 P0002 P0003 VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN P0002 VDD VDD p w=1.37u l=0.18u
MI27-M_u3 Q P0003 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 P0003 N0028 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 P0001 P000 VDD VDD p w=0.96u l=0.18u
MI6 P000 D net74 VDD p w=0.92u l=0.18u
MI7 net74 INCP VDD VDD p w=0.92u l=0.18u
MI52 P0001 INCPB N0028 VDD p w=1.34u l=0.18u
MI54 P0002 INCP N0028 VDD p w=0.42u l=0.18u
MI45 P000 INCPB net86 VDD p w=0.42u l=0.18u
MI43 net86 P0001 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFD2BWP7T D CP Q QN VDD VSS 
MI4 net43 INCPB VSS VSS n w=0.94u l=0.18u
MI5 P000 D net43 VSS n w=0.94u l=0.18u
MI47 P000 INCP net50 VSS n w=0.42u l=0.18u
MI48 net50 P0001 VSS VSS n w=0.42u l=0.18u
MI55 P0002 INCPB N0028 VSS n w=0.42u l=0.18u
MI50 P0001 INCP N0028 VSS n w=0.91u l=0.18u
MI56-M_u2 P0002 P0003 VSS VSS n w=1u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN P0002 VSS VSS n w=2u l=0.18u
MI27_0-M_u2 Q P0003 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q P0003 VSS VSS n w=1u l=0.18u
MI53_0-M_u2 P0003 N0028 VSS VSS n w=1u l=0.18u
MI53_1-M_u2 P0003 N0028 VSS VSS n w=1u l=0.18u
MI13-M_u2 P0001 P000 VSS VSS n w=0.54u l=0.18u
MI56-M_u3 P0002 P0003 VDD VDD p w=1.37u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN P0002 VDD VDD p w=2.605u l=0.18u
MI27_0-M_u3 Q P0003 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q P0003 VDD VDD p w=1.37u l=0.18u
MI53_0-M_u3 P0003 N0028 VDD VDD p w=1.235u l=0.18u
MI53_1-M_u3 P0003 N0028 VDD VDD p w=1.235u l=0.18u
MI13-M_u3 P0001 P000 VDD VDD p w=0.96u l=0.18u
MI6 P000 D net74 VDD p w=0.92u l=0.18u
MI7 net74 INCP VDD VDD p w=0.92u l=0.18u
MI52 P0001 INCPB N0028 VDD p w=1.34u l=0.18u
MI54 P0002 INCP N0028 VDD p w=0.42u l=0.18u
MI45 P000 INCPB net86 VDD p w=0.42u l=0.18u
MI43 net86 P0001 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFKCND0BWP7T D CP CN Q QN VDD VSS 
MI15 net38 CN VSS VSS n w=0.97u l=0.18u
MI12 net64 INCPB net39 VSS n w=0.97u l=0.18u
MI47 net64 INCP net54 VSS n w=0.42u l=0.18u
MI48 net54 net55 VSS VSS n w=0.42u l=0.18u
MI55 net51 INCPB net47 VSS n w=0.42u l=0.18u
MI50 net55 INCP net47 VSS n w=0.91u l=0.18u
MI16 net39 D net38 VSS n w=0.97u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net51 VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q net88 VSS VSS n w=0.5u l=0.18u
MI53-M_u2 net88 net47 VSS VSS n w=0.5u l=0.18u
MI13-M_u2 net55 net64 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net51 net88 VSS VSS n w=0.42u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net51 VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q net88 VDD VDD p w=0.685u l=0.18u
MI53-M_u3 net88 net47 VDD VDD p w=0.685u l=0.18u
MI13-M_u3 net55 net64 VDD VDD p w=0.96u l=0.18u
MI14-M_u3 net51 net88 VDD VDD p w=0.685u l=0.18u
MI17 VDD D net62 VDD p w=0.95u l=0.18u
MI52 net55 INCPB net47 VDD p w=1.34u l=0.18u
MI54 net51 INCP net47 VDD p w=0.42u l=0.18u
MI45 net64 INCPB net73 VDD p w=0.42u l=0.18u
MI43 net73 net55 VDD VDD p w=0.42u l=0.18u
MI18 net62 INCP net64 VDD p w=0.65u l=0.18u
MI19 VDD CN net62 VDD p w=0.42u l=0.18u
.ends
.subckt DFKCND1BWP7T D CP CN Q QN VDD VSS 
MI15 net38 CN VSS VSS n w=0.97u l=0.18u
MI12 net64 INCPB net39 VSS n w=0.97u l=0.18u
MI47 net64 INCP net54 VSS n w=0.42u l=0.18u
MI48 net54 net55 VSS VSS n w=0.42u l=0.18u
MI55 net51 INCPB net47 VSS n w=0.42u l=0.18u
MI50 net55 INCP net47 VSS n w=0.91u l=0.18u
MI16 net39 D net38 VSS n w=0.97u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net51 VSS VSS n w=0.94u l=0.18u
MI27-M_u2 Q net88 VSS VSS n w=1u l=0.18u
MI53-M_u2 net88 net47 VSS VSS n w=1u l=0.18u
MI13-M_u2 net55 net64 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net51 net88 VSS VSS n w=0.42u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net51 VDD VDD p w=1.37u l=0.18u
MI27-M_u3 Q net88 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 net88 net47 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 net55 net64 VDD VDD p w=0.96u l=0.18u
MI14-M_u3 net51 net88 VDD VDD p w=0.685u l=0.18u
MI17 VDD D net62 VDD p w=0.95u l=0.18u
MI52 net55 INCPB net47 VDD p w=1.34u l=0.18u
MI54 net51 INCP net47 VDD p w=0.42u l=0.18u
MI45 net64 INCPB net73 VDD p w=0.42u l=0.18u
MI43 net73 net55 VDD VDD p w=0.42u l=0.18u
MI18 net62 INCP net64 VDD p w=0.65u l=0.18u
MI19 VDD CN net62 VDD p w=0.42u l=0.18u
.ends
.subckt DFKCND2BWP7T D CP CN Q QN VDD VSS 
MI15 net38 CN VSS VSS n w=0.97u l=0.18u
MI12 net64 INCPB net39 VSS n w=0.97u l=0.18u
MI47 net64 INCP net54 VSS n w=0.42u l=0.18u
MI48 net54 net55 VSS VSS n w=0.42u l=0.18u
MI55 net060 INCPB net47 VSS n w=0.42u l=0.18u
MI50 net55 INCP net47 VSS n w=0.91u l=0.18u
MI16 net39 D net38 VSS n w=0.97u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29_0-M_u2 QN net060 VSS VSS n w=1u l=0.18u
MI29_1-M_u2 QN net060 VSS VSS n w=1u l=0.18u
MI27_0-M_u2 Q net076 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q net076 VSS VSS n w=1u l=0.18u
MI53-M_u2 net076 net47 VSS VSS n w=1u l=0.18u
MI13-M_u2 net55 net64 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net060 net076 VSS VSS n w=1u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29_0-M_u3 QN net060 VDD VDD p w=1.3u l=0.18u
MI29_1-M_u3 QN net060 VDD VDD p w=1.3u l=0.18u
MI27_0-M_u3 Q net076 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q net076 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 net076 net47 VDD VDD p w=1.23u l=0.18u
MI13-M_u3 net55 net64 VDD VDD p w=0.96u l=0.18u
MI14-M_u3 net060 net076 VDD VDD p w=1.37u l=0.18u
MI17 VDD D net62 VDD p w=0.95u l=0.18u
MI52 net55 INCPB net47 VDD p w=1.34u l=0.18u
MI54 net060 INCP net47 VDD p w=0.42u l=0.18u
MI45 net64 INCPB net73 VDD p w=0.42u l=0.18u
MI43 net73 net55 VDD VDD p w=0.42u l=0.18u
MI18 net62 INCP net64 VDD p w=0.65u l=0.18u
MI19 VDD CN net62 VDD p w=0.42u l=0.18u
.ends
.subckt DFKCNQD1BWP7T D CP CN Q VDD VSS 
MI15 net38 CN VSS VSS n w=0.97u l=0.18u
MI12 net64 INCPB net39 VSS n w=0.97u l=0.18u
MI47 net64 INCP net54 VSS n w=0.42u l=0.18u
MI48 net54 net55 VSS VSS n w=0.42u l=0.18u
MI50 net55 INCP net049 VSS n w=0.91u l=0.18u
MI16 net39 D net38 VSS n w=0.97u l=0.18u
MI22 net049 INCPB net048 VSS n w=0.42u l=0.18u
MI23 net048 net51 VSS VSS n w=0.42u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q net51 VSS VSS n w=1u l=0.18u
MI53-M_u2 net51 net049 VSS VSS n w=1u l=0.18u
MI13-M_u2 net55 net64 VSS VSS n w=0.54u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q net51 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 net51 net049 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 net55 net64 VDD VDD p w=0.96u l=0.18u
MI17 VDD D net62 VDD p w=0.95u l=0.18u
MI52 net55 INCPB net049 VDD p w=1.34u l=0.18u
MI45 net64 INCPB net73 VDD p w=0.42u l=0.18u
MI43 net73 net55 VDD VDD p w=0.42u l=0.18u
MI18 net62 INCP net64 VDD p w=0.65u l=0.18u
MI25 net049 INCP net084 VDD p w=0.42u l=0.18u
MI26 net084 net51 VDD VDD p w=0.42u l=0.18u
MI19 VDD CN net62 VDD p w=0.42u l=0.18u
.ends
.subckt DFKCNQD2BWP7T D CP CN Q VDD VSS 
MI15 net38 CN VSS VSS n w=0.97u l=0.18u
MI12 net64 INCPB net39 VSS n w=0.97u l=0.18u
MI47 net64 INCP net54 VSS n w=0.42u l=0.18u
MI48 net54 net55 VSS VSS n w=0.42u l=0.18u
MI50 net55 INCP net049 VSS n w=0.91u l=0.18u
MI16 net39 D net38 VSS n w=0.97u l=0.18u
MI22 net049 INCPB net048 VSS n w=0.42u l=0.18u
MI23 net048 net076 VSS VSS n w=0.42u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27_0-M_u2 Q net076 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q net076 VSS VSS n w=1u l=0.18u
MI53-M_u2 net076 net049 VSS VSS n w=1u l=0.18u
MI13-M_u2 net55 net64 VSS VSS n w=0.54u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27_0-M_u3 Q net076 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q net076 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 net076 net049 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 net55 net64 VDD VDD p w=0.96u l=0.18u
MI17 VDD D net62 VDD p w=0.95u l=0.18u
MI52 net55 INCPB net049 VDD p w=1.34u l=0.18u
MI45 net64 INCPB net73 VDD p w=0.42u l=0.18u
MI43 net73 net55 VDD VDD p w=0.42u l=0.18u
MI18 net62 INCP net64 VDD p w=0.65u l=0.18u
MI25 net049 INCP net084 VDD p w=0.42u l=0.18u
MI26 net084 net076 VDD VDD p w=0.42u l=0.18u
MI19 VDD CN net62 VDD p w=0.42u l=0.18u
.ends
.subckt DFKSND0BWP7T D CP SN Q QN VDD VSS 
MI15 net44 D VSS VSS n w=1u l=0.18u
MI12 net64 INCPB net44 VSS n w=0.94u l=0.18u
MI47 net64 INCP net56 VSS n w=0.42u l=0.18u
MI48 net56 net55 VSS VSS n w=0.42u l=0.18u
MI55 net51 INCPB net47 VSS n w=0.42u l=0.18u
MI50 net55 INCP net47 VSS n w=0.91u l=0.18u
MI16 net44 net84 VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net51 VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q net90 VSS VSS n w=0.5u l=0.18u
MI53-M_u2 net90 net47 VSS VSS n w=0.5u l=0.18u
MI13-M_u2 net55 net64 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net51 net90 VSS VSS n w=0.5u l=0.18u
MI20-M_u2 net84 SN VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net51 VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q net90 VDD VDD p w=0.685u l=0.18u
MI53-M_u3 net90 net47 VDD VDD p w=0.685u l=0.18u
MI13-M_u3 net55 net64 VDD VDD p w=0.96u l=0.18u
MI14-M_u3 net51 net90 VDD VDD p w=0.685u l=0.18u
MI20-M_u3 net84 SN VDD VDD p w=0.685u l=0.18u
MI17 net61 D net44 VDD p w=1.37u l=0.18u
MI52 net55 INCPB net47 VDD p w=1.34u l=0.18u
MI54 net51 INCP net47 VDD p w=0.42u l=0.18u
MI45 net64 INCPB net68 VDD p w=0.42u l=0.18u
MI43 net68 net55 VDD VDD p w=0.42u l=0.18u
MI18 net44 INCP net64 VDD p w=0.92u l=0.18u
MI19 VDD net84 net61 VDD p w=1.37u l=0.18u
.ends
.subckt DFKSND1BWP7T D CP SN Q QN VDD VSS 
MI15 net44 D VSS VSS n w=1u l=0.18u
MI12 net64 INCPB net44 VSS n w=0.94u l=0.18u
MI47 net64 INCP net56 VSS n w=0.42u l=0.18u
MI48 net56 net55 VSS VSS n w=0.42u l=0.18u
MI55 net51 INCPB net47 VSS n w=0.42u l=0.18u
MI50 net55 INCP net47 VSS n w=0.91u l=0.18u
MI16 net44 net84 VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net51 VSS VSS n w=0.94u l=0.18u
MI27-M_u2 Q net90 VSS VSS n w=1u l=0.18u
MI53-M_u2 net90 net47 VSS VSS n w=1u l=0.18u
MI13-M_u2 net55 net64 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net51 net90 VSS VSS n w=0.5u l=0.18u
MI20-M_u2 net84 SN VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net51 VDD VDD p w=1.37u l=0.18u
MI27-M_u3 Q net90 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 net90 net47 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 net55 net64 VDD VDD p w=0.96u l=0.18u
MI14-M_u3 net51 net90 VDD VDD p w=0.685u l=0.18u
MI20-M_u3 net84 SN VDD VDD p w=0.685u l=0.18u
MI17 net61 D net44 VDD p w=1.37u l=0.18u
MI52 net55 INCPB net47 VDD p w=1.34u l=0.18u
MI54 net51 INCP net47 VDD p w=0.42u l=0.18u
MI45 net64 INCPB net68 VDD p w=0.42u l=0.18u
MI43 net68 net55 VDD VDD p w=0.42u l=0.18u
MI18 net44 INCP net64 VDD p w=0.92u l=0.18u
MI19 VDD net84 net61 VDD p w=1.37u l=0.18u
.ends
.subckt DFKSND2BWP7T D CP SN Q QN VDD VSS 
MI15 net44 D VSS VSS n w=1u l=0.18u
MI12 net64 INCPB net44 VSS n w=0.94u l=0.18u
MI47 net64 INCP net56 VSS n w=0.42u l=0.18u
MI48 net56 net55 VSS VSS n w=0.42u l=0.18u
MI55 net062 INCPB net47 VSS n w=0.42u l=0.18u
MI50 net55 INCP net47 VSS n w=0.91u l=0.18u
MI16 net44 net84 VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29_0-M_u2 QN net062 VSS VSS n w=1u l=0.18u
MI29_1-M_u2 QN net062 VSS VSS n w=1u l=0.18u
MI27_0-M_u2 Q net90 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q net90 VSS VSS n w=1u l=0.18u
MI53-M_u2 net90 net47 VSS VSS n w=1u l=0.18u
MI13-M_u2 net55 net64 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net062 net90 VSS VSS n w=1u l=0.18u
MI20-M_u2 net84 SN VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29_0-M_u3 QN net062 VDD VDD p w=1.3u l=0.18u
MI29_1-M_u3 QN net062 VDD VDD p w=1.3u l=0.18u
MI27_0-M_u3 Q net90 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q net90 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 net90 net47 VDD VDD p w=1.23u l=0.18u
MI13-M_u3 net55 net64 VDD VDD p w=0.96u l=0.18u
MI14-M_u3 net062 net90 VDD VDD p w=1.37u l=0.18u
MI20-M_u3 net84 SN VDD VDD p w=0.685u l=0.18u
MI17 net61 D net44 VDD p w=1.37u l=0.18u
MI52 net55 INCPB net47 VDD p w=1.34u l=0.18u
MI54 net062 INCP net47 VDD p w=0.42u l=0.18u
MI45 net64 INCPB net68 VDD p w=0.42u l=0.18u
MI43 net68 net55 VDD VDD p w=0.42u l=0.18u
MI18 net44 INCP net64 VDD p w=0.92u l=0.18u
MI19 VDD net84 net61 VDD p w=1.37u l=0.18u
.ends
.subckt DFNCND0BWP7T D CPN CDN Q QN VDD VSS 
MI4 net52 net66 VSS VSS n w=1u l=0.18u
MI15 d1 INCPB net37 VSS n w=0.91u l=0.18u
MI5 d0 D net52 VSS n w=1u l=0.18u
MI18 d3 net66 net37 VSS n w=0.42u l=0.18u
MI47 d0 INCPB net59 VSS n w=0.42u l=0.18u
MI48 net59 CDN net62 VSS n w=0.42u l=0.18u
MI49 net62 d1 VSS VSS n w=0.42u l=0.18u
MI60-M_u4 XI60-net6 CDN VSS VSS n w=0.97u l=0.18u
MI60-M_u3 d2 net37 XI60-net6 VSS n w=0.97u l=0.18u
MI32-M_u2 net66 INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN d3 VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q d2 VSS VSS n w=0.5u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 d3 d2 VSS VSS n w=0.42u l=0.18u
MI60-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI60-M_u1 d2 net37 VDD VDD p w=1.31u l=0.18u
MI32-M_u3 net66 INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN d3 VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q d2 VDD VDD p w=0.685u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI14-M_u3 d3 d2 VDD VDD p w=0.6u l=0.18u
MI6 d0 D net85 VDD p w=1.27u l=0.18u
MI7 net85 INCPB VDD VDD p w=1.27u l=0.18u
MI16 d1 net66 net37 VDD p w=0.62u l=0.18u
MI17 d3 INCPB net37 VDD p w=0.42u l=0.18u
MI45 d0 net66 net98 VDD p w=0.42u l=0.18u
MI43 net98 d1 VDD VDD p w=0.42u l=0.18u
MI44 net98 CDN VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFNCND1BWP7T D CPN CDN Q QN VDD VSS 
MI4 net52 net66 VSS VSS n w=1u l=0.18u
MI15 d1 INCPB net37 VSS n w=0.91u l=0.18u
MI5 d0 D net52 VSS n w=1u l=0.18u
MI18 d3 net66 net37 VSS n w=0.42u l=0.18u
MI47 d0 INCPB net59 VSS n w=0.42u l=0.18u
MI48 net59 CDN net62 VSS n w=0.42u l=0.18u
MI49 net62 d1 VSS VSS n w=0.42u l=0.18u
MI60-M_u4 XI60-net6 CDN VSS VSS n w=0.97u l=0.18u
MI60-M_u3 d2 net37 XI60-net6 VSS n w=0.97u l=0.18u
MI32-M_u2 net66 INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN d3 VSS VSS n w=0.94u l=0.18u
MI27-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 d3 d2 VSS VSS n w=0.42u l=0.18u
MI60-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI60-M_u1 d2 net37 VDD VDD p w=1.37u l=0.18u
MI32-M_u3 net66 INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN d3 VDD VDD p w=0.835u l=0.18u
MI27-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI14-M_u3 d3 d2 VDD VDD p w=0.6u l=0.18u
MI6 d0 D net85 VDD p w=1.27u l=0.18u
MI7 net85 INCPB VDD VDD p w=1.27u l=0.18u
MI16 d1 net66 net37 VDD p w=0.62u l=0.18u
MI17 d3 INCPB net37 VDD p w=0.42u l=0.18u
MI45 d0 net66 net98 VDD p w=0.42u l=0.18u
MI43 net98 d1 VDD VDD p w=0.42u l=0.18u
MI44 net98 CDN VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFNCND2BWP7T D CPN CDN Q QN VDD VSS 
MI4 net52 net66 VSS VSS n w=1u l=0.18u
MI15 d1 INCPB net37 VSS n w=0.91u l=0.18u
MI5 d0 D net52 VSS n w=1u l=0.18u
MI18 d3 net66 net37 VSS n w=0.42u l=0.18u
MI47 d0 INCPB net59 VSS n w=0.42u l=0.18u
MI48 net59 CDN net62 VSS n w=0.42u l=0.18u
MI49 net62 d1 VSS VSS n w=0.42u l=0.18u
MI60-M_u4 XI60-net6 CDN VSS VSS n w=0.97u l=0.18u
MI60-M_u3 d2 net37 XI60-net6 VSS n w=0.97u l=0.18u
MI32-M_u2 net66 INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI29_0-M_u2 QN d3 VSS VSS n w=1u l=0.18u
MI29_1-M_u2 QN d3 VSS VSS n w=1u l=0.18u
MI27_0-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 d3 d2 VSS VSS n w=0.97u l=0.18u
MI60-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI60-M_u1 d2 net37 VDD VDD p w=1.23u l=0.18u
MI32-M_u3 net66 INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI29_0-M_u3 QN d3 VDD VDD p w=1.3u l=0.18u
MI29_1-M_u3 QN d3 VDD VDD p w=1.3u l=0.18u
MI27_0-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI14-M_u3 d3 d2 VDD VDD p w=0.97u l=0.18u
MI6 d0 D net85 VDD p w=1.27u l=0.18u
MI7 net85 INCPB VDD VDD p w=1.27u l=0.18u
MI16 d1 net66 net37 VDD p w=0.62u l=0.18u
MI17 d3 INCPB net37 VDD p w=0.42u l=0.18u
MI45 d0 net66 net98 VDD p w=0.42u l=0.18u
MI43 net98 d1 VDD VDD p w=0.42u l=0.18u
MI44 net98 CDN VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFND0BWP7T D CPN Q QN VDD VSS 
MI4 net43 net55 VSS VSS n w=0.905u l=0.18u
MI5 d0 D net43 VSS n w=1u l=0.18u
MI47 d0 INCPB net50 VSS n w=0.42u l=0.18u
MI48 net50 d1 VSS VSS n w=0.42u l=0.18u
MI55 net67 net55 d2 VSS n w=0.42u l=0.18u
MI50 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI32-M_u2 net55 INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net67 VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI53-M_u2 d3 d2 VSS VSS n w=0.5u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net67 d3 VSS VSS n w=0.5u l=0.18u
MI32-M_u3 net55 INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net67 VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI53-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.97u l=0.18u
MI14-M_u3 net67 d3 VDD VDD p w=0.685u l=0.18u
MI6 d0 D net66 VDD p w=0.94u l=0.18u
MI7 net66 INCPB VDD VDD p w=0.84u l=0.18u
MI52 d1 net55 d2 VDD p w=1.34u l=0.18u
MI54 net67 INCPB d2 VDD p w=0.42u l=0.18u
MI45 d0 net55 net84 VDD p w=0.42u l=0.18u
MI43 net84 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFND1BWP7T D CPN Q QN VDD VSS 
MI4 net43 net55 VSS VSS n w=0.905u l=0.18u
MI5 d0 D net43 VSS n w=1u l=0.18u
MI47 d0 INCPB net50 VSS n w=0.42u l=0.18u
MI48 net50 d1 VSS VSS n w=0.42u l=0.18u
MI55 net67 net55 d2 VSS n w=0.42u l=0.18u
MI50 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI32-M_u2 net55 INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net67 VSS VSS n w=0.94u l=0.18u
MI27-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI53-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net67 d3 VSS VSS n w=0.5u l=0.18u
MI32-M_u3 net55 INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net67 VDD VDD p w=1.37u l=0.18u
MI27-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.97u l=0.18u
MI14-M_u3 net67 d3 VDD VDD p w=0.685u l=0.18u
MI6 d0 D net66 VDD p w=0.94u l=0.18u
MI7 net66 INCPB VDD VDD p w=0.84u l=0.18u
MI52 d1 net55 d2 VDD p w=1.34u l=0.18u
MI54 net67 INCPB d2 VDD p w=0.42u l=0.18u
MI45 d0 net55 net84 VDD p w=0.42u l=0.18u
MI43 net84 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFND2BWP7T D CPN Q QN VDD VSS 
MI4 net43 net55 VSS VSS n w=0.905u l=0.18u
MI5 d0 D net43 VSS n w=1u l=0.18u
MI47 d0 INCPB net50 VSS n w=0.42u l=0.18u
MI48 net50 d1 VSS VSS n w=0.42u l=0.18u
MI55 net053 net55 d2 VSS n w=0.42u l=0.18u
MI50 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI32-M_u2 net55 INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI29_0-M_u2 QN net053 VSS VSS n w=1u l=0.18u
MI29_1-M_u2 QN net053 VSS VSS n w=1u l=0.18u
MI27_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI53-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI14-M_u2 net053 d3 VSS VSS n w=1u l=0.18u
MI32-M_u3 net55 INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI29_0-M_u3 QN net053 VDD VDD p w=1.3u l=0.18u
MI29_1-M_u3 QN net053 VDD VDD p w=1.3u l=0.18u
MI27_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 d3 d2 VDD VDD p w=1.23u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.97u l=0.18u
MI14-M_u3 net053 d3 VDD VDD p w=1.37u l=0.18u
MI6 d0 D net66 VDD p w=0.94u l=0.18u
MI7 net66 INCPB VDD VDD p w=0.84u l=0.18u
MI52 d1 net55 d2 VDD p w=1.34u l=0.18u
MI54 net053 INCPB d2 VDD p w=0.42u l=0.18u
MI45 d0 net55 net84 VDD p w=0.42u l=0.18u
MI43 net84 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFNSND0BWP7T D CPN SDN Q QN VDD VSS 
MI19 net57 net68 VSS VSS n w=1u l=0.18u
MI20 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI21 d0 D net57 VSS n w=1u l=0.18u
MI22 d4 net68 d2 VSS n w=0.42u l=0.18u
MI23 d0 INCPB net44 VSS n w=0.42u l=0.18u
MI24 net44 d1 VSS VSS n w=0.42u l=0.18u
MI31-M_u4 XI31-net6 d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u3 d4 SDN XI31-net6 VSS n w=0.5u l=0.18u
MI32-M_u4 XI32-net6 SDN VSS VSS n w=0.54u l=0.18u
MI32-M_u3 d1 d0 XI32-net6 VSS n w=0.54u l=0.18u
MI25-M_u2 d3 d2 VSS VSS n w=0.5u l=0.18u
MI40-M_u2 net68 INCPB VSS VSS n w=0.5u l=0.18u
MI55-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI57-M_u2 QN d4 VSS VSS n w=0.5u l=0.18u
MI60-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u2 d4 d3 VDD VDD p w=0.685u l=0.18u
MI31-M_u1 d4 SDN VDD VDD p w=0.685u l=0.18u
MI32-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI32-M_u1 d1 d0 VDD VDD p w=0.97u l=0.18u
MI25-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI40-M_u3 net68 INCPB VDD VDD p w=0.685u l=0.18u
MI55-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI57-M_u3 QN d4 VDD VDD p w=0.685u l=0.18u
MI60-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI26 d0 D net82 VDD p w=1.27u l=0.18u
MI28 net82 INCPB VDD VDD p w=1.27u l=0.18u
MI30 d1 net68 d2 VDD p w=1.34u l=0.18u
MI33 d4 INCPB d2 VDD p w=0.42u l=0.18u
MI34 d0 net68 net65 VDD p w=0.42u l=0.18u
MI35 net65 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFNSND1BWP7T D CPN SDN Q QN VDD VSS 
MI19 net57 net68 VSS VSS n w=1u l=0.18u
MI20 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI21 d0 D net57 VSS n w=1u l=0.18u
MI22 d4 net68 d2 VSS n w=0.42u l=0.18u
MI23 d0 INCPB net44 VSS n w=0.42u l=0.18u
MI24 net44 d1 VSS VSS n w=0.42u l=0.18u
MI31-M_u4 XI31-net6 d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u3 d4 SDN XI31-net6 VSS n w=0.5u l=0.18u
MI32-M_u4 XI32-net6 SDN VSS VSS n w=0.54u l=0.18u
MI32-M_u3 d1 d0 XI32-net6 VSS n w=0.54u l=0.18u
MI25-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI40-M_u2 net68 INCPB VSS VSS n w=0.5u l=0.18u
MI55-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI57-M_u2 QN d4 VSS VSS n w=1u l=0.18u
MI60-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI31-M_u2 d4 d3 VDD VDD p w=0.685u l=0.18u
MI31-M_u1 d4 SDN VDD VDD p w=0.685u l=0.18u
MI32-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI32-M_u1 d1 d0 VDD VDD p w=0.97u l=0.18u
MI25-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI40-M_u3 net68 INCPB VDD VDD p w=0.685u l=0.18u
MI55-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI57-M_u3 QN d4 VDD VDD p w=1.37u l=0.18u
MI60-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI26 d0 D net82 VDD p w=1.27u l=0.18u
MI28 net82 INCPB VDD VDD p w=1.27u l=0.18u
MI30 d1 net68 d2 VDD p w=1.34u l=0.18u
MI33 d4 INCPB d2 VDD p w=0.42u l=0.18u
MI34 d0 net68 net65 VDD p w=0.42u l=0.18u
MI35 net65 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFNSND2BWP7T D CPN SDN Q QN VDD VSS 
MI19 net57 net68 VSS VSS n w=1u l=0.18u
MI20 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI21 d0 D net57 VSS n w=1u l=0.18u
MI22 d4 net68 d2 VSS n w=0.42u l=0.18u
MI23 d0 INCPB net44 VSS n w=0.42u l=0.18u
MI24 net44 d1 VSS VSS n w=0.42u l=0.18u
MI31-M_u4 XI31-net6 d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u3 d4 SDN XI31-net6 VSS n w=0.5u l=0.18u
MI32-M_u4 XI32-net6 SDN VSS VSS n w=0.54u l=0.18u
MI32-M_u3 d1 d0 XI32-net6 VSS n w=0.54u l=0.18u
MI25-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI40-M_u2 net68 INCPB VSS VSS n w=0.5u l=0.18u
MI55-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI57_0-M_u2 QN d4 VSS VSS n w=1u l=0.18u
MI57_1-M_u2 QN d4 VSS VSS n w=1u l=0.18u
MI60_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI60_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI31-M_u2 d4 d3 VDD VDD p w=0.685u l=0.18u
MI31-M_u1 d4 SDN VDD VDD p w=0.685u l=0.18u
MI32-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI32-M_u1 d1 d0 VDD VDD p w=0.97u l=0.18u
MI25-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI40-M_u3 net68 INCPB VDD VDD p w=0.685u l=0.18u
MI55-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI57_0-M_u3 QN d4 VDD VDD p w=1.37u l=0.18u
MI57_1-M_u3 QN d4 VDD VDD p w=1.37u l=0.18u
MI60_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI60_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI26 d0 D net82 VDD p w=1.27u l=0.18u
MI28 net82 INCPB VDD VDD p w=1.27u l=0.18u
MI30 d1 net68 d2 VDD p w=1.34u l=0.18u
MI33 d4 INCPB d2 VDD p w=0.42u l=0.18u
MI34 d0 net68 net65 VDD p w=0.42u l=0.18u
MI35 net65 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFQD0BWP7T D CP Q VDD VSS 
MI4 net43 INCPB VSS VSS n w=0.94u l=0.18u
MI5 P000 D net43 VSS n w=0.94u l=0.18u
MI47 P000 INCP net50 VSS n w=0.42u l=0.18u
MI48 net50 P0001 VSS VSS n w=0.42u l=0.18u
MI55 net052 INCPB N0028 VSS n w=0.42u l=0.18u
MI50 P0001 INCP N0028 VSS n w=0.91u l=0.18u
MI56-M_u2 net052 P0003 VSS VSS n w=0.42u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q P0003 VSS VSS n w=0.5u l=0.18u
MI53-M_u2 P0003 N0028 VSS VSS n w=0.5u l=0.18u
MI13-M_u2 P0001 P000 VSS VSS n w=0.54u l=0.18u
MI56-M_u3 net052 P0003 VDD VDD p w=0.42u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q P0003 VDD VDD p w=0.685u l=0.18u
MI53-M_u3 P0003 N0028 VDD VDD p w=0.685u l=0.18u
MI13-M_u3 P0001 P000 VDD VDD p w=0.96u l=0.18u
MI6 P000 D net74 VDD p w=0.92u l=0.18u
MI7 net74 INCP VDD VDD p w=0.92u l=0.18u
MI52 P0001 INCPB N0028 VDD p w=1.34u l=0.18u
MI54 net052 INCP N0028 VDD p w=0.42u l=0.18u
MI45 P000 INCPB net86 VDD p w=0.42u l=0.18u
MI43 net86 P0001 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFQD1BWP7T D CP Q VDD VSS 
MI4 net43 INCPB VSS VSS n w=0.94u l=0.18u
MI5 P000 D net43 VSS n w=0.94u l=0.18u
MI47 P000 INCP net50 VSS n w=0.42u l=0.18u
MI48 net50 P0001 VSS VSS n w=0.42u l=0.18u
MI55 net052 INCPB N0028 VSS n w=0.42u l=0.18u
MI50 P0001 INCP N0028 VSS n w=0.91u l=0.18u
MI56-M_u2 net052 P0003 VSS VSS n w=0.42u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q P0003 VSS VSS n w=1u l=0.18u
MI53-M_u2 P0003 N0028 VSS VSS n w=1u l=0.18u
MI13-M_u2 P0001 P000 VSS VSS n w=0.54u l=0.18u
MI56-M_u3 net052 P0003 VDD VDD p w=0.42u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q P0003 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 P0003 N0028 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 P0001 P000 VDD VDD p w=0.96u l=0.18u
MI6 P000 D net74 VDD p w=0.92u l=0.18u
MI7 net74 INCP VDD VDD p w=0.92u l=0.18u
MI52 P0001 INCPB N0028 VDD p w=1.34u l=0.18u
MI54 net052 INCP N0028 VDD p w=0.42u l=0.18u
MI45 P000 INCPB net86 VDD p w=0.42u l=0.18u
MI43 net86 P0001 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFQD2BWP7T D CP Q VDD VSS 
MI4 net43 INCPB VSS VSS n w=0.94u l=0.18u
MI5 P000 D net43 VSS n w=0.94u l=0.18u
MI47 P000 INCP net50 VSS n w=0.42u l=0.18u
MI48 net50 P0001 VSS VSS n w=0.42u l=0.18u
MI55 net052 INCPB N0028 VSS n w=0.42u l=0.18u
MI50 P0001 INCP N0028 VSS n w=0.91u l=0.18u
MI56-M_u2 net052 P0003 VSS VSS n w=0.42u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27_0-M_u2 Q P0003 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q P0003 VSS VSS n w=1u l=0.18u
MI53-M_u2 P0003 N0028 VSS VSS n w=1u l=0.18u
MI13-M_u2 P0001 P000 VSS VSS n w=0.54u l=0.18u
MI56-M_u3 net052 P0003 VDD VDD p w=0.42u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27_0-M_u3 Q P0003 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q P0003 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 P0003 N0028 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 P0001 P000 VDD VDD p w=0.96u l=0.18u
MI6 P000 D net74 VDD p w=0.92u l=0.18u
MI7 net74 INCP VDD VDD p w=0.92u l=0.18u
MI52 P0001 INCPB N0028 VDD p w=1.34u l=0.18u
MI54 net052 INCP N0028 VDD p w=0.42u l=0.18u
MI45 P000 INCPB net86 VDD p w=0.42u l=0.18u
MI43 net86 P0001 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFSND0BWP7T D CP SDN Q QN VDD VSS 
MI19 net57 INCPB VSS VSS n w=0.94u l=0.18u
MI20 d1 INCP d2 VSS n w=0.91u l=0.18u
MI21 net052 D net57 VSS n w=0.94u l=0.18u
MI22 d4 INCPB d2 VSS n w=0.42u l=0.18u
MI23 net052 INCP net44 VSS n w=0.42u l=0.18u
MI24 net44 d1 VSS VSS n w=0.42u l=0.18u
MI31-M_u4 XI31-net6 d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u3 d4 SDN XI31-net6 VSS n w=0.5u l=0.18u
MI32-M_u4 XI32-net6 SDN VSS VSS n w=0.54u l=0.18u
MI32-M_u3 d1 net052 XI32-net6 VSS n w=0.54u l=0.18u
MI25-M_u2 d3 d2 VSS VSS n w=0.5u l=0.18u
MI40-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI55-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI57-M_u2 QN d4 VSS VSS n w=0.5u l=0.18u
MI60-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u2 d4 d3 VDD VDD p w=0.685u l=0.18u
MI31-M_u1 d4 SDN VDD VDD p w=0.685u l=0.18u
MI32-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI32-M_u1 d1 net052 VDD VDD p w=0.97u l=0.18u
MI25-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI40-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI55-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI57-M_u3 QN d4 VDD VDD p w=0.685u l=0.18u
MI60-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI26 net052 D net82 VDD p w=0.92u l=0.18u
MI28 net82 INCP VDD VDD p w=0.92u l=0.18u
MI30 d1 INCPB d2 VDD p w=1.34u l=0.18u
MI33 d4 INCP d2 VDD p w=0.42u l=0.18u
MI34 net052 INCPB net65 VDD p w=0.42u l=0.18u
MI35 net65 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFSND1BWP7T D CP SDN Q QN VDD VSS 
MI19 net57 INCPB VSS VSS n w=0.94u l=0.18u
MI20 d1 INCP d2 VSS n w=0.91u l=0.18u
MI21 net052 D net57 VSS n w=0.94u l=0.18u
MI22 d4 INCPB d2 VSS n w=0.42u l=0.18u
MI23 net052 INCP net44 VSS n w=0.42u l=0.18u
MI24 net44 d1 VSS VSS n w=0.42u l=0.18u
MI31-M_u4 XI31-net6 d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u3 d4 SDN XI31-net6 VSS n w=0.5u l=0.18u
MI32-M_u4 XI32-net6 SDN VSS VSS n w=0.54u l=0.18u
MI32-M_u3 d1 net052 XI32-net6 VSS n w=0.54u l=0.18u
MI25-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI40-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI55-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI57-M_u2 QN d4 VSS VSS n w=1u l=0.18u
MI60-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI31-M_u2 d4 d3 VDD VDD p w=0.685u l=0.18u
MI31-M_u1 d4 SDN VDD VDD p w=0.685u l=0.18u
MI32-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI32-M_u1 d1 net052 VDD VDD p w=0.97u l=0.18u
MI25-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI40-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI55-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI57-M_u3 QN d4 VDD VDD p w=1.37u l=0.18u
MI60-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI26 net052 D net82 VDD p w=0.92u l=0.18u
MI28 net82 INCP VDD VDD p w=0.92u l=0.18u
MI30 d1 INCPB d2 VDD p w=1.34u l=0.18u
MI33 d4 INCP d2 VDD p w=0.42u l=0.18u
MI34 net052 INCPB net65 VDD p w=0.42u l=0.18u
MI35 net65 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFSND2BWP7T D CP SDN Q QN VDD VSS 
MI19 net57 INCPB VSS VSS n w=0.94u l=0.18u
MI20 d1 INCP d2 VSS n w=0.91u l=0.18u
MI21 net052 D net57 VSS n w=0.94u l=0.18u
MI22 d4 INCPB d2 VSS n w=0.42u l=0.18u
MI23 net052 INCP net44 VSS n w=0.42u l=0.18u
MI24 net44 d1 VSS VSS n w=0.42u l=0.18u
MI31-M_u4 XI31-net6 d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u3 d4 SDN XI31-net6 VSS n w=0.5u l=0.18u
MI32-M_u4 XI32-net6 SDN VSS VSS n w=0.54u l=0.18u
MI32-M_u3 d1 net052 XI32-net6 VSS n w=0.54u l=0.18u
MI25-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI40-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI55-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI57_0-M_u2 QN d4 VSS VSS n w=1u l=0.18u
MI57_1-M_u2 QN d4 VSS VSS n w=1u l=0.18u
MI60_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI60_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI31-M_u2 d4 d3 VDD VDD p w=0.685u l=0.18u
MI31-M_u1 d4 SDN VDD VDD p w=0.685u l=0.18u
MI32-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI32-M_u1 d1 net052 VDD VDD p w=0.97u l=0.18u
MI25-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI40-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI55-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI57_0-M_u3 QN d4 VDD VDD p w=1.37u l=0.18u
MI57_1-M_u3 QN d4 VDD VDD p w=1.37u l=0.18u
MI60_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI60_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI26 net052 D net82 VDD p w=0.92u l=0.18u
MI28 net82 INCP VDD VDD p w=0.92u l=0.18u
MI30 d1 INCPB d2 VDD p w=1.34u l=0.18u
MI33 d4 INCP d2 VDD p w=0.42u l=0.18u
MI34 net052 INCPB net65 VDD p w=0.42u l=0.18u
MI35 net65 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFSNQD1BWP7T D CP SDN Q VDD VSS 
MI19 net57 INCPB VSS VSS n w=0.94u l=0.18u
MI20 d1 INCP d2 VSS n w=0.91u l=0.18u
MI21 net052 D net57 VSS n w=0.94u l=0.18u
MI22 net056 INCPB d2 VSS n w=0.42u l=0.18u
MI23 net052 INCP net44 VSS n w=0.42u l=0.18u
MI24 net44 d1 VSS VSS n w=0.42u l=0.18u
MI31-M_u4 XI31-net6 d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u3 net056 SDN XI31-net6 VSS n w=0.5u l=0.18u
MI32-M_u4 XI32-net6 SDN VSS VSS n w=0.54u l=0.18u
MI32-M_u3 d1 net052 XI32-net6 VSS n w=0.54u l=0.18u
MI25-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI40-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI55-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI60-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI31-M_u2 net056 d3 VDD VDD p w=0.685u l=0.18u
MI31-M_u1 net056 SDN VDD VDD p w=0.685u l=0.18u
MI32-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI32-M_u1 d1 net052 VDD VDD p w=0.97u l=0.18u
MI25-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI40-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI55-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI60-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI26 net052 D net82 VDD p w=0.92u l=0.18u
MI28 net82 INCP VDD VDD p w=0.92u l=0.18u
MI30 d1 INCPB d2 VDD p w=1.34u l=0.18u
MI33 net056 INCP d2 VDD p w=0.42u l=0.18u
MI34 net052 INCPB net65 VDD p w=0.42u l=0.18u
MI35 net65 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFSNQD2BWP7T D CP SDN Q VDD VSS 
MI19 net57 INCPB VSS VSS n w=0.94u l=0.18u
MI20 d1 INCP d2 VSS n w=0.91u l=0.18u
MI21 net052 D net57 VSS n w=0.94u l=0.18u
MI22 net056 INCPB d2 VSS n w=0.42u l=0.18u
MI23 net052 INCP net44 VSS n w=0.42u l=0.18u
MI24 net44 d1 VSS VSS n w=0.42u l=0.18u
MI31-M_u4 XI31-net6 d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u3 net056 SDN XI31-net6 VSS n w=0.5u l=0.18u
MI32-M_u4 XI32-net6 SDN VSS VSS n w=0.54u l=0.18u
MI32-M_u3 d1 net052 XI32-net6 VSS n w=0.54u l=0.18u
MI25-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI40-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI55-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI60_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI60_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI31-M_u2 net056 d3 VDD VDD p w=0.685u l=0.18u
MI31-M_u1 net056 SDN VDD VDD p w=0.685u l=0.18u
MI32-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI32-M_u1 d1 net052 VDD VDD p w=0.97u l=0.18u
MI25-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI40-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI55-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI60_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI60_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI26 net052 D net82 VDD p w=0.92u l=0.18u
MI28 net82 INCP VDD VDD p w=0.92u l=0.18u
MI30 d1 INCPB d2 VDD p w=1.34u l=0.18u
MI33 net056 INCP d2 VDD p w=0.42u l=0.18u
MI34 net052 INCPB net65 VDD p w=0.42u l=0.18u
MI35 net65 d1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt DFXD0BWP7T DA DB SA CP Q QN VDD VSS 
MI47 net66 INCP net75 VSS n w=0.42u l=0.18u
MI26 net66 INCPB net57 VSS n w=0.91u l=0.18u
MI30 net53 DB VSS VSS n w=1u l=0.18u
MI33 net57 SA net63 VSS n w=0.525u l=0.18u
MI18 net76 INCP net68 VSS n w=0.91u l=0.18u
MI17 net72 INCPB net68 VSS n w=0.42u l=0.18u
MI48 net75 net76 VSS VSS n w=0.42u l=0.18u
MI28 net63 DA VSS VSS n w=0.525u l=0.18u
MI34 net57 net84 net53 VSS n w=1u l=0.18u
MI24-M_u2 net72 net90 VSS VSS n w=0.42u l=0.18u
MI23-M_u2 net76 net66 VSS VSS n w=0.54u l=0.18u
MI22-M_u2 net90 net68 VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q net90 VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net72 VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI35-M_u2 net84 SA VSS VSS n w=0.5u l=0.18u
MI24-M_u3 net72 net90 VDD VDD p w=0.685u l=0.18u
MI23-M_u3 net76 net66 VDD VDD p w=0.96u l=0.18u
MI22-M_u3 net90 net68 VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q net90 VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net72 VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI35-M_u3 net84 SA VDD VDD p w=0.685u l=0.18u
MI21 net72 INCP net68 VDD p w=0.42u l=0.18u
MI20 net76 INCPB net68 VDD p w=1.34u l=0.18u
MI43 net116 net76 VDD VDD p w=0.42u l=0.18u
MI45 net66 INCPB net116 VDD p w=0.42u l=0.18u
MI40 net110 DA VDD VDD p w=0.725u l=0.18u
MI36 net57 net84 net110 VDD p w=0.725u l=0.18u
MI37 net104 DB VDD VDD p w=1.23u l=0.18u
MI38 net57 SA net104 VDD p w=1.095u l=0.18u
MI39 net66 INCP net57 VDD p w=0.95u l=0.18u
.ends
.subckt DFXD1BWP7T DA DB SA CP Q QN VDD VSS 
MI47 net66 INCP net75 VSS n w=0.42u l=0.18u
MI26 net66 INCPB net57 VSS n w=0.91u l=0.18u
MI30 net53 DB VSS VSS n w=1u l=0.18u
MI33 net57 SA net63 VSS n w=0.525u l=0.18u
MI18 net76 INCP net68 VSS n w=0.91u l=0.18u
MI17 net72 INCPB net68 VSS n w=0.42u l=0.18u
MI48 net75 net76 VSS VSS n w=0.42u l=0.18u
MI28 net63 DA VSS VSS n w=0.525u l=0.18u
MI34 net57 net84 net53 VSS n w=1u l=0.18u
MI24-M_u2 net72 net90 VSS VSS n w=0.42u l=0.18u
MI23-M_u2 net76 net66 VSS VSS n w=0.54u l=0.18u
MI22-M_u2 net90 net68 VSS VSS n w=1u l=0.18u
MI27-M_u2 Q net90 VSS VSS n w=1u l=0.18u
MI29-M_u2 QN net72 VSS VSS n w=0.94u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI35-M_u2 net84 SA VSS VSS n w=0.5u l=0.18u
MI24-M_u3 net72 net90 VDD VDD p w=0.685u l=0.18u
MI23-M_u3 net76 net66 VDD VDD p w=0.96u l=0.18u
MI22-M_u3 net90 net68 VDD VDD p w=1.37u l=0.18u
MI27-M_u3 Q net90 VDD VDD p w=1.37u l=0.18u
MI29-M_u3 QN net72 VDD VDD p w=1.37u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI35-M_u3 net84 SA VDD VDD p w=0.685u l=0.18u
MI21 net72 INCP net68 VDD p w=0.42u l=0.18u
MI20 net76 INCPB net68 VDD p w=1.34u l=0.18u
MI43 net116 net76 VDD VDD p w=0.42u l=0.18u
MI45 net66 INCPB net116 VDD p w=0.42u l=0.18u
MI40 net110 DA VDD VDD p w=0.725u l=0.18u
MI36 net57 net84 net110 VDD p w=0.725u l=0.18u
MI37 net104 DB VDD VDD p w=1.23u l=0.18u
MI38 net57 SA net104 VDD p w=1.095u l=0.18u
MI39 net66 INCP net57 VDD p w=0.95u l=0.18u
.ends
.subckt DFXD2BWP7T DA DB SA CP Q QN VDD VSS 
MI47 net66 INCP net75 VSS n w=0.42u l=0.18u
MI26 net66 INCPB net57 VSS n w=0.91u l=0.18u
MI30 net53 DB VSS VSS n w=1u l=0.18u
MI33 net57 SA net63 VSS n w=0.525u l=0.18u
MI18 net76 INCP net68 VSS n w=0.91u l=0.18u
MI17 net72 INCPB net68 VSS n w=0.42u l=0.18u
MI48 net75 net76 VSS VSS n w=0.42u l=0.18u
MI28 net63 DA VSS VSS n w=0.525u l=0.18u
MI34 net57 net84 net53 VSS n w=1u l=0.18u
MI24-M_u2 net72 net90 VSS VSS n w=1u l=0.18u
MI23-M_u2 net76 net66 VSS VSS n w=0.54u l=0.18u
MI22-M_u2 net90 net68 VSS VSS n w=1u l=0.18u
MI27_0-M_u2 Q net90 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q net90 VSS VSS n w=1u l=0.18u
MI29_0-M_u2 QN net72 VSS VSS n w=1u l=0.18u
MI29_1-M_u2 QN net72 VSS VSS n w=1u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI35-M_u2 net84 SA VSS VSS n w=0.5u l=0.18u
MI24-M_u3 net72 net90 VDD VDD p w=1.37u l=0.18u
MI23-M_u3 net76 net66 VDD VDD p w=0.96u l=0.18u
MI22-M_u3 net90 net68 VDD VDD p w=1.23u l=0.18u
MI27_0-M_u3 Q net90 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q net90 VDD VDD p w=1.37u l=0.18u
MI29_0-M_u3 QN net72 VDD VDD p w=1.3u l=0.18u
MI29_1-M_u3 QN net72 VDD VDD p w=1.3u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI35-M_u3 net84 SA VDD VDD p w=0.685u l=0.18u
MI21 net72 INCP net68 VDD p w=0.42u l=0.18u
MI20 net76 INCPB net68 VDD p w=1.34u l=0.18u
MI43 net116 net76 VDD VDD p w=0.42u l=0.18u
MI45 net66 INCPB net116 VDD p w=0.42u l=0.18u
MI40 net110 DA VDD VDD p w=0.725u l=0.18u
MI36 net57 net84 net110 VDD p w=0.725u l=0.18u
MI37 net104 DB VDD VDD p w=1.23u l=0.18u
MI38 net57 SA net104 VDD p w=1.095u l=0.18u
MI39 net66 INCP net57 VDD p w=0.95u l=0.18u
.ends
.subckt DFXQD1BWP7T DA DB SA CP Q VDD VSS 
MI47 net66 INCP net75 VSS n w=0.42u l=0.18u
MI26 net66 INCPB net57 VSS n w=0.91u l=0.18u
MI30 net53 DB VSS VSS n w=1u l=0.18u
MI33 net57 SA net63 VSS n w=0.525u l=0.18u
MI18 net76 INCP net68 VSS n w=0.91u l=0.18u
MI17 net72 INCPB net68 VSS n w=0.42u l=0.18u
MI48 net75 net76 VSS VSS n w=0.42u l=0.18u
MI28 net63 DA VSS VSS n w=0.525u l=0.18u
MI34 net57 net84 net53 VSS n w=1u l=0.18u
MI24-M_u2 net72 net90 VSS VSS n w=0.42u l=0.18u
MI23-M_u2 net76 net66 VSS VSS n w=0.54u l=0.18u
MI22-M_u2 net90 net68 VSS VSS n w=1u l=0.18u
MI27-M_u2 Q net90 VSS VSS n w=1u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI35-M_u2 net84 SA VSS VSS n w=0.5u l=0.18u
MI24-M_u3 net72 net90 VDD VDD p w=0.42u l=0.18u
MI23-M_u3 net76 net66 VDD VDD p w=0.96u l=0.18u
MI22-M_u3 net90 net68 VDD VDD p w=1.37u l=0.18u
MI27-M_u3 Q net90 VDD VDD p w=1.37u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI35-M_u3 net84 SA VDD VDD p w=0.685u l=0.18u
MI21 net72 INCP net68 VDD p w=0.42u l=0.18u
MI20 net76 INCPB net68 VDD p w=1.34u l=0.18u
MI43 net116 net76 VDD VDD p w=0.42u l=0.18u
MI45 net66 INCPB net116 VDD p w=0.42u l=0.18u
MI40 net110 DA VDD VDD p w=0.94u l=0.18u
MI36 net57 net84 net110 VDD p w=0.94u l=0.18u
MI37 net104 DB VDD VDD p w=1.23u l=0.18u
MI38 net57 SA net104 VDD p w=1.095u l=0.18u
MI39 net66 INCP net57 VDD p w=0.92u l=0.18u
.ends
.subckt DFXQD2BWP7T DA DB SA CP Q VDD VSS 
MI47 net66 INCP net75 VSS n w=0.42u l=0.18u
MI26 net66 INCPB net57 VSS n w=0.91u l=0.18u
MI30 net53 DB VSS VSS n w=1u l=0.18u
MI33 net57 SA net63 VSS n w=0.525u l=0.18u
MI18 net76 INCP net68 VSS n w=0.91u l=0.18u
MI17 net72 INCPB net68 VSS n w=0.42u l=0.18u
MI48 net75 net76 VSS VSS n w=0.42u l=0.18u
MI28 net63 DA VSS VSS n w=0.525u l=0.18u
MI34 net57 net84 net53 VSS n w=1u l=0.18u
MI24-M_u2 net72 net90 VSS VSS n w=0.42u l=0.18u
MI23-M_u2 net76 net66 VSS VSS n w=0.54u l=0.18u
MI22-M_u2 net90 net68 VSS VSS n w=1u l=0.18u
MI27_0-M_u2 Q net90 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q net90 VSS VSS n w=1u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI35-M_u2 net84 SA VSS VSS n w=0.5u l=0.18u
MI24-M_u3 net72 net90 VDD VDD p w=0.42u l=0.18u
MI23-M_u3 net76 net66 VDD VDD p w=0.96u l=0.18u
MI22-M_u3 net90 net68 VDD VDD p w=1.37u l=0.18u
MI27_0-M_u3 Q net90 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q net90 VDD VDD p w=1.37u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI35-M_u3 net84 SA VDD VDD p w=0.685u l=0.18u
MI21 net72 INCP net68 VDD p w=0.42u l=0.18u
MI20 net76 INCPB net68 VDD p w=1.34u l=0.18u
MI43 net116 net76 VDD VDD p w=0.42u l=0.18u
MI45 net66 INCPB net116 VDD p w=0.42u l=0.18u
MI40 net110 DA VDD VDD p w=0.94u l=0.18u
MI36 net57 net84 net110 VDD p w=0.94u l=0.18u
MI37 net104 DB VDD VDD p w=1.23u l=0.18u
MI38 net57 SA net104 VDD p w=1.095u l=0.18u
MI39 net66 INCP net57 VDD p w=0.92u l=0.18u
.ends
.subckt EDFCND0BWP7T D E CP CDN Q QN VDD VSS 
MI132 d0 INCPB net124 VSS n w=0.74u l=0.18u
MI133 net116 d3 VSS VSS n w=0.42u l=0.18u
MI49 net89 d1 VSS VSS n w=0.42u l=0.18u
MI48 net92 CDN net89 VSS n w=0.42u l=0.18u
MI47 d0 INCP net92 VSS n w=0.42u l=0.18u
MI18 d3 INCPB net98 VSS n w=0.42u l=0.18u
MI146 net124 E net088 VSS n w=0.57u l=0.18u
MI15 d1 INCP net98 VSS n w=0.91u l=0.18u
MI135 net088 D VSS VSS n w=0.57u l=0.18u
MI136 net124 net119 net116 VSS n w=0.42u l=0.18u
MI144-M_u4 XI144-net6 CDN VSS VSS n w=0.93u l=0.18u
MI144-M_u3 d2 net98 XI144-net6 VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI27-M_u2 Q d2 VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN d3 VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI14-M_u2 d3 d2 VSS VSS n w=0.42u l=0.18u
MI137-M_u2 net119 E VSS VSS n w=0.5u l=0.18u
MI144-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI144-M_u1 d2 net98 VDD VDD p w=1.03u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI27-M_u3 Q d2 VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN d3 VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI14-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI137-M_u3 net119 E VDD VDD p w=0.685u l=0.18u
MI44 net79 CDN VDD VDD p w=0.42u l=0.18u
MI43 net79 d1 VDD VDD p w=0.42u l=0.18u
MI45 d0 INCPB net79 VDD p w=0.42u l=0.18u
MI17 d3 INCP net98 VDD p w=0.42u l=0.18u
MI16 d1 INCPB net98 VDD p w=0.62u l=0.18u
MI138 d0 INCP net124 VDD p w=0.78u l=0.18u
MI139 net64 D VDD VDD p w=0.75u l=0.18u
MI141 net124 E net129 VDD p w=0.42u l=0.18u
MI140 net129 d3 VDD VDD p w=0.42u l=0.18u
MI145 net124 net119 net64 VDD p w=0.75u l=0.18u
.ends
.subckt EDFCND1BWP7T D E CP CDN Q QN VDD VSS 
MI132 d0 INCPB net124 VSS n w=0.74u l=0.18u
MI133 net116 d3 VSS VSS n w=0.42u l=0.18u
MI49 net89 d1 VSS VSS n w=0.42u l=0.18u
MI48 net92 CDN net89 VSS n w=0.42u l=0.18u
MI47 d0 INCP net92 VSS n w=0.42u l=0.18u
MI18 d3 INCPB net98 VSS n w=0.42u l=0.18u
MI146 net124 E net088 VSS n w=0.57u l=0.18u
MI15 d1 INCP net98 VSS n w=0.91u l=0.18u
MI135 net088 D VSS VSS n w=0.57u l=0.18u
MI136 net124 net119 net116 VSS n w=0.42u l=0.18u
MI144-M_u4 XI144-net6 CDN VSS VSS n w=0.93u l=0.18u
MI144-M_u3 d2 net98 XI144-net6 VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI27-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI29-M_u2 QN d3 VSS VSS n w=0.94u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI14-M_u2 d3 d2 VSS VSS n w=0.42u l=0.18u
MI137-M_u2 net119 E VSS VSS n w=0.5u l=0.18u
MI144-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI144-M_u1 d2 net98 VDD VDD p w=1.03u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI27-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI29-M_u3 QN d3 VDD VDD p w=1.37u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI14-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI137-M_u3 net119 E VDD VDD p w=0.685u l=0.18u
MI44 net79 CDN VDD VDD p w=0.42u l=0.18u
MI43 net79 d1 VDD VDD p w=0.42u l=0.18u
MI45 d0 INCPB net79 VDD p w=0.42u l=0.18u
MI17 d3 INCP net98 VDD p w=0.42u l=0.18u
MI16 d1 INCPB net98 VDD p w=0.62u l=0.18u
MI138 d0 INCP net124 VDD p w=0.78u l=0.18u
MI139 net64 D VDD VDD p w=0.75u l=0.18u
MI141 net124 E net129 VDD p w=0.42u l=0.18u
MI140 net129 d3 VDD VDD p w=0.42u l=0.18u
MI145 net124 net119 net64 VDD p w=0.75u l=0.18u
.ends
.subckt EDFCND2BWP7T D E CP CDN Q QN VDD VSS 
MI132 d0 INCPB net124 VSS n w=0.74u l=0.18u
MI133 net116 d3 VSS VSS n w=0.42u l=0.18u
MI49 net89 d1 VSS VSS n w=0.42u l=0.18u
MI48 net92 CDN net89 VSS n w=0.42u l=0.18u
MI47 d0 INCP net92 VSS n w=0.42u l=0.18u
MI18 d3 INCPB net98 VSS n w=0.42u l=0.18u
MI146 net124 E net088 VSS n w=0.57u l=0.18u
MI15 d1 INCP net98 VSS n w=0.91u l=0.18u
MI135 net088 D VSS VSS n w=0.57u l=0.18u
MI136 net124 net119 net116 VSS n w=0.42u l=0.18u
MI144-M_u4 XI144-net6 CDN VSS VSS n w=0.93u l=0.18u
MI144-M_u3 d2 net98 XI144-net6 VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI27_0-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI29_0-M_u2 QN d3 VSS VSS n w=1u l=0.18u
MI29_1-M_u2 QN d3 VSS VSS n w=1u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI14-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI137-M_u2 net119 E VSS VSS n w=0.5u l=0.18u
MI144-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI144-M_u1 d2 net98 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI27_0-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI29_0-M_u3 QN d3 VDD VDD p w=1.37u l=0.18u
MI29_1-M_u3 QN d3 VDD VDD p w=1.37u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI14-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI137-M_u3 net119 E VDD VDD p w=0.685u l=0.18u
MI44 net79 CDN VDD VDD p w=0.42u l=0.18u
MI43 net79 d1 VDD VDD p w=0.42u l=0.18u
MI45 d0 INCPB net79 VDD p w=0.42u l=0.18u
MI17 d3 INCP net98 VDD p w=0.42u l=0.18u
MI16 d1 INCPB net98 VDD p w=0.62u l=0.18u
MI138 d0 INCP net124 VDD p w=0.78u l=0.18u
MI139 net64 D VDD VDD p w=0.75u l=0.18u
MI141 net124 E net129 VDD p w=0.42u l=0.18u
MI140 net129 d3 VDD VDD p w=0.42u l=0.18u
MI145 net124 net119 net64 VDD p w=0.75u l=0.18u
.ends
.subckt EDFCNQD1BWP7T D E CP CDN Q VDD VSS 
MI132 d0 INCPB net124 VSS n w=0.74u l=0.18u
MI133 net116 net065 VSS VSS n w=0.42u l=0.18u
MI49 net89 d1 VSS VSS n w=0.42u l=0.18u
MI48 net92 CDN net89 VSS n w=0.42u l=0.18u
MI47 d0 INCP net92 VSS n w=0.42u l=0.18u
MI18 net065 INCPB net98 VSS n w=0.42u l=0.18u
MI146 net124 E net088 VSS n w=0.57u l=0.18u
MI15 d1 INCP net98 VSS n w=0.91u l=0.18u
MI135 net088 D VSS VSS n w=0.57u l=0.18u
MI136 net124 net119 net116 VSS n w=0.42u l=0.18u
MI144-M_u4 XI144-net6 CDN VSS VSS n w=0.93u l=0.18u
MI144-M_u3 d2 net98 XI144-net6 VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI27-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI14-M_u2 net065 d2 VSS VSS n w=0.42u l=0.18u
MI137-M_u2 net119 E VSS VSS n w=0.5u l=0.18u
MI144-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI144-M_u1 d2 net98 VDD VDD p w=1.03u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI27-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI14-M_u3 net065 d2 VDD VDD p w=0.42u l=0.18u
MI137-M_u3 net119 E VDD VDD p w=0.685u l=0.18u
MI44 net79 CDN VDD VDD p w=0.42u l=0.18u
MI43 net79 d1 VDD VDD p w=0.42u l=0.18u
MI45 d0 INCPB net79 VDD p w=0.42u l=0.18u
MI17 net065 INCP net98 VDD p w=0.42u l=0.18u
MI16 d1 INCPB net98 VDD p w=0.62u l=0.18u
MI138 d0 INCP net124 VDD p w=0.78u l=0.18u
MI139 net64 D VDD VDD p w=0.75u l=0.18u
MI141 net124 E net129 VDD p w=0.42u l=0.18u
MI140 net129 net065 VDD VDD p w=0.42u l=0.18u
MI145 net124 net119 net64 VDD p w=0.75u l=0.18u
.ends
.subckt EDFCNQD2BWP7T D E CP CDN Q VDD VSS 
MI132 d0 INCPB net124 VSS n w=0.74u l=0.18u
MI133 net116 net065 VSS VSS n w=0.42u l=0.18u
MI49 net89 d1 VSS VSS n w=0.42u l=0.18u
MI48 net92 CDN net89 VSS n w=0.42u l=0.18u
MI47 d0 INCP net92 VSS n w=0.42u l=0.18u
MI18 net065 INCPB net98 VSS n w=0.42u l=0.18u
MI146 net124 E net088 VSS n w=0.57u l=0.18u
MI15 d1 INCP net98 VSS n w=0.91u l=0.18u
MI135 net088 D VSS VSS n w=0.57u l=0.18u
MI136 net124 net119 net116 VSS n w=0.42u l=0.18u
MI144-M_u4 XI144-net6 CDN VSS VSS n w=0.93u l=0.18u
MI144-M_u3 d2 net98 XI144-net6 VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI27_0-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI14-M_u2 net065 d2 VSS VSS n w=0.42u l=0.18u
MI137-M_u2 net119 E VSS VSS n w=0.5u l=0.18u
MI144-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI144-M_u1 d2 net98 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI27_0-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI14-M_u3 net065 d2 VDD VDD p w=0.42u l=0.18u
MI137-M_u3 net119 E VDD VDD p w=0.685u l=0.18u
MI44 net79 CDN VDD VDD p w=0.42u l=0.18u
MI43 net79 d1 VDD VDD p w=0.42u l=0.18u
MI45 d0 INCPB net79 VDD p w=0.42u l=0.18u
MI17 net065 INCP net98 VDD p w=0.42u l=0.18u
MI16 d1 INCPB net98 VDD p w=0.62u l=0.18u
MI138 d0 INCP net124 VDD p w=0.78u l=0.18u
MI139 net64 D VDD VDD p w=0.75u l=0.18u
MI141 net124 E net129 VDD p w=0.42u l=0.18u
MI140 net129 net065 VDD VDD p w=0.42u l=0.18u
MI145 net124 net119 net64 VDD p w=0.75u l=0.18u
.ends
.subckt EDFD0BWP7T D E CP Q QN VDD VSS 
MI81 net92 net103 net98 VSS n w=0.42u l=0.18u
MI80 net081 D VSS VSS n w=0.57u l=0.18u
MI63 net117 INCP net85 VSS n w=0.42u l=0.18u
MI64 net85 net84 VSS VSS n w=0.42u l=0.18u
MI55 net99 INCPB net76 VSS n w=0.42u l=0.18u
MI65 net84 INCP net76 VSS n w=0.91u l=0.18u
MI78 net98 net99 VSS VSS n w=0.42u l=0.18u
MI77 net117 INCPB net92 VSS n w=0.91u l=0.18u
MI89 net92 E net081 VSS n w=0.57u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net99 VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q net58 VSS VSS n w=0.5u l=0.18u
MI73-M_u2 net58 net76 VSS VSS n w=0.5u l=0.18u
MI74-M_u2 net84 net117 VSS VSS n w=0.54u l=0.18u
MI75-M_u2 net99 net58 VSS VSS n w=0.42u l=0.18u
MI82-M_u2 net103 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net99 VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q net58 VDD VDD p w=0.685u l=0.18u
MI73-M_u3 net58 net76 VDD VDD p w=0.685u l=0.18u
MI74-M_u3 net84 net117 VDD VDD p w=0.785u l=0.18u
MI75-M_u3 net99 net58 VDD VDD p w=0.685u l=0.18u
MI82-M_u3 net103 E VDD VDD p w=0.685u l=0.18u
MI90 net92 net103 net59 VDD p w=0.75u l=0.18u
MI67 net84 INCPB net76 VDD p w=1.34u l=0.18u
MI68 net99 INCP net76 VDD p w=0.42u l=0.18u
MI69 net117 INCPB net69 VDD p w=0.42u l=0.18u
MI70 net69 net84 VDD VDD p w=0.42u l=0.18u
MI86 net92 E net110 VDD p w=0.42u l=0.18u
MI85 net110 net99 VDD VDD p w=0.42u l=0.18u
MI84 net59 D VDD VDD p w=0.75u l=0.18u
MI83 net117 INCP net92 VDD p w=0.62u l=0.18u
.ends
.subckt EDFD1BWP7T D E CP Q QN VDD VSS 
MI81 net92 net103 net98 VSS n w=0.42u l=0.18u
MI80 net081 D VSS VSS n w=0.57u l=0.18u
MI63 net117 INCP net85 VSS n w=0.42u l=0.18u
MI64 net85 net84 VSS VSS n w=0.42u l=0.18u
MI55 net99 INCPB net76 VSS n w=0.42u l=0.18u
MI65 net84 INCP net76 VSS n w=0.91u l=0.18u
MI78 net98 net99 VSS VSS n w=0.42u l=0.18u
MI77 net117 INCPB net92 VSS n w=0.91u l=0.18u
MI89 net92 E net081 VSS n w=0.57u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net99 VSS VSS n w=0.94u l=0.18u
MI27-M_u2 Q net58 VSS VSS n w=1u l=0.18u
MI73-M_u2 net58 net76 VSS VSS n w=1u l=0.18u
MI74-M_u2 net84 net117 VSS VSS n w=0.54u l=0.18u
MI75-M_u2 net99 net58 VSS VSS n w=0.42u l=0.18u
MI82-M_u2 net103 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net99 VDD VDD p w=1.37u l=0.18u
MI27-M_u3 Q net58 VDD VDD p w=1.37u l=0.18u
MI73-M_u3 net58 net76 VDD VDD p w=1.37u l=0.18u
MI74-M_u3 net84 net117 VDD VDD p w=0.785u l=0.18u
MI75-M_u3 net99 net58 VDD VDD p w=0.685u l=0.18u
MI82-M_u3 net103 E VDD VDD p w=0.685u l=0.18u
MI90 net92 net103 net59 VDD p w=0.75u l=0.18u
MI67 net84 INCPB net76 VDD p w=1.34u l=0.18u
MI68 net99 INCP net76 VDD p w=0.42u l=0.18u
MI69 net117 INCPB net69 VDD p w=0.42u l=0.18u
MI70 net69 net84 VDD VDD p w=0.42u l=0.18u
MI86 net92 E net110 VDD p w=0.42u l=0.18u
MI85 net110 net99 VDD VDD p w=0.42u l=0.18u
MI84 net59 D VDD VDD p w=0.75u l=0.18u
MI83 net117 INCP net92 VDD p w=0.62u l=0.18u
.ends
.subckt EDFD2BWP7T D E CP Q QN VDD VSS 
MI81 net92 net103 net98 VSS n w=0.42u l=0.18u
MI80 net081 D VSS VSS n w=0.57u l=0.18u
MI63 net117 INCP net85 VSS n w=0.42u l=0.18u
MI64 net85 net84 VSS VSS n w=0.42u l=0.18u
MI55 net99 INCPB net76 VSS n w=0.42u l=0.18u
MI65 net84 INCP net76 VSS n w=0.91u l=0.18u
MI78 net98 net99 VSS VSS n w=0.42u l=0.18u
MI77 net117 INCPB net92 VSS n w=0.91u l=0.18u
MI89 net92 E net081 VSS n w=0.57u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29_0-M_u2 QN net99 VSS VSS n w=1u l=0.18u
MI29_1-M_u2 QN net99 VSS VSS n w=1u l=0.18u
MI27_0-M_u2 Q net091 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q net091 VSS VSS n w=1u l=0.18u
MI73-M_u2 net091 net76 VSS VSS n w=1u l=0.18u
MI74-M_u2 net84 net117 VSS VSS n w=0.54u l=0.18u
MI75-M_u2 net99 net091 VSS VSS n w=1u l=0.18u
MI82-M_u2 net103 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29_0-M_u3 QN net99 VDD VDD p w=1.37u l=0.18u
MI29_1-M_u3 QN net99 VDD VDD p w=1.37u l=0.18u
MI27_0-M_u3 Q net091 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q net091 VDD VDD p w=1.37u l=0.18u
MI73-M_u3 net091 net76 VDD VDD p w=1.37u l=0.18u
MI74-M_u3 net84 net117 VDD VDD p w=0.785u l=0.18u
MI75-M_u3 net99 net091 VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net103 E VDD VDD p w=0.685u l=0.18u
MI90 net92 net103 net59 VDD p w=0.75u l=0.18u
MI67 net84 INCPB net76 VDD p w=1.34u l=0.18u
MI68 net99 INCP net76 VDD p w=0.42u l=0.18u
MI69 net117 INCPB net69 VDD p w=0.42u l=0.18u
MI70 net69 net84 VDD VDD p w=0.42u l=0.18u
MI86 net92 E net110 VDD p w=0.42u l=0.18u
MI85 net110 net99 VDD VDD p w=0.42u l=0.18u
MI84 net59 D VDD VDD p w=0.75u l=0.18u
MI83 net117 INCP net92 VDD p w=0.62u l=0.18u
.ends
.subckt EDFKCND0BWP7T D E CP CN Q QN VDD VSS 
MI47 net90 INCP net77 VSS n w=0.42u l=0.18u
MI63 net77 net82 VSS VSS n w=0.42u l=0.18u
MI64 net103 INCPB net86 VSS n w=0.42u l=0.18u
MI65 net82 INCP net86 VSS n w=0.42u l=0.18u
MI76 net98 CN VSS VSS n w=1u l=0.18u
MI74 net96 D net99 VSS n w=0.57u l=0.18u
MI73 net99 E net98 VSS n w=0.57u l=0.18u
MI72 net104 net103 net98 VSS n w=0.42u l=0.18u
MI75 net96 net107 net104 VSS n w=0.42u l=0.18u
MI87 net90 INCPB net96 VSS n w=0.91u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net103 VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q net56 VSS VSS n w=0.5u l=0.18u
MI68-M_u2 net56 net86 VSS VSS n w=0.5u l=0.18u
MI13-M_u2 net82 net90 VSS VSS n w=0.635u l=0.18u
MI14-M_u2 net103 net56 VSS VSS n w=0.5u l=0.18u
MI77-M_u2 net107 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net103 VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q net56 VDD VDD p w=0.685u l=0.18u
MI68-M_u3 net56 net86 VDD VDD p w=0.685u l=0.18u
MI13-M_u3 net82 net90 VDD VDD p w=0.97u l=0.18u
MI14-M_u3 net103 net56 VDD VDD p w=0.685u l=0.18u
MI77-M_u3 net107 E VDD VDD p w=0.685u l=0.18u
MI52 net82 INCPB net86 VDD p w=0.905u l=0.18u
MI66 net103 INCP net86 VDD p w=0.42u l=0.18u
MI45 net90 INCPB net70 VDD p w=0.42u l=0.18u
MI67 net70 net82 VDD VDD p w=0.42u l=0.18u
MI78 net96 D net120 VDD p w=0.72u l=0.18u
MI82 net96 CN VDD VDD p w=0.42u l=0.18u
MI81 net120 net107 VDD VDD p w=0.72u l=0.18u
MI80 net96 E net111 VDD p w=0.42u l=0.18u
MI79 net111 net103 VDD VDD p w=0.42u l=0.18u
MI86 net96 INCP net90 VDD p w=0.785u l=0.18u
.ends
.subckt EDFKCND1BWP7T D E CP CN Q QN VDD VSS 
MI47 net90 INCP net77 VSS n w=0.42u l=0.18u
MI63 net77 net82 VSS VSS n w=0.42u l=0.18u
MI64 net103 INCPB net86 VSS n w=0.42u l=0.18u
MI65 net82 INCP net86 VSS n w=0.635u l=0.18u
MI76 net98 CN VSS VSS n w=1u l=0.18u
MI74 net96 D net99 VSS n w=0.57u l=0.18u
MI73 net99 E net98 VSS n w=0.57u l=0.18u
MI72 net104 net103 net98 VSS n w=0.42u l=0.18u
MI75 net96 net107 net104 VSS n w=0.42u l=0.18u
MI87 net90 INCPB net96 VSS n w=0.91u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29-M_u2 QN net103 VSS VSS n w=1u l=0.18u
MI27-M_u2 Q net56 VSS VSS n w=1u l=0.18u
MI68-M_u2 net56 net86 VSS VSS n w=0.665u l=0.18u
MI13-M_u2 net82 net90 VSS VSS n w=0.635u l=0.18u
MI14-M_u2 net103 net56 VSS VSS n w=0.5u l=0.18u
MI77-M_u2 net107 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29-M_u3 QN net103 VDD VDD p w=1.235u l=0.18u
MI27-M_u3 Q net56 VDD VDD p w=1.37u l=0.18u
MI68-M_u3 net56 net86 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 net82 net90 VDD VDD p w=0.97u l=0.18u
MI14-M_u3 net103 net56 VDD VDD p w=0.685u l=0.18u
MI77-M_u3 net107 E VDD VDD p w=0.685u l=0.18u
MI52 net82 INCPB net86 VDD p w=1.215u l=0.18u
MI66 net103 INCP net86 VDD p w=0.42u l=0.18u
MI45 net90 INCPB net70 VDD p w=0.42u l=0.18u
MI67 net70 net82 VDD VDD p w=0.42u l=0.18u
MI78 net96 D net120 VDD p w=0.72u l=0.18u
MI82 net96 CN VDD VDD p w=0.42u l=0.18u
MI81 net120 net107 VDD VDD p w=0.72u l=0.18u
MI80 net96 E net111 VDD p w=0.42u l=0.18u
MI79 net111 net103 VDD VDD p w=0.42u l=0.18u
MI86 net96 INCP net90 VDD p w=0.65u l=0.18u
.ends
.subckt EDFKCND2BWP7T D E CP CN Q QN VDD VSS 
MI47 net90 INCP net77 VSS n w=0.42u l=0.18u
MI63 net77 net82 VSS VSS n w=0.42u l=0.18u
MI64 net103 INCPB net86 VSS n w=0.42u l=0.18u
MI65 net82 INCP net86 VSS n w=0.635u l=0.18u
MI76 net98 CN VSS VSS n w=1u l=0.18u
MI74 net96 D net99 VSS n w=0.57u l=0.18u
MI73 net99 E net98 VSS n w=0.57u l=0.18u
MI72 net104 net103 net98 VSS n w=0.42u l=0.18u
MI75 net96 net107 net104 VSS n w=0.42u l=0.18u
MI87 net90 INCPB net96 VSS n w=0.91u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI29_0-M_u2 QN net103 VSS VSS n w=1u l=0.18u
MI29_1-M_u2 QN net103 VSS VSS n w=1u l=0.18u
MI27_0-M_u2 Q net56 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q net56 VSS VSS n w=1u l=0.18u
MI68-M_u2 net56 net86 VSS VSS n w=0.665u l=0.18u
MI13-M_u2 net82 net90 VSS VSS n w=0.635u l=0.18u
MI14-M_u2 net103 net56 VSS VSS n w=0.5u l=0.18u
MI77-M_u2 net107 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI29_0-M_u3 QN net103 VDD VDD p w=1.37u l=0.18u
MI29_1-M_u3 QN net103 VDD VDD p w=1.37u l=0.18u
MI27_0-M_u3 Q net56 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q net56 VDD VDD p w=1.37u l=0.18u
MI68-M_u3 net56 net86 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 net82 net90 VDD VDD p w=0.97u l=0.18u
MI14-M_u3 net103 net56 VDD VDD p w=0.685u l=0.18u
MI77-M_u3 net107 E VDD VDD p w=0.685u l=0.18u
MI52 net82 INCPB net86 VDD p w=1.215u l=0.18u
MI66 net103 INCP net86 VDD p w=0.42u l=0.18u
MI45 net90 INCPB net70 VDD p w=0.42u l=0.18u
MI67 net70 net82 VDD VDD p w=0.42u l=0.18u
MI78 net96 D net120 VDD p w=0.72u l=0.18u
MI82 net96 CN VDD VDD p w=0.42u l=0.18u
MI81 net120 net107 VDD VDD p w=0.72u l=0.18u
MI80 net96 E net111 VDD p w=0.42u l=0.18u
MI79 net111 net103 VDD VDD p w=0.42u l=0.18u
MI86 net96 INCP net90 VDD p w=0.65u l=0.18u
.ends
.subckt EDFKCNQD1BWP7T D E CP CN Q VDD VSS 
MI47 net90 INCP net77 VSS n w=0.42u l=0.18u
MI63 net77 net82 VSS VSS n w=0.42u l=0.18u
MI64 net103 INCPB net86 VSS n w=0.42u l=0.18u
MI65 net82 INCP net86 VSS n w=0.635u l=0.18u
MI76 net98 CN VSS VSS n w=1u l=0.18u
MI74 net96 D net99 VSS n w=0.57u l=0.18u
MI73 net99 E net98 VSS n w=0.57u l=0.18u
MI72 net104 net103 net98 VSS n w=0.42u l=0.18u
MI75 net96 net107 net104 VSS n w=0.42u l=0.18u
MI87 net90 INCPB net96 VSS n w=0.91u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q net56 VSS VSS n w=1u l=0.18u
MI68-M_u2 net56 net86 VSS VSS n w=0.665u l=0.18u
MI13-M_u2 net82 net90 VSS VSS n w=0.97u l=0.18u
MI14-M_u2 net103 net56 VSS VSS n w=0.42u l=0.18u
MI77-M_u2 net107 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q net56 VDD VDD p w=1.37u l=0.18u
MI68-M_u3 net56 net86 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 net82 net90 VDD VDD p w=0.97u l=0.18u
MI14-M_u3 net103 net56 VDD VDD p w=0.42u l=0.18u
MI77-M_u3 net107 E VDD VDD p w=0.685u l=0.18u
MI52 net82 INCPB net86 VDD p w=1.215u l=0.18u
MI66 net103 INCP net86 VDD p w=0.42u l=0.18u
MI45 net90 INCPB net70 VDD p w=0.42u l=0.18u
MI67 net70 net82 VDD VDD p w=0.42u l=0.18u
MI78 net96 D net120 VDD p w=0.72u l=0.18u
MI82 net96 CN VDD VDD p w=0.42u l=0.18u
MI81 net120 net107 VDD VDD p w=0.72u l=0.18u
MI80 net96 E net111 VDD p w=0.42u l=0.18u
MI79 net111 net103 VDD VDD p w=0.42u l=0.18u
MI86 net96 INCP net90 VDD p w=0.65u l=0.18u
.ends
.subckt EDFKCNQD2BWP7T D E CP CN Q VDD VSS 
MI47 net90 INCP net77 VSS n w=0.42u l=0.18u
MI63 net77 net82 VSS VSS n w=0.42u l=0.18u
MI64 net103 INCPB net86 VSS n w=0.42u l=0.18u
MI65 net82 INCP net86 VSS n w=0.42u l=0.18u
MI76 net98 CN VSS VSS n w=1u l=0.18u
MI74 net96 D net99 VSS n w=0.57u l=0.18u
MI73 net99 E net98 VSS n w=0.57u l=0.18u
MI72 net104 net103 net98 VSS n w=0.42u l=0.18u
MI75 net96 net107 net104 VSS n w=0.42u l=0.18u
MI87 net90 INCPB net96 VSS n w=0.91u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27_0-M_u2 Q net56 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q net56 VSS VSS n w=1u l=0.18u
MI68-M_u2 net56 net86 VSS VSS n w=1u l=0.18u
MI13-M_u2 net82 net90 VSS VSS n w=0.97u l=0.18u
MI14-M_u2 net103 net56 VSS VSS n w=0.42u l=0.18u
MI77-M_u2 net107 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27_0-M_u3 Q net56 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q net56 VDD VDD p w=1.37u l=0.18u
MI68-M_u3 net56 net86 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 net82 net90 VDD VDD p w=0.97u l=0.18u
MI14-M_u3 net103 net56 VDD VDD p w=0.42u l=0.18u
MI77-M_u3 net107 E VDD VDD p w=0.685u l=0.18u
MI52 net82 INCPB net86 VDD p w=1.34u l=0.18u
MI66 net103 INCP net86 VDD p w=0.42u l=0.18u
MI45 net90 INCPB net70 VDD p w=0.42u l=0.18u
MI67 net70 net82 VDD VDD p w=0.42u l=0.18u
MI78 net96 D net120 VDD p w=0.72u l=0.18u
MI82 net96 CN VDD VDD p w=0.42u l=0.18u
MI81 net120 net107 VDD VDD p w=0.72u l=0.18u
MI80 net96 E net111 VDD p w=0.42u l=0.18u
MI79 net111 net103 VDD VDD p w=0.42u l=0.18u
MI86 net96 INCP net90 VDD p w=0.95u l=0.18u
.ends
.subckt EDFQD0BWP7T D E CP Q VDD VSS 
MI81 net92 net103 net98 VSS n w=0.42u l=0.18u
MI80 net081 D VSS VSS n w=0.57u l=0.18u
MI63 net117 INCP net85 VSS n w=0.42u l=0.18u
MI64 net85 net84 VSS VSS n w=0.42u l=0.18u
MI55 net99 INCPB net76 VSS n w=0.42u l=0.18u
MI65 net84 INCP net76 VSS n w=0.91u l=0.18u
MI78 net98 net99 VSS VSS n w=0.42u l=0.18u
MI77 net117 INCPB net92 VSS n w=0.91u l=0.18u
MI89 net92 E net081 VSS n w=0.57u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q net58 VSS VSS n w=0.5u l=0.18u
MI73-M_u2 net58 net76 VSS VSS n w=0.5u l=0.18u
MI74-M_u2 net84 net117 VSS VSS n w=0.54u l=0.18u
MI75-M_u2 net99 net58 VSS VSS n w=0.42u l=0.18u
MI82-M_u2 net103 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q net58 VDD VDD p w=0.685u l=0.18u
MI73-M_u3 net58 net76 VDD VDD p w=0.685u l=0.18u
MI74-M_u3 net84 net117 VDD VDD p w=0.785u l=0.18u
MI75-M_u3 net99 net58 VDD VDD p w=0.42u l=0.18u
MI82-M_u3 net103 E VDD VDD p w=0.685u l=0.18u
MI90 net92 net103 net59 VDD p w=0.75u l=0.18u
MI67 net84 INCPB net76 VDD p w=1.34u l=0.18u
MI68 net99 INCP net76 VDD p w=0.42u l=0.18u
MI69 net117 INCPB net69 VDD p w=0.42u l=0.18u
MI70 net69 net84 VDD VDD p w=0.42u l=0.18u
MI86 net92 E net110 VDD p w=0.42u l=0.18u
MI85 net110 net99 VDD VDD p w=0.42u l=0.18u
MI84 net59 D VDD VDD p w=0.75u l=0.18u
MI83 net117 INCP net92 VDD p w=0.62u l=0.18u
.ends
.subckt EDFQD1BWP7T D E CP Q VDD VSS 
MI81 net92 net103 net98 VSS n w=0.42u l=0.18u
MI80 net081 D VSS VSS n w=0.57u l=0.18u
MI63 net117 INCP net85 VSS n w=0.42u l=0.18u
MI64 net85 net84 VSS VSS n w=0.42u l=0.18u
MI55 net99 INCPB net76 VSS n w=0.42u l=0.18u
MI65 net84 INCP net76 VSS n w=0.91u l=0.18u
MI78 net98 net99 VSS VSS n w=0.42u l=0.18u
MI77 net117 INCPB net92 VSS n w=0.91u l=0.18u
MI89 net92 E net081 VSS n w=0.57u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27-M_u2 Q net58 VSS VSS n w=1u l=0.18u
MI73-M_u2 net58 net76 VSS VSS n w=1u l=0.18u
MI74-M_u2 net84 net117 VSS VSS n w=0.54u l=0.18u
MI75-M_u2 net99 net58 VSS VSS n w=0.42u l=0.18u
MI82-M_u2 net103 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27-M_u3 Q net58 VDD VDD p w=1.37u l=0.18u
MI73-M_u3 net58 net76 VDD VDD p w=1.37u l=0.18u
MI74-M_u3 net84 net117 VDD VDD p w=0.785u l=0.18u
MI75-M_u3 net99 net58 VDD VDD p w=0.42u l=0.18u
MI82-M_u3 net103 E VDD VDD p w=0.685u l=0.18u
MI90 net92 net103 net59 VDD p w=0.75u l=0.18u
MI67 net84 INCPB net76 VDD p w=1.34u l=0.18u
MI68 net99 INCP net76 VDD p w=0.42u l=0.18u
MI69 net117 INCPB net69 VDD p w=0.42u l=0.18u
MI70 net69 net84 VDD VDD p w=0.42u l=0.18u
MI86 net92 E net110 VDD p w=0.42u l=0.18u
MI85 net110 net99 VDD VDD p w=0.42u l=0.18u
MI84 net59 D VDD VDD p w=0.75u l=0.18u
MI83 net117 INCP net92 VDD p w=0.62u l=0.18u
.ends
.subckt EDFQD2BWP7T D E CP Q VDD VSS 
MI81 net92 net103 net98 VSS n w=0.42u l=0.18u
MI80 net081 D VSS VSS n w=0.57u l=0.18u
MI63 net117 INCP net85 VSS n w=0.42u l=0.18u
MI64 net85 net84 VSS VSS n w=0.42u l=0.18u
MI55 net99 INCPB net76 VSS n w=0.42u l=0.18u
MI65 net84 INCP net76 VSS n w=0.91u l=0.18u
MI78 net98 net99 VSS VSS n w=0.42u l=0.18u
MI77 net117 INCPB net92 VSS n w=0.91u l=0.18u
MI89 net92 E net081 VSS n w=0.57u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI27_0-M_u2 Q net087 VSS VSS n w=1u l=0.18u
MI27_1-M_u2 Q net087 VSS VSS n w=1u l=0.18u
MI73-M_u2 net087 net76 VSS VSS n w=1u l=0.18u
MI74-M_u2 net84 net117 VSS VSS n w=0.54u l=0.18u
MI75-M_u2 net99 net087 VSS VSS n w=0.42u l=0.18u
MI82-M_u2 net103 E VSS VSS n w=0.5u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI27_0-M_u3 Q net087 VDD VDD p w=1.37u l=0.18u
MI27_1-M_u3 Q net087 VDD VDD p w=1.37u l=0.18u
MI73-M_u3 net087 net76 VDD VDD p w=1.37u l=0.18u
MI74-M_u3 net84 net117 VDD VDD p w=0.785u l=0.18u
MI75-M_u3 net99 net087 VDD VDD p w=0.42u l=0.18u
MI82-M_u3 net103 E VDD VDD p w=0.685u l=0.18u
MI90 net92 net103 net59 VDD p w=0.75u l=0.18u
MI67 net84 INCPB net76 VDD p w=1.34u l=0.18u
MI68 net99 INCP net76 VDD p w=0.42u l=0.18u
MI69 net117 INCPB net69 VDD p w=0.42u l=0.18u
MI70 net69 net84 VDD VDD p w=0.42u l=0.18u
MI86 net92 E net110 VDD p w=0.42u l=0.18u
MI85 net110 net99 VDD VDD p w=0.42u l=0.18u
MI84 net59 D VDD VDD p w=0.75u l=0.18u
MI83 net117 INCP net92 VDD p w=0.62u l=0.18u
.ends
.subckt FA1D0BWP7T A B CI S CO VDD VSS 
MI19 net54 net32 net046 VSS n w=0.84u l=0.18u
MI36 net046 net67 VSS VSS n w=0.84u l=0.18u
MI38 net0108 net34 VSS VSS n w=0.88u l=0.18u
MI29 net32 net0112 net0108 VSS n w=0.88u l=0.18u
MU18-M_u2 S net54 VSS VSS n w=0.5u l=0.18u
MU1-M_u2 net34 A VSS VSS n w=0.88u l=0.18u
MU3-M_u2 net0112 B VSS VSS n w=0.425u l=0.18u
MU28-M_u2 CO net24 VSS VSS n w=0.5u l=0.18u
MU26-M_u2 net67 CI VSS VSS n w=0.84u l=0.18u
MU4-M_u2 net44 net32 VSS VSS n w=0.905u l=0.18u
MU17-M_u2 net67 net44 net54 VSS n w=0.465u l=0.18u
MI14-M_u2 net34 B net32 VSS n w=0.5u l=0.18u
MU27-M_u2 net0112 net44 net24 VSS n w=0.545u l=0.18u
MU25-M_u2 net67 net32 net24 VSS n w=0.7u l=0.18u
MI17 net055 net67 VDD VDD p w=1.16u l=0.18u
MI25 net54 net44 net055 VDD p w=1u l=0.18u
MI37 net32 B net0121 VDD p w=1.02u l=0.18u
MI32 net0121 net34 VDD VDD p w=1.18u l=0.18u
MU18-M_u3 S net54 VDD VDD p w=0.685u l=0.18u
MU1-M_u3 net34 A VDD VDD p w=1.18u l=0.18u
MU3-M_u3 net0112 B VDD VDD p w=0.655u l=0.18u
MU28-M_u3 CO net24 VDD VDD p w=0.685u l=0.18u
MU26-M_u3 net67 CI VDD VDD p w=1u l=0.18u
MU4-M_u3 net44 net32 VDD VDD p w=1.275u l=0.18u
MU17-M_u3 net67 net32 net54 VDD p w=0.88u l=0.18u
MI14-M_u3 net34 net0112 net32 VDD p w=0.725u l=0.18u
MU27-M_u3 net0112 net32 net24 VDD p w=1.01u l=0.18u
MU25-M_u3 net67 net44 net24 VDD p w=1.035u l=0.18u
.ends
.subckt FA1D1BWP7T A B CI S CO VDD VSS 
MI20 net54 net32 net049 VSS n w=0.84u l=0.18u
MI21 net049 net67 VSS VSS n w=0.84u l=0.18u
MI12_0-M_u2 net64 net34 VSS VSS n w=0.9225u l=0.18u
MI12_1-M_u2 net64 net34 VSS VSS n w=0.9225u l=0.18u
MU18-M_u2 S net54 VSS VSS n w=1u l=0.18u
MU1_0-M_u2 net34 A VSS VSS n w=1u l=0.18u
MU1_1-M_u2 net34 A VSS VSS n w=1u l=0.18u
MU3-M_u2 net36 B VSS VSS n w=0.425u l=0.18u
MU28-M_u2 CO net24 VSS VSS n w=1u l=0.18u
MU26_0-M_u2 net67 CI VSS VSS n w=0.84u l=0.18u
MU26_1-M_u2 net67 CI VSS VSS n w=0.84u l=0.18u
MU4-M_u2 net44 net32 VSS VSS n w=0.905u l=0.18u
MU17-M_u2 net67 net44 net54 VSS n w=0.465u l=0.18u
MI14-M_u2 net34 B net32 VSS n w=0.5u l=0.18u
MI13-M_u2 net64 net36 net32 VSS n w=0.88u l=0.18u
MU27-M_u2 net36 net44 net24 VSS n w=0.545u l=0.18u
MU25-M_u2 net67 net32 net24 VSS n w=0.7u l=0.18u
MI19 VDD net67 net045 VDD p w=1.16u l=0.18u
MI18 net045 net44 net54 VDD p w=1u l=0.18u
MI12_0-M_u3 net64 net34 VDD VDD p w=1.37u l=0.18u
MI12_1-M_u3 net64 net34 VDD VDD p w=1.37u l=0.18u
MU18-M_u3 S net54 VDD VDD p w=1.025u l=0.18u
MU1_0-M_u3 net34 A VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 net34 A VDD VDD p w=1.37u l=0.18u
MU3-M_u3 net36 B VDD VDD p w=0.655u l=0.18u
MU28-M_u3 CO net24 VDD VDD p w=1.37u l=0.18u
MU26_0-M_u3 net67 CI VDD VDD p w=1u l=0.18u
MU26_1-M_u3 net67 CI VDD VDD p w=1u l=0.18u
MU4-M_u3 net44 net32 VDD VDD p w=1.275u l=0.18u
MU17-M_u3 net67 net32 net54 VDD p w=0.88u l=0.18u
MI14-M_u3 net34 net36 net32 VDD p w=0.725u l=0.18u
MI13-M_u3 net64 B net32 VDD p w=1.04u l=0.18u
MU27-M_u3 net36 net32 net24 VDD p w=1.01u l=0.18u
MU25-M_u3 net67 net44 net24 VDD p w=1.035u l=0.18u
.ends
.subckt FA1D2BWP7T A B CI S CO VDD VSS 
MI20 net54 net32 net049 VSS n w=0.84u l=0.18u
MI21 net049 net67 VSS VSS n w=0.84u l=0.18u
MI12_0-M_u2 net64 net34 VSS VSS n w=0.9225u l=0.18u
MI12_1-M_u2 net64 net34 VSS VSS n w=0.9225u l=0.18u
MU18_0-M_u2 S net54 VSS VSS n w=0.5u l=0.18u
MU18_1-M_u2 S net54 VSS VSS n w=0.5u l=0.18u
MU1_0-M_u2 net34 A VSS VSS n w=1u l=0.18u
MU1_1-M_u2 net34 A VSS VSS n w=1u l=0.18u
MU3-M_u2 net36 B VSS VSS n w=0.425u l=0.18u
MU28_0-M_u2 CO net24 VSS VSS n w=1u l=0.18u
MU28_1-M_u2 CO net24 VSS VSS n w=1u l=0.18u
MU26_0-M_u2 net67 CI VSS VSS n w=0.84u l=0.18u
MU26_1-M_u2 net67 CI VSS VSS n w=0.84u l=0.18u
MU4-M_u2 net44 net32 VSS VSS n w=0.905u l=0.18u
MU17-M_u2 net67 net44 net54 VSS n w=0.465u l=0.18u
MI14-M_u2 net34 B net32 VSS n w=0.5u l=0.18u
MI13-M_u2 net64 net36 net32 VSS n w=0.88u l=0.18u
MU27-M_u2 net36 net44 net24 VSS n w=0.545u l=0.18u
MU25-M_u2 net67 net32 net24 VSS n w=0.7u l=0.18u
MI19 VDD net67 net045 VDD p w=1.16u l=0.18u
MI18 net045 net44 net54 VDD p w=1u l=0.18u
MI12_0-M_u3 net64 net34 VDD VDD p w=1.37u l=0.18u
MI12_1-M_u3 net64 net34 VDD VDD p w=1.37u l=0.18u
MU18_0-M_u3 S net54 VDD VDD p w=0.5125u l=0.18u
MU18_1-M_u3 S net54 VDD VDD p w=0.5125u l=0.18u
MU1_0-M_u3 net34 A VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 net34 A VDD VDD p w=1.37u l=0.18u
MU3-M_u3 net36 B VDD VDD p w=0.655u l=0.18u
MU28_0-M_u3 CO net24 VDD VDD p w=1.37u l=0.18u
MU28_1-M_u3 CO net24 VDD VDD p w=1.37u l=0.18u
MU26_0-M_u3 net67 CI VDD VDD p w=1u l=0.18u
MU26_1-M_u3 net67 CI VDD VDD p w=1u l=0.18u
MU4-M_u3 net44 net32 VDD VDD p w=1.275u l=0.18u
MU17-M_u3 net67 net32 net54 VDD p w=0.88u l=0.18u
MI14-M_u3 net34 net36 net32 VDD p w=0.725u l=0.18u
MI13-M_u3 net64 B net32 VDD p w=1.04u l=0.18u
MU27-M_u3 net36 net32 net24 VDD p w=1.01u l=0.18u
MU25-M_u3 net67 net44 net24 VDD p w=1.035u l=0.18u
.ends
.subckt GAN2D1BWP7T A1 A2 Z VDD VSS 
MI1 VSS net6 VSS VSS n w=1u l=0.18u
M_u3-M_u2 Z net6 VSS VSS n w=1u l=0.18u
M_u2-M_u4 X_u2-net6 A2 VSS VSS n w=1u l=0.18u
M_u2-M_u3 net6 A1 X_u2-net6 VSS n w=1u l=0.18u
MI2 VDD net6 VDD VDD p w=1.37u l=0.18u
M_u3-M_u3 Z net6 VDD VDD p w=1.37u l=0.18u
M_u2-M_u2 net6 A2 VDD VDD p w=1.37u l=0.18u
M_u2-M_u1 net6 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GAN2D2BWP7T A1 A2 Z VDD VSS 
M_u3-M_u2 Z net10 VSS VSS n w=2u l=0.18u
M_u2-M_u4 X_u2-net6 A2 VSS VSS n w=1u l=0.18u
M_u2-M_u3 net10 A1 X_u2-net6 VSS n w=1u l=0.18u
M_u3-M_u3 Z net10 VDD VDD p w=2.74u l=0.18u
M_u2-M_u2 net10 A2 VDD VDD p w=1.37u l=0.18u
M_u2-M_u1 net10 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GAOI21D1BWP7T A1 A2 B ZN VDD VSS 
MI2 ZN A1 net27 VSS n w=1u l=0.18u
MI3 net27 A2 VSS VSS n w=1u l=0.18u
MI5 ZN B VSS VSS n w=1u l=0.18u
M_u7 ZN B VSS VSS n w=1u l=0.18u
MI4 net13 B VDD VDD p w=1.37u l=0.18u
M_u4 net13 A2 ZN VDD p w=1.37u l=0.18u
M_u2 net13 B VDD VDD p w=1.37u l=0.18u
M_u3 net13 A1 ZN VDD p w=1.37u l=0.18u
.ends
.subckt GAOI21D2BWP7T A1 A2 B ZN VDD VSS 
MI2 ZN A1 p0 VSS n w=1u l=0.18u
MI12 p0 A2 VSS VSS n w=1u l=0.18u
MI13 ZN A1 net23 VSS n w=1u l=0.18u
MI14 net23 A2 VSS VSS n w=1u l=0.18u
MI11_0 ZN B VSS VSS n w=1u l=0.18u
MI11_1 ZN B VSS VSS n w=1u l=0.18u
MI8 ZN A2 net74 VDD p w=2.74u l=0.18u
M_u2 net74 B VDD VDD p w=2.74u l=0.18u
MI9 ZN A1 net74 VDD p w=2.74u l=0.18u
.ends
.subckt GAOI22D1BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI16 ZN B1 net29 VSS n w=1u l=0.18u
MI15 net29 B2 VSS VSS n w=1u l=0.18u
MI20 net23 A2 VSS VSS n w=1u l=0.18u
MI19 ZN A1 net23 VSS n w=1u l=0.18u
MI13 net20 A1 ZN VDD p w=1.37u l=0.18u
M_u4 VDD B1 net20 VDD p w=1.37u l=0.18u
MI12 net20 A2 ZN VDD p w=1.37u l=0.18u
MI11 VDD B2 net20 VDD p w=1.37u l=0.18u
.ends
.subckt GBUFFD1BWP7T I Z VDD VSS 
MI1-M_u2 Z net6 VSS VSS n w=1u l=0.18u
MI2-M_u2 net6 I VSS VSS n w=1u l=0.18u
MI1-M_u3 Z net6 VDD VDD p w=1.37u l=0.18u
MI2-M_u3 net6 I VDD VDD p w=1.37u l=0.18u
.ends
.subckt GBUFFD2BWP7T I Z VDD VSS 
MI0-M_u2 net8 I VSS VSS n w=1u l=0.18u
M_u2-M_u2 net8 I VSS VSS n w=1u l=0.18u
M_u3_0-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z net8 VSS VSS n w=1u l=0.18u
MI0-M_u3 net8 I VDD VDD p w=1.37u l=0.18u
M_u2-M_u3 net8 I VDD VDD p w=1.37u l=0.18u
M_u3_0-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GBUFFD3BWP7T I Z VDD VSS 
M_u3_0-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u3_2-M_u2 Z net8 VSS VSS n w=1u l=0.18u
M_u2-M_u2 net8 I VSS VSS n w=1u l=0.18u
M_u3_0-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u3_2-M_u3 Z net8 VDD VDD p w=1.37u l=0.18u
M_u2-M_u3 net8 I VDD VDD p w=1.37u l=0.18u
.ends
.subckt GBUFFD8BWP7T I Z VDD VSS 
MI1-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u2_0-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u2_1-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u2_2-M_u2 n0 I VSS VSS n w=1u l=0.18u
M_u7_0-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_1-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_2-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_3-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_4-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_5-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_6-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_7-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MI1-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u2_0-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u2_1-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u2_2-M_u3 n0 I VDD VDD p w=1.37u l=0.18u
M_u7_0-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_1-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_2-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_3-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_4-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_5-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_6-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_7-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GDCAP10BWP7T VDD VSS 
MI4 VSS net016 VSS VSS n w=10u l=0.18u
M_u2 net016 net8 VSS VSS n w=10u l=0.18u
MI3 VDD net8 VDD VDD p w=13.7u l=0.18u
M_u1 net8 net016 VDD VDD p w=13.7u l=0.18u
.ends
.subckt GDCAP2BWP7T VDD VSS 
MI5 net13 net16 VSS VSS n w=2u l=0.18u
MI4 VSS net13 VSS VSS n w=2u l=0.18u
MI1 net16 net13 VDD VDD p w=2.74u l=0.18u
MI3 VDD net16 VDD VDD p w=2.74u l=0.18u
.ends
.subckt GDCAP3BWP7T VDD VSS 
MI5 net7 net10 VSS VSS n w=3u l=0.18u
MI4 VSS net7 VSS VSS n w=3u l=0.18u
MI3 VDD net10 VDD VDD p w=4.11u l=0.18u
MI1 net10 net7 VDD VDD p w=4.11u l=0.18u
.ends
.subckt GDCAP4BWP7T VDD VSS 
MI5 net7 net10 VSS VSS n w=4u l=0.18u
MI4 VSS net7 VSS VSS n w=4u l=0.18u
MI3 VDD net10 VDD VDD p w=5.48u l=0.18u
MI1 net10 net7 VDD VDD p w=5.48u l=0.18u
.ends
.subckt GDCAPBWP7T VDD VSS 
MI4 VSS net16 VSS VSS n w=1u l=0.18u
MI5 net16 net13 VSS VSS n w=1u l=0.18u
MI3 VDD net13 VDD VDD p w=1.37u l=0.18u
MI1 net13 net16 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GDFCNQD1BWP7T D CP CDN Q VDD VSS 
MI4 net52 D VSS VSS n w=1u l=0.18u
MI15 d1 CP d2 VSS n w=1u l=0.18u
MI5 d0 net075 net52 VSS n w=1u l=0.18u
MI18 net101 net072 d2 VSS n w=1u l=0.18u
MI47 d0 CP net59 VSS n w=1u l=0.18u
MI48 net59 d1 net62 VSS n w=1u l=0.18u
MI49 net62 CDN VSS VSS n w=1u l=0.18u
MI21-M_u4 XI21-net6 d2 VSS VSS n w=1u l=0.18u
MI21-M_u3 d3 CDN XI21-net6 VSS n w=1u l=0.18u
MI22-M_u2 net075 CP VSS VSS n w=1u l=0.18u
MI31-M_u2 net072 CP VSS VSS n w=1u l=0.18u
MI27-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI13-M_u2 d1 d0 VSS VSS n w=1u l=0.18u
MI14-M_u2 net101 d3 VSS VSS n w=1u l=0.18u
MI21-M_u2 d3 d2 VDD VDD p w=1.37u l=0.18u
MI21-M_u1 d3 CDN VDD VDD p w=1.37u l=0.18u
MI22-M_u3 net075 CP VDD VDD p w=1.37u l=0.18u
MI31-M_u3 net072 CP VDD VDD p w=1.37u l=0.18u
MI27-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI13-M_u3 d1 d0 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net101 d3 VDD VDD p w=1.37u l=0.18u
MI6 d0 CP net85 VDD p w=1.37u l=0.18u
MI7 net85 D VDD VDD p w=1.37u l=0.18u
MI16 d1 net072 d2 VDD p w=1.37u l=0.18u
MI17 net101 CP d2 VDD p w=1.37u l=0.18u
MI45 d0 net075 net98 VDD p w=1.37u l=0.18u
MI43 net98 d1 VDD VDD p w=1.37u l=0.18u
MI44 net98 CDN VDD VDD p w=1.37u l=0.18u
.ends
.subckt GDFQD1BWP7T D CP Q VDD VSS 
MI4 net66 D VSS VSS n w=1u l=0.18u
MI57 SLI INCPB net043 VSS n w=1u l=0.18u
MI58 net043 SLO VSS VSS n w=1u l=0.18u
MI5 MLI INCPB net66 VSS n w=1u l=0.18u
MI47 MLI INCP net50 VSS n w=1u l=0.18u
MI48 net50 MLO VSS VSS n w=1u l=0.18u
MI50 MLO INCP SLI VSS n w=1u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=1u l=0.18u
MI31-M_u2 INCPB CP VSS VSS n w=1u l=0.18u
MI27-M_u2 Q SLO VSS VSS n w=1u l=0.18u
MI53-M_u2 SLO SLI VSS VSS n w=1u l=0.18u
MI13-M_u2 MLO MLI VSS VSS n w=1u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=1.37u l=0.18u
MI31-M_u3 INCPB CP VDD VDD p w=1.37u l=0.18u
MI27-M_u3 Q SLO VDD VDD p w=1.37u l=0.18u
MI53-M_u3 SLO SLI VDD VDD p w=1.37u l=0.18u
MI13-M_u3 MLO MLI VDD VDD p w=1.37u l=0.18u
MI6 MLI INCP net66 VDD p w=1.37u l=0.18u
MI7 net66 D VDD VDD p w=1.37u l=0.18u
MI61 net071 SLO VDD VDD p w=1.37u l=0.18u
MI60 SLI INCP net071 VDD p w=1.37u l=0.18u
MI52 MLO INCPB SLI VDD p w=1.37u l=0.18u
MI45 MLI INCPB net84 VDD p w=1.37u l=0.18u
MI43 net84 MLO VDD VDD p w=1.37u l=0.18u
.ends
.subckt GFILL10BWP7T VDD VSS 
MI22 net0154 net032 net0154 vss n w=1u l=0.18u
MI23 net032 net018 net0154 vss n w=1u l=0.18u
MI24 net0148 net032 net0148 vss n w=1u l=0.18u
MI25 net032 net018 net0148 vss n w=1u l=0.18u
MI26 net0142 net032 net0142 vss n w=1u l=0.18u
MI27 net032 net018 net0142 vss n w=1u l=0.18u
MI28 net0136 net032 net0136 vss n w=1u l=0.18u
MI29 net032 net018 net0136 vss n w=1u l=0.18u
MI37 net0121 net032 net0121 vss n w=1u l=0.18u
MI36 net032 net018 net0121 vss n w=1u l=0.18u
MI35 net0127 net032 net0127 vss n w=1u l=0.18u
MI34 net032 net018 net0127 vss n w=1u l=0.18u
MI10 net064 net032 net064 vss n w=1u l=0.18u
MI11 net032 net018 net064 vss n w=1u l=0.18u
MI12 net058 net032 net058 vss n w=1u l=0.18u
MI13 net032 net018 net058 vss n w=1u l=0.18u
MI4 net030 net032 net030 vss n w=1u l=0.18u
MI5 net032 net018 net030 vss n w=1u l=0.18u
M_u2 net11 net032 net11 vss n w=1u l=0.18u
MI1 net032 net018 net11 vss n w=1u l=0.18u
MI14 net018 net032 net096 vdd p w=1.37u l=0.18u
MI15 net096 net018 net096 vdd p w=1.37u l=0.18u
MI16 net018 net032 net090 vdd p w=1.37u l=0.18u
MI17 net090 net018 net090 vdd p w=1.37u l=0.18u
MI18 net018 net032 net084 vdd p w=1.37u l=0.18u
MI19 net084 net018 net084 vdd p w=1.37u l=0.18u
MI20 net018 net032 net078 vdd p w=1.37u l=0.18u
MI21 net078 net018 net078 vdd p w=1.37u l=0.18u
MI33 net018 net032 net063 vdd p w=1.37u l=0.18u
MI32 net063 net018 net063 vdd p w=1.37u l=0.18u
MI30 net069 net018 net069 vdd p w=1.37u l=0.18u
MI31 net018 net032 net069 vdd p w=1.37u l=0.18u
MI6 net018 net032 net042 vdd p w=1.37u l=0.18u
MI7 net042 net018 net042 vdd p w=1.37u l=0.18u
MI8 net018 net032 net036 vdd p w=1.37u l=0.18u
MI9 net036 net018 net036 vdd p w=1.37u l=0.18u
MI2 net018 net032 net020 vdd p w=1.37u l=0.18u
MI3 net020 net018 net020 vdd p w=1.37u l=0.18u
M_u3 net018 net032 net6 vdd p w=1.37u l=0.18u
MI0 net6 net018 net6 vdd p w=1.37u l=0.18u
.ends
.subckt GFILL2BWP7T VDD VSS 
MI4 net030 net032 net030 vss n w=1u l=0.18u
MI5 net032 net018 net030 vss n w=1u l=0.18u
M_u2 net11 net032 net11 vss n w=1u l=0.18u
MI1 net032 net018 net11 vss n w=1u l=0.18u
MI2 net018 net032 net020 vdd p w=1.37u l=0.18u
MI3 net020 net018 net020 vdd p w=1.37u l=0.18u
M_u3 net018 net032 net6 vdd p w=1.37u l=0.18u
MI0 net6 net018 net6 vdd p w=1.37u l=0.18u
.ends
.subckt GFILL3BWP7T VDD VSS 
MI8 net074 net076 net074 vss n w=1u l=0.18u
MI9 net076 net056 net074 vss n w=1u l=0.18u
MI4 net030 net076 net030 vss n w=1u l=0.18u
MI5 net076 net056 net030 vss n w=1u l=0.18u
M_u2 net11 net076 net11 vss n w=1u l=0.18u
MI1 net076 net056 net11 vss n w=1u l=0.18u
MI6 net056 net076 net058 vdd p w=1.37u l=0.18u
MI7 net058 net056 net058 vdd p w=1.37u l=0.18u
MI2 net056 net076 net020 vdd p w=1.37u l=0.18u
MI3 net020 net056 net020 vdd p w=1.37u l=0.18u
M_u3 net056 net076 net6 vdd p w=1.37u l=0.18u
MI0 net6 net056 net6 vdd p w=1.37u l=0.18u
.ends
.subckt GFILL4BWP7T VDD VSS 
MI10 net064 net032 net064 vss n w=1u l=0.18u
MI11 net032 net018 net064 vss n w=1u l=0.18u
MI12 net058 net032 net058 vss n w=1u l=0.18u
MI13 net032 net018 net058 vss n w=1u l=0.18u
MI4 net030 net032 net030 vss n w=1u l=0.18u
MI5 net032 net018 net030 vss n w=1u l=0.18u
M_u2 net11 net032 net11 vss n w=1u l=0.18u
MI1 net032 net018 net11 vss n w=1u l=0.18u
MI6 net018 net032 net042 vdd p w=1.37u l=0.18u
MI7 net042 net018 net042 vdd p w=1.37u l=0.18u
MI8 net018 net032 net036 vdd p w=1.37u l=0.18u
MI9 net036 net018 net036 vdd p w=1.37u l=0.18u
MI2 net018 net032 net020 vdd p w=1.37u l=0.18u
MI3 net020 net018 net020 vdd p w=1.37u l=0.18u
M_u3 net018 net032 net6 vdd p w=1.37u l=0.18u
MI0 net6 net018 net6 vdd p w=1.37u l=0.18u
.ends
.subckt GFILLBWP7T VDD VSS 
M_u2 net11 net12 net11 vss n w=1u l=0.18u
MI1 net12 net4 net11 vss n w=1u l=0.18u
M_u3 net4 net12 net6 vdd p w=1.37u l=0.18u
MI0 net6 net4 net6 vdd p w=1.37u l=0.18u
.ends
.subckt GINVD1BWP7T I ZN VDD VSS 
MI1 VSS I VSS VSS n w=1u l=0.18u
MU1-M_u2 ZN I VSS VSS n w=1u l=0.18u
MI2 VDD I VDD VDD p w=1.37u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt GINVD2BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=2u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=2.74u l=0.18u
.ends
.subckt GINVD3BWP7T I ZN VDD VSS 
MI1 VSS I VSS VSS n w=1u l=0.18u
MU1-M_u2 ZN I VSS VSS n w=3u l=0.18u
MI2 VDD I VDD VDD p w=1.37u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=4.11u l=0.18u
.ends
.subckt GINVD8BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=8u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=10.96u l=0.18u
.ends
.subckt GMUX2D1BWP7T I0 I1 S Z VDD VSS 
MI15-M_u2 net6 S VSS VSS n w=1u l=0.18u
MU29-M_u2 Z net28 VSS VSS n w=1u l=0.18u
M_u2 net026 I0 VSS VSS n w=1u l=0.18u
MI17 net28 net6 net026 VSS n w=1u l=0.18u
MI23 net056 I1 VSS VSS n w=1u l=0.18u
MI24 net28 S net056 VSS n w=1u l=0.18u
MI15-M_u3 net6 S VDD VDD p w=1.37u l=0.18u
MU29-M_u3 Z net28 VDD VDD p w=1.37u l=0.18u
MI21 net28 net6 net045 VDD p w=1.37u l=0.18u
M_u1 net021 I0 VDD VDD p w=1.37u l=0.18u
MI16 net28 S net021 VDD p w=1.37u l=0.18u
MI22 net045 I1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GMUX2D2BWP7T I0 I1 S Z VDD VSS 
MI15-M_u2 net043 S VSS VSS n w=1u l=0.18u
MU29_0-M_u2 Z net026 VSS VSS n w=1u l=0.18u
MU29_1-M_u2 Z net026 VSS VSS n w=1u l=0.18u
MI26 net023 I1 VSS VSS n w=1u l=0.18u
MI23 net023 I1 VSS VSS n w=1u l=0.18u
MI24 net026 S net023 VSS n w=1u l=0.18u
MI17 net026 net043 net029 VSS n w=1u l=0.18u
M_u2 net029 I0 VSS VSS n w=1u l=0.18u
MI15-M_u3 net043 S VDD VDD p w=1.37u l=0.18u
MU29_0-M_u3 Z net026 VDD VDD p w=1.37u l=0.18u
MU29_1-M_u3 Z net026 VDD VDD p w=1.37u l=0.18u
MI25 net042 I1 VDD VDD p w=1.37u l=0.18u
MI21 net026 net043 net042 VDD p w=1.37u l=0.18u
M_u1 net036 I0 VDD VDD p w=1.37u l=0.18u
MI22 net042 I1 VDD VDD p w=1.37u l=0.18u
MI16 net026 S net036 VDD p w=1.37u l=0.18u
.ends
.subckt GMUX2ND1BWP7T I0 I1 S ZN VDD VSS 
MI15-M_u2 net045 S VSS VSS n w=1u l=0.18u
MI16-M_u2 net48 net28 VSS VSS n w=1u l=0.18u
MU29-M_u2 ZN net48 VSS VSS n w=1u l=0.18u
MI27 net025 I1 VSS VSS n w=1u l=0.18u
MI25 net28 S net025 VSS n w=1u l=0.18u
M_u2 net031 I0 VSS VSS n w=1u l=0.18u
MI24 net025 I1 VSS VSS n w=1u l=0.18u
MI23 net28 net045 net031 VSS n w=1u l=0.18u
MI15-M_u3 net045 S VDD VDD p w=1.37u l=0.18u
MI16-M_u3 net48 net28 VDD VDD p w=1.37u l=0.18u
MU29-M_u3 ZN net48 VDD VDD p w=1.37u l=0.18u
MI26 net044 I1 VDD VDD p w=1.37u l=0.18u
M_u1 net038 I0 VDD VDD p w=1.37u l=0.18u
MI17 net28 S net038 VDD p w=1.37u l=0.18u
MI22 net044 I1 VDD VDD p w=1.37u l=0.18u
MI21 net28 net045 net044 VDD p w=1.37u l=0.18u
.ends
.subckt GMUX2ND2BWP7T I0 I1 S ZN VDD VSS 
MI15-M_u2 net045 S VSS VSS n w=1u l=0.18u
MI16-M_u2 net27 net28 VSS VSS n w=1u l=0.18u
MU29_0-M_u2 ZN net27 VSS VSS n w=1u l=0.18u
MU29_1-M_u2 ZN net27 VSS VSS n w=1u l=0.18u
MI25 net28 S net025 VSS n w=1u l=0.18u
M_u2 net031 I0 VSS VSS n w=1u l=0.18u
MI24 net025 I1 VSS VSS n w=1u l=0.18u
MI17 net28 net045 net031 VSS n w=1u l=0.18u
MI15-M_u3 net045 S VDD VDD p w=1.37u l=0.18u
MI16-M_u3 net27 net28 VDD VDD p w=1.37u l=0.18u
MU29_0-M_u3 ZN net27 VDD VDD p w=1.37u l=0.18u
MU29_1-M_u3 ZN net27 VDD VDD p w=1.37u l=0.18u
M_u1 net038 I0 VDD VDD p w=1.37u l=0.18u
MI22 net28 S net038 VDD p w=1.37u l=0.18u
MI23 net044 I1 VDD VDD p w=1.37u l=0.18u
MI21 net28 net045 net044 VDD p w=1.37u l=0.18u
.ends
.subckt GND2D1BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 XI1-net6 A1 VSS VSS n w=1u l=0.18u
MI1-M_u3 ZN A2 XI1-net6 VSS n w=1u l=0.18u
MI1-M_u2 ZN A1 VDD VDD p w=1.37u l=0.18u
MI1-M_u1 ZN A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GND2D2BWP7T A1 A2 ZN VDD VSS 
MU3_0-M_u4 XU3_0-net6 A2 VSS VSS n w=1u l=0.18u
MU3_0-M_u3 ZN A1 XU3_0-net6 VSS n w=1u l=0.18u
MU3_1-M_u4 XU3_1-net6 A2 VSS VSS n w=1u l=0.18u
MU3_1-M_u3 ZN A1 XU3_1-net6 VSS n w=1u l=0.18u
MU3_0-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
MU3_0-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
MU3_1-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
MU3_1-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GND2D3BWP7T A1 A2 ZN VDD VSS 
MI2_0 net19 A2 VSS VSS n w=1u l=0.18u
MI2_1 net19 A2 VSS VSS n w=1u l=0.18u
MI2_2 net19 A2 VSS VSS n w=1u l=0.18u
MI3_0 ZN A1 net19 VSS n w=1u l=0.18u
MI3_1 ZN A1 net19 VSS n w=1u l=0.18u
MI3_2 ZN A1 net19 VSS n w=1u l=0.18u
MI4_0 ZN A2 VDD VDD p w=1.37u l=0.18u
MI4_1 ZN A2 VDD VDD p w=1.37u l=0.18u
MI4_2 ZN A2 VDD VDD p w=1.37u l=0.18u
MI5_0 ZN A1 VDD VDD p w=1.37u l=0.18u
MI5_1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI5_2 ZN A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GND3D1BWP7T A1 A2 A3 ZN VDD VSS 
MI1-M_u4 ZN A3 XI1-net10 VSS n w=1u l=0.18u
MI1-M_u5 XI1-net10 A2 XI1-net13 VSS n w=1u l=0.18u
MI1-M_u6_0 XI1-net13 A1 VSS VSS n w=1u l=0.18u
MI1-M_u6_1 XI1-net13 A1 VSS VSS n w=1u l=0.18u
MI1-M_u3_0 ZN A1 VDD VDD p w=1.37u l=0.18u
MI1-M_u3_1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI1-M_u1 ZN A3 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GND3D2BWP7T A1 A2 A3 ZN VDD VSS 
MI0_0-M_u4 ZN A1 XI0_0-net10 VSS n w=1u l=0.18u
MI0_0-M_u5 XI0_0-net10 A2 XI0_0-net13 VSS n w=1u l=0.18u
MI0_0-M_u6 XI0_0-net13 A3 VSS VSS n w=1u l=0.18u
MI0_1-M_u4 ZN A1 XI0_1-net10 VSS n w=1u l=0.18u
MI0_1-M_u5 XI0_1-net10 A2 XI0_1-net13 VSS n w=1u l=0.18u
MI0_1-M_u6 XI0_1-net13 A3 VSS VSS n w=1u l=0.18u
MI0_0-M_u3 ZN A3 VDD VDD p w=1.37u l=0.18u
MI0_0-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI0_0-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
MI0_1-M_u3 ZN A3 VDD VDD p w=1.37u l=0.18u
MI0_1-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI0_1-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GNR2D1BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A2 VSS VSS n w=1u l=0.18u
MI1-M_u3 ZN A1 VSS VSS n w=1u l=0.18u
MI1-M_u1 XI1-net8 A1 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 ZN A2 XI1-net8 VDD p w=1.37u l=0.18u
.ends
.subckt GNR2D2BWP7T A1 A2 ZN VDD VSS 
MI2-M_u4 ZN A2 VSS VSS n w=1u l=0.18u
MI2-M_u3 ZN A1 VSS VSS n w=1u l=0.18u
MI1-M_u4 ZN A2 VSS VSS n w=1u l=0.18u
MI1-M_u3 ZN A1 VSS VSS n w=1u l=0.18u
MI2-M_u1 XI2-net8 A1 VDD VDD p w=1.37u l=0.18u
MI2-M_u2 ZN A2 XI2-net8 VDD p w=1.37u l=0.18u
MI1-M_u1 XI1-net8 A1 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 ZN A2 XI1-net8 VDD p w=1.37u l=0.18u
.ends
.subckt GNR3D1BWP7T A1 A2 A3 ZN VDD VSS 
M_u4 ZN A3 VSS VSS n w=1u l=0.18u
MI5 ZN A3 VSS VSS n w=1u l=0.18u
MI2 ZN A2 VSS VSS n w=1u l=0.18u
MI3 ZN A1 VSS VSS n w=1u l=0.18u
MI4 net025 A3 VDD VDD p w=1.37u l=0.18u
M_u1 net025 A3 VDD VDD p w=1.37u l=0.18u
MI0 net028 A2 net025 VDD p w=1.37u l=0.18u
MI1 ZN A1 net028 VDD p w=1.37u l=0.18u
.ends
.subckt GNR3D2BWP7T A1 A2 A3 ZN VDD VSS 
M_u4_0 ZN A3 VSS VSS n w=1u l=0.18u
M_u4_1 ZN A3 VSS VSS n w=1u l=0.18u
MI7_0 ZN A1 VSS VSS n w=1u l=0.18u
MI7_1 ZN A1 VSS VSS n w=1u l=0.18u
MI6_0 ZN A2 VSS VSS n w=1u l=0.18u
MI6_1 ZN A2 VSS VSS n w=1u l=0.18u
M_u1 net70 A3 VDD VDD p w=2.74u l=0.18u
MI20 net67 A2 net70 VDD p w=2.74u l=0.18u
MI21 ZN A1 net67 VDD p w=2.74u l=0.18u
.ends
.subckt GOAI21D1BWP7T A1 A2 B ZN VDD VSS 
MI0 net15 B VSS VSS n w=1u l=0.18u
M_u2 ZN A1 net15 VSS n w=1u l=0.18u
M_u3 ZN A2 net15 VSS n w=1u l=0.18u
M_u4 net15 B VSS VSS n w=1u l=0.18u
MI1 ZN B VDD VDD p w=1.37u l=0.18u
M_u9 ZN B VDD VDD p w=1.37u l=0.18u
MI16-MI12 ZN A1 XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GOAI21D2BWP7T A1 A2 B ZN VDD VSS 
M_u2 ZN A1 net15 VSS n w=2u l=0.18u
M_u3 ZN A2 net15 VSS n w=2u l=0.18u
M_u4 net15 B VSS VSS n w=2u l=0.18u
M_u9 ZN B VDD VDD p w=2.74u l=0.18u
MI16_0-MI12 ZN A1 XI16_0-net11 VDD p w=1.37u l=0.18u
MI16_0-MI13 XI16_0-net11 A2 VDD VDD p w=1.37u l=0.18u
MI16_1-MI12 ZN A1 XI16_1-net11 VDD p w=1.37u l=0.18u
MI16_1-MI13 XI16_1-net11 A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GOR2D1BWP7T A1 A2 Z VDD VSS 
MI1 VSS net7 VSS VSS n w=1u l=0.18u
MU1-M_u2 Z net7 VSS VSS n w=1u l=0.18u
M_u7-M_u4 net7 A1 VSS VSS n w=1u l=0.18u
M_u7-M_u3 net7 A2 VSS VSS n w=1u l=0.18u
MI2 VDD net7 VDD VDD p w=1.37u l=0.18u
MU1-M_u3 Z net7 VDD VDD p w=1.37u l=0.18u
M_u7-M_u1 X_u7-net8 A2 VDD VDD p w=1.37u l=0.18u
M_u7-M_u2 net7 A1 X_u7-net8 VDD p w=1.37u l=0.18u
.ends
.subckt GOR2D2BWP7T A1 A2 Z VDD VSS 
MU1_0-M_u2 Z net9 VSS VSS n w=1u l=0.18u
MU1_1-M_u2 Z net9 VSS VSS n w=1u l=0.18u
M_u7-M_u4 net9 A1 VSS VSS n w=1u l=0.18u
M_u7-M_u3 net9 A2 VSS VSS n w=1u l=0.18u
MU1_0-M_u3 Z net9 VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 Z net9 VDD VDD p w=1.37u l=0.18u
M_u7-M_u1 X_u7-net8 A2 VDD VDD p w=1.37u l=0.18u
M_u7-M_u2 net9 A1 X_u7-net8 VDD p w=1.37u l=0.18u
.ends
.subckt GSDFCNQD1BWP7T SI D SE CP CDN Q VDD VSS 
MI150 net62 net098 net070 VSS n w=1u l=0.18u
MI149 d1 CP net070 VSS n w=1u l=0.18u
MI165 net63 CDN VSS VSS n w=1u l=0.18u
MI164 net82 d1 net63 VSS n w=1u l=0.18u
MI47 d0 CP net82 VSS n w=1u l=0.18u
MI169 net177 net120 net69 VSS n w=1u l=0.18u
MI77 d0 INCPB net177 VSS n w=1u l=0.18u
MI161 net67 SI VSS VSS n w=1u l=0.18u
MI160 net177 SE net67 VSS n w=1u l=0.18u
MI158-M_u4 XI158-net6 net070 VSS VSS n w=1u l=0.18u
MI158-M_u3 d3 CDN XI158-net6 VSS n w=1u l=0.18u
MI166-M_u2 INCPB CP VSS VSS n w=1u l=0.18u
MI174-M_u2 net098 CP VSS VSS n w=1u l=0.18u
MI152-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI153-M_u2 net62 d3 VSS VSS n w=1u l=0.18u
MI85-M_u2 d1 d0 VSS VSS n w=1u l=0.18u
MI173-M_u2 net69 D VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=1u l=0.18u
MI158-M_u2 d3 net070 VDD VDD p w=1.37u l=0.18u
MI158-M_u1 d3 CDN VDD VDD p w=1.37u l=0.18u
MI166-M_u3 INCPB CP VDD VDD p w=1.37u l=0.18u
MI174-M_u3 net098 CP VDD VDD p w=1.37u l=0.18u
MI152-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI153-M_u3 net62 d3 VDD VDD p w=1.37u l=0.18u
MI85-M_u3 d1 d0 VDD VDD p w=1.37u l=0.18u
MI173-M_u3 net69 D VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=1.37u l=0.18u
MI155 net62 CP net070 VDD p w=1.37u l=0.18u
MI170 net132 SE net69 VDD p w=1.37u l=0.18u
MI163 d0 INCPB net166 VDD p w=1.37u l=0.18u
MI162 net166 d1 VDD VDD p w=1.37u l=0.18u
MI71 net132 net120 net142 VDD p w=1.37u l=0.18u
MI74 d0 CP net132 VDD p w=1.37u l=0.18u
MI75 net142 SI VDD VDD p w=1.37u l=0.18u
MI44 net166 CDN VDD VDD p w=1.37u l=0.18u
MI154 d1 net098 net070 VDD p w=1.37u l=0.18u
.ends
.subckt GTIEHBWP7T Z VDD VSS 
MI1 net6 net6 VSS VSS n w=1u l=0.18u
M_u2 net6 net6 VSS VSS n w=1u l=0.18u
MI0 Z net6 VDD VDD p w=1.37u l=0.18u
M_u1 Z net6 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GTIELBWP7T ZN VDD VSS 
MI1 ZN net6 VSS VSS n w=1u l=0.18u
M_u2 ZN net6 VSS VSS n w=1u l=0.18u
MI0 net6 net6 VDD VDD p w=1.37u l=0.18u
M_u1 net6 net6 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GXNR2D1BWP7T A1 A2 ZN VDD VSS 
M_u6-M_u2 net4 A1 net14 VSS n w=1u l=0.18u
MI57 net14 net10 net025 VSS n w=1u l=0.18u
MI58 net025 net4 VSS VSS n w=1u l=0.18u
M_u2-M_u2 net4 A2 VSS VSS n w=1u l=0.18u
M_u4-M_u2 ZN net14 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net10 A1 VSS VSS n w=1u l=0.18u
M_u6-M_u3 net4 net10 net14 VDD p w=1.37u l=0.18u
M_u2-M_u3 net4 A2 VDD VDD p w=1.37u l=0.18u
M_u4-M_u3 ZN net14 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net10 A1 VDD VDD p w=1.37u l=0.18u
MI61 net018 net4 VDD VDD p w=1.37u l=0.18u
MI60 net14 A1 net018 VDD p w=1.37u l=0.18u
.ends
.subckt GXNR2D2BWP7T A1 A2 ZN VDD VSS 
M_u6-M_u2 net4 A1 net14 VSS n w=1u l=0.18u
MI57 net14 net10 net017 VSS n w=1u l=0.18u
MI58 net017 net4 VSS VSS n w=1u l=0.18u
MI0-M_u2 net4 A2 VSS VSS n w=1u l=0.18u
M_u2-M_u2 net4 A2 VSS VSS n w=1u l=0.18u
M_u4_0-M_u2 ZN net14 VSS VSS n w=1u l=0.18u
M_u4_1-M_u2 ZN net14 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net10 A1 VSS VSS n w=1u l=0.18u
M_u6-M_u3 net4 net10 net14 VDD p w=1.37u l=0.18u
MI61 net024 net4 VDD VDD p w=1.37u l=0.18u
MI60 net14 A1 net024 VDD p w=1.37u l=0.18u
MI0-M_u3 net4 A2 VDD VDD p w=1.37u l=0.18u
M_u2-M_u3 net4 A2 VDD VDD p w=1.37u l=0.18u
M_u4_0-M_u3 ZN net14 VDD VDD p w=1.37u l=0.18u
M_u4_1-M_u3 ZN net14 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net10 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt GXOR2D1BWP7T A1 A2 Z VDD VSS 
M_u6-M_u2 net4 net045 net14 VSS n w=1u l=0.18u
MI58 net024 net4 VSS VSS n w=1u l=0.18u
MI57 net14 A1 net024 VSS n w=1u l=0.18u
M_u2-M_u2 net4 A2 VSS VSS n w=1u l=0.18u
M_u4-M_u2 Z net14 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net045 A1 VSS VSS n w=1u l=0.18u
M_u6-M_u3 net4 A1 net14 VDD p w=1.37u l=0.18u
M_u2-M_u3 net4 A2 VDD VDD p w=1.37u l=0.18u
M_u4-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net045 A1 VDD VDD p w=1.37u l=0.18u
MI61 net018 net4 VDD VDD p w=1.37u l=0.18u
MI60 net14 net045 net018 VDD p w=1.37u l=0.18u
.ends
.subckt GXOR2D2BWP7T A1 A2 Z VDD VSS 
M_u6-M_u2 net4 net043 net14 VSS n w=1u l=0.18u
MI57 net14 A1 net024 VSS n w=1u l=0.18u
MI58 net024 net4 VSS VSS n w=1u l=0.18u
MI1-M_u2 net4 A2 VSS VSS n w=1u l=0.18u
M_u2-M_u2 net4 A2 VSS VSS n w=1u l=0.18u
M_u4_0-M_u2 Z net14 VSS VSS n w=1u l=0.18u
M_u4_1-M_u2 Z net14 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net043 A1 VSS VSS n w=1u l=0.18u
M_u6-M_u3 net4 A1 net14 VDD p w=1.37u l=0.18u
MI1-M_u3 net4 A2 VDD VDD p w=1.37u l=0.18u
M_u2-M_u3 net4 A2 VDD VDD p w=1.37u l=0.18u
M_u4_0-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
M_u4_1-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net043 A1 VDD VDD p w=1.37u l=0.18u
MI61 net017 net4 VDD VDD p w=1.37u l=0.18u
MI60 net14 net043 net017 VDD p w=1.37u l=0.18u
.ends
.subckt HA1D0BWP7T A B S CO VDD VSS 
MI2 net21 B net023 VSS n w=0.62u l=0.18u
MI3 net023 net11 VSS VSS n w=0.88u l=0.18u
MU9-M_u4 XU9-net6 B VSS VSS n w=0.685u l=0.18u
MU9-M_u3 net23 A XU9-net6 VSS n w=0.685u l=0.18u
MU4-M_u2 S net21 VSS VSS n w=0.5u l=0.18u
MU3-M_u2 net7 B VSS VSS n w=0.5u l=0.18u
MU1-M_u2 net11 A VSS VSS n w=1u l=0.18u
MU5-M_u2 CO net23 VSS VSS n w=0.5u l=0.18u
MU8-M_u2 net11 net7 net21 VSS n w=0.55u l=0.18u
MI0 net034 net11 VDD VDD p w=1.37u l=0.18u
MI6 net21 net7 net034 VDD p w=1.37u l=0.18u
MU9-M_u2 net23 B VDD VDD p w=0.685u l=0.18u
MU9-M_u1 net23 A VDD VDD p w=0.685u l=0.18u
MU4-M_u3 S net21 VDD VDD p w=0.685u l=0.18u
MU3-M_u3 net7 B VDD VDD p w=0.685u l=0.18u
MU1-M_u3 net11 A VDD VDD p w=1.37u l=0.18u
MU5-M_u3 CO net23 VDD VDD p w=0.685u l=0.18u
MU8-M_u3 net11 B net21 VDD p w=0.92u l=0.18u
.ends
.subckt HA1D1BWP7T A B S CO VDD VSS 
MU8-M_u2 net11 net042 net21 VSS n w=0.55u l=0.18u
MI2 net21 B net036 VSS n w=0.62u l=0.18u
MI3 net036 net11 VSS VSS n w=0.88u l=0.18u
MU9-M_u4 XU9-net6 B VSS VSS n w=1u l=0.18u
MU9-M_u3 net23 A XU9-net6 VSS n w=1u l=0.18u
MU3-M_u2 net042 B VSS VSS n w=0.5u l=0.18u
MU4-M_u2 S net21 VSS VSS n w=1u l=0.18u
MU1_0-M_u2 net11 A VSS VSS n w=1u l=0.18u
MU1_1-M_u2 net11 A VSS VSS n w=1u l=0.18u
MU5-M_u2 CO net23 VSS VSS n w=1u l=0.18u
MU8-M_u3 net11 B net21 VDD p w=0.92u l=0.18u
MI0 net029 net11 VDD VDD p w=1.37u l=0.18u
MI6 net21 net042 net029 VDD p w=1.37u l=0.18u
MU9-M_u2 net23 B VDD VDD p w=1.37u l=0.18u
MU9-M_u1 net23 A VDD VDD p w=1.28u l=0.18u
MU3-M_u3 net042 B VDD VDD p w=0.685u l=0.18u
MU4-M_u3 S net21 VDD VDD p w=1.37u l=0.18u
MU1_0-M_u3 net11 A VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 net11 A VDD VDD p w=1.37u l=0.18u
MU5-M_u3 CO net23 VDD VDD p w=1.37u l=0.18u
.ends
.subckt HA1D2BWP7T A B S CO VDD VSS 
MI20 net38 B net025 VSS n w=0.62u l=0.18u
MI21 net025 net39 VSS VSS n w=0.88u l=0.18u
MU9-M_u4 XU9-net6 B VSS VSS n w=1u l=0.18u
MU9-M_u3 net23 A XU9-net6 VSS n w=1u l=0.18u
MU4_0-M_u2 S net38 VSS VSS n w=1u l=0.18u
MU4_1-M_u2 S net38 VSS VSS n w=1u l=0.18u
MU3-M_u2 net36 B VSS VSS n w=0.5u l=0.18u
MU1_0-M_u2 net39 A VSS VSS n w=1u l=0.18u
MU1_1-M_u2 net39 A VSS VSS n w=1u l=0.18u
MU5_0-M_u2 CO net23 VSS VSS n w=1u l=0.18u
MU5_1-M_u2 CO net23 VSS VSS n w=1u l=0.18u
MI1-M_u2 net39 net36 net38 VSS n w=0.55u l=0.18u
MI19 VDD net39 net030 VDD p w=1.37u l=0.18u
MI18 net030 net36 net38 VDD p w=1.37u l=0.18u
MU9-M_u2 net23 B VDD VDD p w=1.37u l=0.18u
MU9-M_u1 net23 A VDD VDD p w=1.28u l=0.18u
MU4_0-M_u3 S net38 VDD VDD p w=1.37u l=0.18u
MU4_1-M_u3 S net38 VDD VDD p w=1.37u l=0.18u
MU3-M_u3 net36 B VDD VDD p w=0.685u l=0.18u
MU1_0-M_u3 net39 A VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 net39 A VDD VDD p w=1.37u l=0.18u
MU5_0-M_u3 CO net23 VDD VDD p w=1.37u l=0.18u
MU5_1-M_u3 CO net23 VDD VDD p w=1.37u l=0.18u
MI1-M_u3 net39 B net38 VDD p w=0.92u l=0.18u
.ends
.subckt IAO21D0BWP7T A1 A2 B ZN VDD VSS 
MU37-M_u4 net11 A1 VSS VSS n w=0.42u l=0.18u
MU37-M_u3 net11 A2 VSS VSS n w=0.42u l=0.18u
MU39-M_u4 ZN B VSS VSS n w=0.5u l=0.18u
MU39-M_u3 ZN net11 VSS VSS n w=0.5u l=0.18u
MU37-M_u1 XU37-net8 A2 VDD VDD p w=0.42u l=0.18u
MU37-M_u2 net11 A1 XU37-net8 VDD p w=0.42u l=0.18u
MU39-M_u1 XU39-net8 net11 VDD VDD p w=0.685u l=0.18u
MU39-M_u2 ZN B XU39-net8 VDD p w=0.685u l=0.18u
.ends
.subckt IAO21D1BWP7T A1 A2 B ZN VDD VSS 
MU37-M_u4 net11 A1 VSS VSS n w=0.57u l=0.18u
MU37-M_u3 net11 A2 VSS VSS n w=0.57u l=0.18u
MU39-M_u4 ZN B VSS VSS n w=1u l=0.18u
MU39-M_u3 ZN net11 VSS VSS n w=1u l=0.18u
MU37-M_u1 XU37-net8 A2 VDD VDD p w=0.81u l=0.18u
MU37-M_u2 net11 A1 XU37-net8 VDD p w=0.81u l=0.18u
MU39-M_u1 XU39-net8 net11 VDD VDD p w=1.37u l=0.18u
MU39-M_u2 ZN B XU39-net8 VDD p w=1.37u l=0.18u
.ends
.subckt IAO21D2BWP7T A1 A2 B ZN VDD VSS 
MU37-M_u4 net11 A1 VSS VSS n w=1u l=0.18u
MU37-M_u3 net11 A2 VSS VSS n w=1u l=0.18u
MU39_0-M_u4 ZN B VSS VSS n w=1u l=0.18u
MU39_0-M_u3 ZN net11 VSS VSS n w=1u l=0.18u
MU39_1-M_u4 ZN B VSS VSS n w=1u l=0.18u
MU39_1-M_u3 ZN net11 VSS VSS n w=1u l=0.18u
MU37-M_u1 XU37-net8 A2 VDD VDD p w=1.37u l=0.18u
MU37-M_u2 net11 A1 XU37-net8 VDD p w=1.37u l=0.18u
MU39_0-M_u1 XU39_0-net8 net11 VDD VDD p w=1.37u l=0.18u
MU39_0-M_u2 ZN B XU39_0-net8 VDD p w=1.37u l=0.18u
MU39_1-M_u1 XU39_1-net8 net11 VDD VDD p w=1.37u l=0.18u
MU39_1-M_u2 ZN B XU39_1-net8 VDD p w=1.37u l=0.18u
.ends
.subckt IAO22D0BWP7T A1 A2 B1 B2 ZN VDD VSS 
MU37-M_u4 net42 A1 VSS VSS n w=0.42u l=0.18u
MU37-M_u3 net42 A2 VSS VSS n w=0.42u l=0.18u
MI2 ZN B1 net34 VSS n w=0.5u l=0.18u
MI3 net34 B2 VSS VSS n w=0.5u l=0.18u
M_u7 ZN net42 VSS VSS n w=0.5u l=0.18u
MU37-M_u1 XU37-net8 A2 VDD VDD p w=0.42u l=0.18u
MU37-M_u2 net42 A1 XU37-net8 VDD p w=0.42u l=0.18u
M_u4 net32 net42 ZN VDD p w=0.685u l=0.18u
M_u2 net32 B1 VDD VDD p w=0.685u l=0.18u
M_u3 VDD B2 net32 VDD p w=0.685u l=0.18u
.ends
.subckt IAO22D1BWP7T A1 A2 B1 B2 ZN VDD VSS 
MU37-M_u4 net42 A1 VSS VSS n w=0.77u l=0.18u
MU37-M_u3 net42 A2 VSS VSS n w=0.77u l=0.18u
MI2 ZN B1 net34 VSS n w=1u l=0.18u
MI3 net34 B2 VSS VSS n w=1u l=0.18u
M_u7 ZN net42 VSS VSS n w=1u l=0.18u
MU37-M_u1 XU37-net8 A2 VDD VDD p w=1.17u l=0.18u
MU37-M_u2 net42 A1 XU37-net8 VDD p w=1.17u l=0.18u
M_u4 net32 net42 ZN VDD p w=1.37u l=0.18u
M_u2 net32 B1 VDD VDD p w=1.37u l=0.18u
M_u3 VDD B2 net32 VDD p w=1.37u l=0.18u
.ends
.subckt IAO22D2BWP7T A1 A2 B1 B2 ZN VDD VSS 
MU52 net32 net6 net23 VSS n w=1u l=0.18u
MU54 net23 A1 VSS VSS n w=1u l=0.18u
MU53 net23 A2 VSS VSS n w=1u l=0.18u
MU50-M_u4 XU50-net6 B1 VSS VSS n w=0.5u l=0.18u
MU50-M_u3 net6 B2 XU50-net6 VSS n w=0.5u l=0.18u
MU51_0-M_u2 ZN net32 VSS VSS n w=1u l=0.18u
MU51_1-M_u2 ZN net32 VSS VSS n w=1u l=0.18u
MU50-M_u2 net6 B1 VDD VDD p w=0.685u l=0.18u
MU50-M_u1 net6 B2 VDD VDD p w=0.685u l=0.18u
MU51_0-M_u3 ZN net32 VDD VDD p w=1.37u l=0.18u
MU51_1-M_u3 ZN net32 VDD VDD p w=1.37u l=0.18u
MI16-MI12 net32 A2 XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 A1 VDD VDD p w=1.37u l=0.18u
MU47 net32 net6 VDD VDD p w=1.37u l=0.18u
.ends
.subckt IIND4D0BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI21-M_u5 ZN net25 XI21-net23 VSS n w=0.5u l=0.18u
MI21-M_u6 XI21-net23 B1 XI21-net26 VSS n w=0.5u l=0.18u
MI21-M_u7 XI21-net26 B2 XI21-net29 VSS n w=0.5u l=0.18u
MI21-M_u8 XI21-net29 net23 VSS VSS n w=0.5u l=0.18u
MI19-M_u2 net25 A1 VSS VSS n w=0.42u l=0.18u
MI20-M_u2 net23 A2 VSS VSS n w=0.42u l=0.18u
MI21-M_u4 ZN net23 VDD VDD p w=0.685u l=0.18u
MI21-M_u3 ZN B2 VDD VDD p w=0.685u l=0.18u
MI21-M_u2 ZN B1 VDD VDD p w=0.685u l=0.18u
MI21-M_u1 ZN net25 VDD VDD p w=0.685u l=0.18u
MI19-M_u3 net25 A1 VDD VDD p w=0.42u l=0.18u
MI20-M_u3 net23 A2 VDD VDD p w=0.42u l=0.18u
.ends
.subckt IIND4D1BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI21-M_u5 ZN net25 XI21-net23 VSS n w=1u l=0.18u
MI21-M_u6 XI21-net23 B1 XI21-net26 VSS n w=1u l=0.18u
MI21-M_u7 XI21-net26 B2 XI21-net29 VSS n w=1u l=0.18u
MI21-M_u8 XI21-net29 net23 VSS VSS n w=1u l=0.18u
MI19-M_u2 net25 A1 VSS VSS n w=0.5u l=0.18u
MI20-M_u2 net23 A2 VSS VSS n w=0.5u l=0.18u
MI21-M_u4 ZN net23 VDD VDD p w=1.37u l=0.18u
MI21-M_u3 ZN B2 VDD VDD p w=1.37u l=0.18u
MI21-M_u2 ZN B1 VDD VDD p w=1.37u l=0.18u
MI21-M_u1 ZN net25 VDD VDD p w=1.37u l=0.18u
MI19-M_u3 net25 A1 VDD VDD p w=0.685u l=0.18u
MI20-M_u3 net23 A2 VDD VDD p w=0.685u l=0.18u
.ends
.subckt IIND4D2BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI25-M_u2 net97 A2 VSS VSS n w=1u l=0.18u
MI24-M_u2 net48 A1 VSS VSS n w=1u l=0.18u
MI29 net044 B1 net048 VSS n w=2u l=0.18u
MU53 ZN net48 net044 VSS n w=2u l=0.18u
MI30 net048 B2 net047 VSS n w=2u l=0.18u
MI31 net047 net97 VSS VSS n w=2u l=0.18u
MI25-M_u3 net97 A2 VDD VDD p w=1.37u l=0.18u
MI24-M_u3 net48 A1 VDD VDD p w=1.37u l=0.18u
MI27_0 ZN B1 VDD VDD p w=1.37u l=0.18u
MI27_1 ZN B1 VDD VDD p w=1.37u l=0.18u
MI2_0 ZN net97 VDD VDD p w=1.37u l=0.18u
MI2_1 ZN net97 VDD VDD p w=1.37u l=0.18u
MI26_0 ZN B2 VDD VDD p w=1.37u l=0.18u
MI26_1 ZN B2 VDD VDD p w=1.37u l=0.18u
MI28_0 ZN net48 VDD VDD p w=1.37u l=0.18u
MI28_1 ZN net48 VDD VDD p w=1.37u l=0.18u
.ends
.subckt IINR4D0BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI27 ZN B1 VSS VSS n w=0.5u l=0.18u
MI16 ZN net42 VSS VSS n w=0.5u l=0.18u
MI28 ZN B2 VSS VSS n w=0.5u l=0.18u
MI26 ZN net33 VSS VSS n w=0.5u l=0.18u
MI29-M_u2 net33 A2 VSS VSS n w=0.42u l=0.18u
MI11-M_u2 net42 A1 VSS VSS n w=0.42u l=0.18u
MI29-M_u3 net33 A2 VDD VDD p w=0.42u l=0.18u
MI11-M_u3 net42 A1 VDD VDD p w=0.42u l=0.18u
MI22 p0 B2 VDD VDD p w=1.37u l=0.18u
MI24 p2 net33 p1 VDD p w=1.37u l=0.18u
MI23 p1 B1 p0 VDD p w=1.37u l=0.18u
MI25 ZN net42 p2 VDD p w=1.37u l=0.18u
.ends
.subckt IINR4D1BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI25 ZN B2 VSS VSS n w=1u l=0.18u
MI16 ZN net43 VSS VSS n w=1u l=0.18u
MI23 ZN net41 VSS VSS n w=0.7u l=0.18u
MI24 ZN B1 VSS VSS n w=1u l=0.18u
MI36-M_u2 net43 A1 VSS VSS n w=0.5u l=0.18u
MI37-M_u2 net41 A2 VSS VSS n w=0.5u l=0.18u
MI36-M_u3 net43 A1 VDD VDD p w=0.685u l=0.18u
MI37-M_u3 net41 A2 VDD VDD p w=0.685u l=0.18u
MI22 net68 B2 VDD VDD p w=1.37u l=0.18u
MI32 net55 B2 VDD VDD p w=1.37u l=0.18u
MI27 net58 net41 net49 VDD p w=1.37u l=0.18u
MI26 net49 B1 net68 VDD p w=1.37u l=0.18u
MI31 net54 B1 net55 VDD p w=1.37u l=0.18u
MI28 ZN net43 net58 VDD p w=1.37u l=0.18u
MI29 ZN net43 net48 VDD p w=1.37u l=0.18u
MI30 net48 net41 net54 VDD p w=1.37u l=0.18u
.ends
.subckt IINR4D2BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI38_0 ZN B2 VSS VSS n w=1u l=0.18u
MI38_1 ZN B2 VSS VSS n w=1u l=0.18u
MI37_0 ZN B1 VSS VSS n w=1u l=0.18u
MI37_1 ZN B1 VSS VSS n w=1u l=0.18u
MI16_0 ZN net39 VSS VSS n w=1u l=0.18u
MI16_1 ZN net39 VSS VSS n w=1u l=0.18u
MI36_0 ZN net22 VSS VSS n w=1u l=0.18u
MI36_1 ZN net22 VSS VSS n w=1u l=0.18u
MI49-M_u2 net39 A1 VSS VSS n w=1u l=0.18u
MI50-M_u2 net22 A2 VSS VSS n w=1u l=0.18u
MI49-M_u3 net39 A1 VDD VDD p w=1.37u l=0.18u
MI50-M_u3 net22 A2 VDD VDD p w=1.37u l=0.18u
MI39 net55 B2 VDD VDD p w=5.48u l=0.18u
MI40 net59 B1 net55 VDD p w=5.48u l=0.18u
MI41 ZN net39 net58 VDD p w=5.48u l=0.18u
MI42 net58 net22 net59 VDD p w=5.48u l=0.18u
.ends
.subckt IND2D0BWP7T A1 B1 ZN VDD VSS 
MI2-M_u2 net13 A1 VSS VSS n w=0.42u l=0.18u
MI13 net16 net13 VSS VSS n w=0.5u l=0.18u
MI12 ZN B1 net16 VSS n w=0.5u l=0.18u
MI2-M_u3 net13 A1 VDD VDD p w=0.42u l=0.18u
M_u16 VDD net13 ZN VDD p w=0.685u l=0.18u
MI11 VDD B1 ZN VDD p w=0.685u l=0.18u
.ends
.subckt IND2D1BWP7T A1 B1 ZN VDD VSS 
MI2-M_u2 net13 A1 VSS VSS n w=0.5u l=0.18u
MI13 net16 net13 VSS VSS n w=1u l=0.18u
MI12 ZN B1 net16 VSS n w=1u l=0.18u
MI2-M_u3 net13 A1 VDD VDD p w=0.685u l=0.18u
M_u16 VDD net13 ZN VDD p w=1.37u l=0.18u
MI11 VDD B1 ZN VDD p w=1.37u l=0.18u
.ends
.subckt IND2D2BWP7T A1 B1 ZN VDD VSS 
MI13-M_u2 net017 A1 VSS VSS n w=1u l=0.18u
MI10 ZN B1 net20 VSS n w=1u l=0.18u
MI11 net20 net017 VSS VSS n w=1u l=0.18u
MI4 net22 net017 VSS VSS n w=1u l=0.18u
MI12 ZN B1 net22 VSS n w=1u l=0.18u
MI13-M_u3 net017 A1 VDD VDD p w=1.37u l=0.18u
M_u16 VDD net017 ZN VDD p w=2.74u l=0.18u
MI3 VDD B1 ZN VDD p w=2.74u l=0.18u
.ends
.subckt IND2D4BWP7T A1 B1 ZN VDD VSS 
MI2_0-M_u2 p0 A1 VSS VSS n w=1u l=0.18u
MI2_1-M_u2 p0 A1 VSS VSS n w=1u l=0.18u
MI7 ZN B1 net26 VSS n w=1u l=0.18u
MI8 net29 p0 VSS VSS n w=1u l=0.18u
MI9 net26 p0 VSS VSS n w=1u l=0.18u
MI10 ZN B1 net29 VSS n w=1u l=0.18u
MI5 ZN B1 net41 VSS n w=1u l=0.18u
MI13 net38 p0 VSS VSS n w=1u l=0.18u
MI4 net41 p0 VSS VSS n w=1u l=0.18u
MI12 ZN B1 net38 VSS n w=1u l=0.18u
MI2_0-M_u3 p0 A1 VDD VDD p w=1.37u l=0.18u
MI2_1-M_u3 p0 A1 VDD VDD p w=1.37u l=0.18u
M_u16_0 VDD p0 ZN VDD p w=1.37u l=0.18u
M_u16_1 VDD p0 ZN VDD p w=1.37u l=0.18u
M_u16_2 VDD p0 ZN VDD p w=1.37u l=0.18u
M_u16_3 VDD p0 ZN VDD p w=1.37u l=0.18u
MI11_0 VDD B1 ZN VDD p w=1.37u l=0.18u
MI11_1 VDD B1 ZN VDD p w=1.37u l=0.18u
MI11_2 VDD B1 ZN VDD p w=1.37u l=0.18u
MI11_3 VDD B1 ZN VDD p w=1.37u l=0.18u
.ends
.subckt IND3D0BWP7T A1 B1 B2 ZN VDD VSS 
MI5-M_u2 net30 A1 VSS VSS n w=0.42u l=0.18u
MI12 ZN B2 net23 VSS n w=0.5u l=0.18u
MI11 net20 net30 VSS VSS n w=0.5u l=0.18u
MI10 net23 B1 net20 VSS n w=0.5u l=0.18u
MI5-M_u3 net30 A1 VDD VDD p w=0.42u l=0.18u
MI9 VDD B2 ZN VDD p w=0.685u l=0.18u
MI8 VDD B1 ZN VDD p w=0.685u l=0.18u
MI4 VDD net30 ZN VDD p w=0.685u l=0.18u
.ends
.subckt IND3D1BWP7T A1 B1 B2 ZN VDD VSS 
MI5-M_u2 net30 A1 VSS VSS n w=0.5u l=0.18u
MI12 ZN B2 net23 VSS n w=1u l=0.18u
MI7 net20 net30 VSS VSS n w=1u l=0.18u
MI6 net23 B1 net20 VSS n w=1u l=0.18u
MI5-M_u3 net30 A1 VDD VDD p w=0.685u l=0.18u
MI11 VDD B2 ZN VDD p w=1.37u l=0.18u
M_u16 VDD B1 ZN VDD p w=0.835u l=0.18u
MI4 VDD net30 ZN VDD p w=1.37u l=0.18u
.ends
.subckt IND3D2BWP7T A1 B1 B2 ZN VDD VSS 
MI5-M_u2 net30 A1 VSS VSS n w=1u l=0.18u
MI17 net32 B1 net29 VSS n w=2u l=0.18u
MI16 net29 net30 VSS VSS n w=2u l=0.18u
MI18 ZN B2 net32 VSS n w=2u l=0.18u
MI5-M_u3 net30 A1 VDD VDD p w=1.37u l=0.18u
MI9_0 VDD B2 ZN VDD p w=1.37u l=0.18u
MI9_1 VDD B2 ZN VDD p w=1.37u l=0.18u
MI8_0 VDD B1 ZN VDD p w=1.37u l=0.18u
MI8_1 VDD B1 ZN VDD p w=1.37u l=0.18u
MI4_0 VDD net30 ZN VDD p w=1.37u l=0.18u
MI4_1 VDD net30 ZN VDD p w=1.37u l=0.18u
.ends
.subckt IND4D0BWP7T A1 B1 B2 B3 ZN VDD VSS 
MI11-M_u2 net20 A1 VSS VSS n w=0.42u l=0.18u
MU53 ZN B3 p0 VSS n w=0.5u l=0.18u
MI17 p2 net20 VSS VSS n w=0.5u l=0.18u
MI16 p1 B1 p2 VSS n w=0.5u l=0.18u
MI15 p0 B2 p1 VSS n w=0.5u l=0.18u
MI11-M_u3 net20 A1 VDD VDD p w=0.42u l=0.18u
MI12 ZN B1 VDD VDD p w=0.685u l=0.18u
MI14 ZN B3 VDD VDD p w=0.685u l=0.18u
MI13 ZN B2 VDD VDD p w=0.685u l=0.18u
MI18 ZN net20 VDD VDD p w=0.685u l=0.18u
.ends
.subckt IND4D1BWP7T A1 B1 B2 B3 ZN VDD VSS 
MI11-M_u2 net20 A1 VSS VSS n w=0.5u l=0.18u
MI10 p2 net20 VSS VSS n w=1u l=0.18u
MI8 p0 B2 p1 VSS n w=1u l=0.18u
MI9 p1 B1 p2 VSS n w=1u l=0.18u
MU53 ZN B3 p0 VSS n w=1u l=0.18u
MI11-M_u3 net20 A1 VDD VDD p w=0.685u l=0.18u
MI18 ZN net20 VDD VDD p w=1.37u l=0.18u
MI5 ZN B1 VDD VDD p w=1.37u l=0.18u
MI6 ZN B2 VDD VDD p w=1.37u l=0.18u
MI7 ZN B3 VDD VDD p w=1.37u l=0.18u
.ends
.subckt IND4D2BWP7T A1 B1 B2 B3 ZN VDD VSS 
MI11-M_u2 net020 A1 VSS VSS n w=1u l=0.18u
MU53 ZN B3 p0 VSS n w=2u l=0.18u
MI21 p0 B2 p1 VSS n w=2u l=0.18u
MI22 p1 B1 p2 VSS n w=2u l=0.18u
MI23 p2 net020 VSS VSS n w=2u l=0.18u
MI11-M_u3 net020 A1 VDD VDD p w=1.37u l=0.18u
MI19 ZN B2 VDD VDD p w=2.66u l=0.18u
MI18 ZN B1 VDD VDD p w=2.66u l=0.18u
MI17 ZN net020 VDD VDD p w=2.74u l=0.18u
MI20 ZN B3 VDD VDD p w=2.74u l=0.18u
.ends
.subckt INR2D0BWP7T A1 B1 ZN VDD VSS 
MU1-M_u4 ZN B1 VSS VSS n w=0.5u l=0.18u
MU1-M_u3 ZN net4 VSS VSS n w=0.5u l=0.18u
MU6-M_u2 net4 A1 VSS VSS n w=0.42u l=0.18u
MU1-M_u1 XU1-net8 net4 VDD VDD p w=0.685u l=0.18u
MU1-M_u2 ZN B1 XU1-net8 VDD p w=0.685u l=0.18u
MU6-M_u3 net4 A1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt INR2D1BWP7T A1 B1 ZN VDD VSS 
MU1-M_u4 ZN B1 VSS VSS n w=1u l=0.18u
MU1-M_u3 ZN net4 VSS VSS n w=1u l=0.18u
MU6-M_u2 net4 A1 VSS VSS n w=0.5u l=0.18u
MU1-M_u1 XU1-net8 net4 VDD VDD p w=1.37u l=0.18u
MU1-M_u2 ZN B1 XU1-net8 VDD p w=1.37u l=0.18u
MU6-M_u3 net4 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt INR2D2BWP7T A1 B1 ZN VDD VSS 
MU1_0-M_u4 ZN B1 VSS VSS n w=1u l=0.18u
MU1_0-M_u3 ZN net4 VSS VSS n w=1u l=0.18u
MU1_1-M_u4 ZN B1 VSS VSS n w=1u l=0.18u
MU1_1-M_u3 ZN net4 VSS VSS n w=1u l=0.18u
MU6-M_u2 net4 A1 VSS VSS n w=1u l=0.18u
MU1_0-M_u1 XU1_0-net8 net4 VDD VDD p w=1.37u l=0.18u
MU1_0-M_u2 ZN B1 XU1_0-net8 VDD p w=1.37u l=0.18u
MU1_1-M_u1 XU1_1-net8 net4 VDD VDD p w=1.37u l=0.18u
MU1_1-M_u2 ZN B1 XU1_1-net8 VDD p w=1.37u l=0.18u
MU6-M_u3 net4 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt INR2D4BWP7T A1 B1 ZN VDD VSS 
MI13 ZN p0 VSS VSS n w=1u l=0.18u
MI9 ZN B1 VSS VSS n w=1u l=0.18u
MI12 ZN p0 VSS VSS n w=1u l=0.18u
MI11 ZN p0 VSS VSS n w=1u l=0.18u
MI8 ZN B1 VSS VSS n w=1u l=0.18u
M_u4 ZN B1 VSS VSS n w=1u l=0.18u
MI10 ZN B1 VSS VSS n w=1u l=0.18u
M_u3 ZN p0 VSS VSS n w=1u l=0.18u
MU6_0-M_u2 p0 A1 VSS VSS n w=1u l=0.18u
MU6_1-M_u2 p0 A1 VSS VSS n w=1u l=0.18u
MI3 net052 p0 VDD VDD p w=1.37u l=0.18u
MI4 net043 p0 VDD VDD p w=1.37u l=0.18u
M_u1 net12 p0 VDD VDD p w=1.37u l=0.18u
M_u2 ZN B1 net12 VDD p w=1.37u l=0.18u
MI2 ZN B1 net052 VDD p w=1.37u l=0.18u
MI6 ZN B1 net040 VDD p w=1.37u l=0.18u
MI7 net040 p0 VDD VDD p w=1.37u l=0.18u
MI5 ZN B1 net043 VDD p w=1.37u l=0.18u
MU6_0-M_u3 p0 A1 VDD VDD p w=1.37u l=0.18u
MU6_1-M_u3 p0 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt INR2XD0BWP7T A1 B1 ZN VDD VSS 
MU1-M_u4 ZN B1 VSS VSS n w=0.5u l=0.18u
MU1-M_u3 ZN net4 VSS VSS n w=0.5u l=0.18u
MU6-M_u2 net4 A1 VSS VSS n w=0.5u l=0.18u
MU1-M_u1 XU1-net8 net4 VDD VDD p w=1.37u l=0.18u
MU1-M_u2 ZN B1 XU1-net8 VDD p w=1.37u l=0.18u
MU6-M_u3 net4 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt INR2XD1BWP7T A1 B1 ZN VDD VSS 
MU1-M_u4 ZN B1 VSS VSS n w=1u l=0.18u
MU1-M_u3 ZN net4 VSS VSS n w=1u l=0.18u
MU6-M_u2 net4 A1 VSS VSS n w=1u l=0.18u
MU1-M_u1 XU1-net8 net4 VDD VDD p w=2.74u l=0.18u
MU1-M_u2 ZN B1 XU1-net8 VDD p w=2.74u l=0.18u
MU6-M_u3 net4 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt INR2XD2BWP7T A1 B1 ZN VDD VSS 
MU1_0-M_u4 ZN B1 VSS VSS n w=0.5u l=0.18u
MU1_0-M_u3 ZN net4 VSS VSS n w=0.5u l=0.18u
MU1_1-M_u4 ZN B1 VSS VSS n w=0.5u l=0.18u
MU1_1-M_u3 ZN net4 VSS VSS n w=0.5u l=0.18u
MU1_2-M_u4 ZN B1 VSS VSS n w=0.5u l=0.18u
MU1_2-M_u3 ZN net4 VSS VSS n w=0.5u l=0.18u
MU1_3-M_u4 ZN B1 VSS VSS n w=0.5u l=0.18u
MU1_3-M_u3 ZN net4 VSS VSS n w=0.5u l=0.18u
MU6-M_u2 net4 A1 VSS VSS n w=1u l=0.18u
MU1_0-M_u1 XU1_0-net8 net4 VDD VDD p w=1.37u l=0.18u
MU1_0-M_u2 ZN B1 XU1_0-net8 VDD p w=1.37u l=0.18u
MU1_1-M_u1 XU1_1-net8 net4 VDD VDD p w=1.37u l=0.18u
MU1_1-M_u2 ZN B1 XU1_1-net8 VDD p w=1.37u l=0.18u
MU1_2-M_u1 XU1_2-net8 net4 VDD VDD p w=1.37u l=0.18u
MU1_2-M_u2 ZN B1 XU1_2-net8 VDD p w=1.37u l=0.18u
MU1_3-M_u1 XU1_3-net8 net4 VDD VDD p w=1.37u l=0.18u
MU1_3-M_u2 ZN B1 XU1_3-net8 VDD p w=1.37u l=0.18u
MU6-M_u3 net4 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt INR2XD4BWP7T A1 B1 ZN VDD VSS 
M_u2 ZN p0 VSS VSS n w=3.99u l=0.18u
MI14 ZN B1 VSS VSS n w=3.99u l=0.18u
MI5-M_u2 p0 A1 VSS VSS n w=2u l=0.18u
MI5-M_u3 p0 A1 VDD VDD p w=2.74u l=0.18u
MI12 net051 B1 VDD VDD p w=10.7u l=0.18u
MI13 ZN p0 net051 VDD p w=10.7u l=0.18u
.ends
.subckt INR3D0BWP7T A1 B1 B2 ZN VDD VSS 
MU9-M_u6 ZN B2 VSS VSS n w=0.5u l=0.18u
MU9-M_u5 ZN B1 VSS VSS n w=0.5u l=0.18u
MU9-M_u4 ZN net12 VSS VSS n w=0.5u l=0.18u
MU47-M_u2 net12 A1 VSS VSS n w=0.42u l=0.18u
MU9-M_u1 XU9-net9 net12 VDD VDD p w=1.37u l=0.18u
MU9-M_u2 XU9-net12 B1 XU9-net9 VDD p w=1.37u l=0.18u
MU9-M_u3 ZN B2 XU9-net12 VDD p w=1.37u l=0.18u
MU47-M_u3 net12 A1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt INR3D1BWP7T A1 B1 B2 ZN VDD VSS 
M_u4 ZN net12 VSS VSS n w=1u l=0.18u
MI3 ZN B1 VSS VSS n w=1u l=0.18u
MI4 ZN B2 VSS VSS n w=1u l=0.18u
MU47-M_u2 net12 A1 VSS VSS n w=1u l=0.18u
MU47-M_u3 net12 A1 VDD VDD p w=1.37u l=0.18u
MI7 net26 net12 VDD VDD p w=1.245u l=0.18u
MI6 net29 B1 net26 VDD p w=1.245u l=0.18u
M_u1 net35 net12 VDD VDD p w=1.245u l=0.18u
MI1 net32 B1 net35 VDD p w=1.245u l=0.18u
MI2 ZN B2 net32 VDD p w=1.245u l=0.18u
MI5 ZN B2 net29 VDD p w=1.245u l=0.18u
.ends
.subckt INR3D2BWP7T A1 B1 B2 ZN VDD VSS 
MU9-M_u6 ZN B2 VSS VSS n w=2u l=0.18u
MU9-M_u5 ZN B1 VSS VSS n w=2u l=0.18u
MU9-M_u4 ZN net16 VSS VSS n w=2u l=0.18u
MU47-M_u2 net16 A1 VSS VSS n w=1u l=0.18u
MU9-M_u1 XU9-net9 net16 VDD VDD p w=2.74u l=0.18u
MU9-M_u2 XU9-net12 B1 XU9-net9 VDD p w=2.74u l=0.18u
MU9-M_u3 ZN B2 XU9-net12 VDD p w=2.74u l=0.18u
MU47-M_u3 net16 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt INR4D0BWP7T A1 B1 B2 B3 ZN VDD VSS 
MU8-M_u4 ZN net15 VSS VSS n w=0.5u l=0.18u
MU8-M_u3 ZN B1 VSS VSS n w=0.5u l=0.18u
MU8-M_u5 ZN B2 VSS VSS n w=0.5u l=0.18u
MU8-M_u8 ZN B3 VSS VSS n w=0.5u l=0.18u
MU47-M_u2 net15 A1 VSS VSS n w=0.42u l=0.18u
MU8-M_u7 ZN B3 XU8-net7 VDD p w=1.37u l=0.18u
MU8-M_u6 XU8-net7 B2 XU8-net10 VDD p w=1.37u l=0.18u
MU8-M_u2 XU8-net10 B1 XU8-net13 VDD p w=1.37u l=0.18u
MU8-M_u1 XU8-net13 net15 VDD VDD p w=1.37u l=0.18u
MU47-M_u3 net15 A1 VDD VDD p w=0.42u l=0.18u
.ends
.subckt INR4D1BWP7T A1 B1 B2 B3 ZN VDD VSS 
MI3 ZN B2 VSS VSS n w=0.7u l=0.18u
MI2 ZN B1 VSS VSS n w=0.7u l=0.18u
MI1 ZN net039 VSS VSS n w=0.7u l=0.18u
MI5 ZN B3 VSS VSS n w=0.7u l=0.18u
MU47-M_u2 net039 A1 VSS VSS n w=0.5u l=0.18u
MU47-M_u3 net039 A1 VDD VDD p w=0.685u l=0.18u
MI28 ZN B3 net18 VDD p w=1.37u l=0.18u
MI26 net21 B1 net39 VDD p w=1.37u l=0.18u
MI30 net27 net039 net36 VDD p w=1.37u l=0.18u
MI31 net36 B1 net33 VDD p w=1.37u l=0.18u
MI32 net33 B2 VDD VDD p w=1.37u l=0.18u
MI29 ZN B3 net27 VDD p w=1.37u l=0.18u
MI7 net39 B2 VDD VDD p w=1.37u l=0.18u
MI27 net18 net039 net21 VDD p w=1.37u l=0.18u
.ends
.subckt INR4D2BWP7T A1 B1 B2 B3 ZN VDD VSS 
MI15_0 ZN net15 VSS VSS n w=1u l=0.18u
MI15_1 ZN net15 VSS VSS n w=1u l=0.18u
MI14_0 ZN B1 VSS VSS n w=1u l=0.18u
MI14_1 ZN B1 VSS VSS n w=1u l=0.18u
MI13_0 ZN B2 VSS VSS n w=1u l=0.18u
MI13_1 ZN B2 VSS VSS n w=1u l=0.18u
MI5_0 ZN B3 VSS VSS n w=1u l=0.18u
MI5_1 ZN B3 VSS VSS n w=1u l=0.18u
MU47-M_u2 net15 A1 VSS VSS n w=1u l=0.18u
MU47-M_u3 net15 A1 VDD VDD p w=1.37u l=0.18u
MI8 ZN B3 net18 VDD p w=5.48u l=0.18u
MI4 net21 B1 net39 VDD p w=5.48u l=0.18u
MI7 net39 net15 VDD VDD p w=5.48u l=0.18u
MI6 net18 B2 net21 VDD p w=5.48u l=0.18u
.ends
.subckt INVD0BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=0.5u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=0.685u l=0.18u
.ends
.subckt INVD10BWP7T I ZN VDD VSS 
MU1_0-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_1-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_2-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_3-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_4-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_5-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_6-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_7-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_8-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_9-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_0-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_2-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_3-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_4-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_5-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_6-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_7-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_8-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_9-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt INVD12BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=12u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=16.44u l=0.18u
.ends
.subckt INVD1BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt INVD1P5BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=1.5u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=2.055u l=0.18u
.ends
.subckt INVD2BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=2u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=2.74u l=0.18u
.ends
.subckt INVD2P5BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=2.465u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=3.425u l=0.18u
.ends
.subckt INVD3BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=3u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=4.11u l=0.18u
.ends
.subckt INVD4BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=4u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=5.48u l=0.18u
.ends
.subckt INVD5BWP7T I ZN VDD VSS 
MU1_0-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_1-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_2-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_3-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_4-M_u2 ZN I VSS VSS n w=1u l=0.18u
MU1_0-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_2-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_3-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
MU1_4-M_u3 ZN I VDD VDD p w=1.37u l=0.18u
.ends
.subckt INVD6BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=6u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=8.22u l=0.18u
.ends
.subckt INVD8BWP7T I ZN VDD VSS 
MU1-M_u2 ZN I VSS VSS n w=8u l=0.18u
MU1-M_u3 ZN I VDD VDD p w=10.96u l=0.18u
.ends
.subckt IOA21D0BWP7T A1 A2 B ZN VDD VSS 
MU35-M_u4 XU35-net6 A2 VSS VSS n w=0.42u l=0.18u
MU35-M_u3 net5 A1 XU35-net6 VSS n w=0.42u l=0.18u
MU36-M_u4 XU36-net6 net5 VSS VSS n w=0.5u l=0.18u
MU36-M_u3 ZN B XU36-net6 VSS n w=0.5u l=0.18u
MU35-M_u2 net5 A2 VDD VDD p w=0.42u l=0.18u
MU35-M_u1 net5 A1 VDD VDD p w=0.42u l=0.18u
MU36-M_u2 ZN net5 VDD VDD p w=0.685u l=0.18u
MU36-M_u1 ZN B VDD VDD p w=0.685u l=0.18u
.ends
.subckt IOA21D1BWP7T A1 A2 B ZN VDD VSS 
MU35-M_u4 XU35-net6 A2 VSS VSS n w=0.5u l=0.18u
MU35-M_u3 net5 A1 XU35-net6 VSS n w=0.5u l=0.18u
MU36-M_u4 XU36-net6 net5 VSS VSS n w=1u l=0.18u
MU36-M_u3 ZN B XU36-net6 VSS n w=1u l=0.18u
MU35-M_u2 net5 A2 VDD VDD p w=0.685u l=0.18u
MU35-M_u1 net5 A1 VDD VDD p w=0.685u l=0.18u
MU36-M_u2 ZN net5 VDD VDD p w=1.37u l=0.18u
MU36-M_u1 ZN B VDD VDD p w=1.37u l=0.18u
.ends
.subckt IOA21D2BWP7T A1 A2 B ZN VDD VSS 
MU35-M_u4 XU35-net6 A2 VSS VSS n w=1u l=0.18u
MU35-M_u3 net5 A1 XU35-net6 VSS n w=1u l=0.18u
MU36_0-M_u4 XU36_0-net6 net5 VSS VSS n w=1u l=0.18u
MU36_0-M_u3 ZN B XU36_0-net6 VSS n w=1u l=0.18u
MU36_1-M_u4 XU36_1-net6 net5 VSS VSS n w=1u l=0.18u
MU36_1-M_u3 ZN B XU36_1-net6 VSS n w=1u l=0.18u
MU35-M_u2 net5 A2 VDD VDD p w=1.37u l=0.18u
MU35-M_u1 net5 A1 VDD VDD p w=1.37u l=0.18u
MU36_0-M_u2 ZN net5 VDD VDD p w=1.37u l=0.18u
MU36_0-M_u1 ZN B VDD VDD p w=1.37u l=0.18u
MU36_1-M_u2 ZN net5 VDD VDD p w=1.37u l=0.18u
MU36_1-M_u1 ZN B VDD VDD p w=1.37u l=0.18u
.ends
.subckt IOA22D0BWP7T A1 A2 B1 B2 ZN VDD VSS 
MU26 ZN net6 net17 VSS n w=0.5u l=0.18u
MU29 net17 B2 VSS VSS n w=0.5u l=0.18u
MU24 net17 B1 VSS VSS n w=0.5u l=0.18u
MU35-M_u4 XU35-net6 A1 VSS VSS n w=0.42u l=0.18u
MU35-M_u3 net6 A2 XU35-net6 VSS n w=0.42u l=0.18u
MU35-M_u2 net6 A1 VDD VDD p w=0.42u l=0.18u
MU35-M_u1 net6 A2 VDD VDD p w=0.42u l=0.18u
MU30 ZN net6 VDD VDD p w=0.685u l=0.18u
MI16-MI12 ZN B2 XI16-net11 VDD p w=0.685u l=0.18u
MI16-MI13 XI16-net11 B1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt IOA22D1BWP7T A1 A2 B1 B2 ZN VDD VSS 
MU26 ZN net6 net17 VSS n w=1u l=0.18u
MU29 net17 B2 VSS VSS n w=1u l=0.18u
MU24 net17 B1 VSS VSS n w=1u l=0.18u
MU35-M_u4 XU35-net6 A1 VSS VSS n w=0.685u l=0.18u
MU35-M_u3 net6 A2 XU35-net6 VSS n w=0.685u l=0.18u
MU35-M_u2 net6 A1 VDD VDD p w=0.685u l=0.18u
MU35-M_u1 net6 A2 VDD VDD p w=0.685u l=0.18u
MU30 ZN net6 VDD VDD p w=1.37u l=0.18u
MI16-MI12 ZN B2 XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 B1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt IOA22D2BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI4 net27 A2 VSS VSS n w=1u l=0.18u
MI3 net30 A1 net27 VSS n w=1u l=0.18u
MU51 net30 net6 VSS VSS n w=1u l=0.18u
MU37_0-M_u2 ZN net30 VSS VSS n w=1u l=0.18u
MU37_1-M_u2 ZN net30 VSS VSS n w=1u l=0.18u
MU56-M_u4 net6 B1 VSS VSS n w=0.5u l=0.18u
MU56-M_u3 net6 B2 VSS VSS n w=0.5u l=0.18u
MU37_0-M_u3 ZN net30 VDD VDD p w=1.37u l=0.18u
MU37_1-M_u3 ZN net30 VDD VDD p w=1.37u l=0.18u
MU56-M_u1 XU56-net8 B2 VDD VDD p w=1.37u l=0.18u
MU56-M_u2 net6 B1 XU56-net8 VDD p w=1.37u l=0.18u
MI2 net30 net6 net16 VDD p w=1.37u l=0.18u
MU50 net16 A2 VDD VDD p w=1.37u l=0.18u
MI1 net16 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt LHCND1BWP7T D E CDN Q QN VDD VSS 
MI6 net46 net071 net45 VSS n w=0.535u l=0.18u
MI10 net51 CDN VSS VSS n w=0.42u l=0.18u
MI8 net45 D net40 VSS n w=0.535u l=0.18u
MI29 net48 net36 net51 VSS n w=0.42u l=0.18u
MI5 net46 net63 net48 VSS n w=0.42u l=0.18u
MI9 net40 CDN VSS VSS n w=0.78u l=0.18u
MI7-M_u2 net071 net63 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net61 net36 VSS VSS n w=1u l=0.18u
MI12-M_u2 QN net36 VSS VSS n w=1u l=0.18u
MI11-M_u2 Q net61 VSS VSS n w=1u l=0.18u
MI14-M_u2 net63 E VSS VSS n w=0.5u l=0.18u
MI4-M_u2 net36 net46 VSS VSS n w=1u l=0.18u
MI30 net46 CDN VDD VDD p w=0.685u l=0.18u
MI21 net46 net63 net70 VDD p w=0.975u l=0.18u
MI17 VDD net36 net73 VDD p w=0.42u l=0.18u
MI24 net70 D VDD VDD p w=0.975u l=0.18u
MI18 net46 net071 net73 VDD p w=0.42u l=0.18u
MI7-M_u3 net071 net63 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net61 net36 VDD VDD p w=1.37u l=0.18u
MI12-M_u3 QN net36 VDD VDD p w=1.37u l=0.18u
MI11-M_u3 Q net61 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net63 E VDD VDD p w=0.685u l=0.18u
MI4-M_u3 net36 net46 VDD VDD p w=1.37u l=0.18u
.ends
.subckt LHCND2BWP7T D E CDN Q QN VDD VSS 
MI6 net46 net077 net45 VSS n w=0.535u l=0.18u
MI10 net51 CDN VSS VSS n w=0.42u l=0.18u
MI8 net45 D net40 VSS n w=0.535u l=0.18u
MI29 net48 net36 net51 VSS n w=0.42u l=0.18u
MI5 net46 net63 net48 VSS n w=0.42u l=0.18u
MI9 net40 CDN VSS VSS n w=0.535u l=0.18u
MI7-M_u2 Q net61 VSS VSS n w=2u l=0.18u
MI13-M_u2 QN net36 VSS VSS n w=2u l=0.18u
MI15-M_u2 net077 net63 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net61 net36 VSS VSS n w=1u l=0.18u
MI14-M_u2 net63 E VSS VSS n w=0.5u l=0.18u
MI4-M_u2 net36 net46 VSS VSS n w=1u l=0.18u
MI30 net46 CDN VDD VDD p w=0.685u l=0.18u
MI21 net46 net63 net70 VDD p w=0.975u l=0.18u
MI17 VDD net36 net73 VDD p w=0.42u l=0.18u
MI24 net70 D VDD VDD p w=0.975u l=0.18u
MI18 net46 net077 net73 VDD p w=0.42u l=0.18u
MI7-M_u3 Q net61 VDD VDD p w=2.74u l=0.18u
MI13-M_u3 QN net36 VDD VDD p w=2.74u l=0.18u
MI15-M_u3 net077 net63 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net61 net36 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net63 E VDD VDD p w=0.685u l=0.18u
MI4-M_u3 net36 net46 VDD VDD p w=1.37u l=0.18u
.ends
.subckt LHCNQD1BWP7T D E CDN Q VDD VSS 
MI6 net46 net071 net45 VSS n w=0.535u l=0.18u
MI10 net51 CDN VSS VSS n w=0.42u l=0.18u
MI8 net45 D net40 VSS n w=0.535u l=0.18u
MI29 net48 net36 net51 VSS n w=0.42u l=0.18u
MI5 net46 net63 net48 VSS n w=0.42u l=0.18u
MI9 net40 CDN VSS VSS n w=0.78u l=0.18u
MI7-M_u2 net071 net63 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net61 net36 VSS VSS n w=1u l=0.18u
MI11-M_u2 Q net61 VSS VSS n w=1u l=0.18u
MI14-M_u2 net63 E VSS VSS n w=0.5u l=0.18u
MI4-M_u2 net36 net46 VSS VSS n w=1u l=0.18u
MI30 net46 CDN VDD VDD p w=0.685u l=0.18u
MI21 net46 net63 net70 VDD p w=0.975u l=0.18u
MI17 VDD net36 net73 VDD p w=0.42u l=0.18u
MI24 net70 D VDD VDD p w=0.975u l=0.18u
MI18 net46 net071 net73 VDD p w=0.42u l=0.18u
MI7-M_u3 net071 net63 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net61 net36 VDD VDD p w=1.37u l=0.18u
MI11-M_u3 Q net61 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net63 E VDD VDD p w=0.685u l=0.18u
MI4-M_u3 net36 net46 VDD VDD p w=1.37u l=0.18u
.ends
.subckt LHCNQD2BWP7T D E CDN Q VDD VSS 
MI6 net46 net077 net45 VSS n w=0.535u l=0.18u
MI10 net51 CDN VSS VSS n w=0.42u l=0.18u
MI8 net45 D net40 VSS n w=0.535u l=0.18u
MI29 net48 net36 net51 VSS n w=0.42u l=0.18u
MI5 net46 net63 net48 VSS n w=0.42u l=0.18u
MI9 net40 CDN VSS VSS n w=0.535u l=0.18u
MI7-M_u2 Q net61 VSS VSS n w=2u l=0.18u
MI15-M_u2 net077 net63 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net61 net36 VSS VSS n w=1u l=0.18u
MI14-M_u2 net63 E VSS VSS n w=0.5u l=0.18u
MI4-M_u2 net36 net46 VSS VSS n w=1u l=0.18u
MI30 net46 CDN VDD VDD p w=0.685u l=0.18u
MI21 net46 net63 net70 VDD p w=0.975u l=0.18u
MI17 VDD net36 net73 VDD p w=0.42u l=0.18u
MI24 net70 D VDD VDD p w=0.975u l=0.18u
MI18 net46 net077 net73 VDD p w=0.42u l=0.18u
MI7-M_u3 Q net61 VDD VDD p w=2.74u l=0.18u
MI15-M_u3 net077 net63 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net61 net36 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net63 E VDD VDD p w=0.685u l=0.18u
MI4-M_u3 net36 net46 VDD VDD p w=1.37u l=0.18u
.ends
.subckt LHD1BWP7T D E Q QN VDD VSS 
MI2-M_u2 net11 E VSS VSS n w=0.5u l=0.18u
MU24-M_u2 QN net20 VSS VSS n w=1u l=0.18u
MU23-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU29-M_u2 net34 net11 VSS VSS n w=0.5u l=0.18u
MU30-M_u2 net20 net15 VSS VSS n w=1u l=0.18u
MU32-MU3 net15 net34 XU32-net16 VSS n w=0.68u l=0.18u
MU32-MU4 XU32-net16 D VSS VSS n w=0.78u l=0.18u
MU22-MU3 net15 net11 XU22-net16 VSS n w=0.42u l=0.18u
MU22-MU4 XU22-net16 net20 VSS VSS n w=0.42u l=0.18u
MI2-M_u3 net11 E VDD VDD p w=0.685u l=0.18u
MU24-M_u3 QN net20 VDD VDD p w=1.37u l=0.18u
MU23-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU29-M_u3 net34 net11 VDD VDD p w=0.685u l=0.18u
MU30-M_u3 net20 net15 VDD VDD p w=1.37u l=0.18u
MU32-MU2 net15 net11 XU32-net6 VDD p w=1.12u l=0.18u
MU32-MU1 XU32-net6 D VDD VDD p w=1.12u l=0.18u
MU22-MU2 net15 net34 XU22-net6 VDD p w=0.42u l=0.18u
MU22-MU1 XU22-net6 net20 VDD VDD p w=0.42u l=0.18u
.ends
.subckt LHD2BWP7T D E Q QN VDD VSS 
MI2-M_u2 net11 E VSS VSS n w=0.5u l=0.18u
MU24_0-M_u2 QN net20 VSS VSS n w=1u l=0.18u
MU24_1-M_u2 QN net20 VSS VSS n w=1u l=0.18u
MU23_0-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU23_1-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU29-M_u2 net34 net11 VSS VSS n w=0.5u l=0.18u
MU30-M_u2 net20 net15 VSS VSS n w=1u l=0.18u
MU32-MU3 net15 net34 XU32-net16 VSS n w=0.68u l=0.18u
MU32-MU4 XU32-net16 D VSS VSS n w=0.78u l=0.18u
MU22-MU3 net15 net11 XU22-net16 VSS n w=0.42u l=0.18u
MU22-MU4 XU22-net16 net20 VSS VSS n w=0.42u l=0.18u
MI2-M_u3 net11 E VDD VDD p w=0.685u l=0.18u
MU24_0-M_u3 QN net20 VDD VDD p w=1.37u l=0.18u
MU24_1-M_u3 QN net20 VDD VDD p w=1.37u l=0.18u
MU23_0-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU23_1-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU29-M_u3 net34 net11 VDD VDD p w=0.685u l=0.18u
MU30-M_u3 net20 net15 VDD VDD p w=1.37u l=0.18u
MU32-MU2 net15 net11 XU32-net6 VDD p w=1.12u l=0.18u
MU32-MU1 XU32-net6 D VDD VDD p w=1.12u l=0.18u
MU22-MU2 net15 net34 XU22-net6 VDD p w=0.42u l=0.18u
MU22-MU1 XU22-net6 net20 VDD VDD p w=0.42u l=0.18u
.ends
.subckt LHQD1BWP7T D E Q VDD VSS 
MI2-M_u2 net11 E VSS VSS n w=0.5u l=0.18u
MU23-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU29-M_u2 net34 net11 VSS VSS n w=0.5u l=0.18u
MU30-M_u2 net20 net15 VSS VSS n w=1u l=0.18u
MU32-MU3 net15 net34 XU32-net16 VSS n w=0.68u l=0.18u
MU32-MU4 XU32-net16 D VSS VSS n w=0.78u l=0.18u
MU22-MU3 net15 net11 XU22-net16 VSS n w=0.42u l=0.18u
MU22-MU4 XU22-net16 net20 VSS VSS n w=0.42u l=0.18u
MI2-M_u3 net11 E VDD VDD p w=0.685u l=0.18u
MU23-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU29-M_u3 net34 net11 VDD VDD p w=0.685u l=0.18u
MU30-M_u3 net20 net15 VDD VDD p w=1.37u l=0.18u
MU32-MU2 net15 net11 XU32-net6 VDD p w=1.12u l=0.18u
MU32-MU1 XU32-net6 D VDD VDD p w=1.12u l=0.18u
MU22-MU2 net15 net34 XU22-net6 VDD p w=0.42u l=0.18u
MU22-MU1 XU22-net6 net20 VDD VDD p w=0.42u l=0.18u
.ends
.subckt LHQD2BWP7T D E Q VDD VSS 
MI2-M_u2 net11 E VSS VSS n w=0.5u l=0.18u
MU23_0-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU23_1-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU29-M_u2 net34 net11 VSS VSS n w=0.5u l=0.18u
MU30-M_u2 net20 net15 VSS VSS n w=1u l=0.18u
MU32-MU3 net15 net34 XU32-net16 VSS n w=0.68u l=0.18u
MU32-MU4 XU32-net16 D VSS VSS n w=0.78u l=0.18u
MU22-MU3 net15 net11 XU22-net16 VSS n w=0.42u l=0.18u
MU22-MU4 XU22-net16 net20 VSS VSS n w=0.42u l=0.18u
MI2-M_u3 net11 E VDD VDD p w=0.685u l=0.18u
MU23_0-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU23_1-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU29-M_u3 net34 net11 VDD VDD p w=0.685u l=0.18u
MU30-M_u3 net20 net15 VDD VDD p w=1.37u l=0.18u
MU32-MU2 net15 net11 XU32-net6 VDD p w=1.12u l=0.18u
MU32-MU1 XU32-net6 D VDD VDD p w=1.12u l=0.18u
MU22-MU2 net15 net34 XU22-net6 VDD p w=0.42u l=0.18u
MU22-MU1 XU22-net6 net20 VDD VDD p w=0.42u l=0.18u
.ends
.subckt LHSND1BWP7T D E SDN Q QN VDD VSS 
MI6 net46 net062 net45 VSS n w=0.53u l=0.18u
MI8 net45 D VSS VSS n w=0.53u l=0.18u
MI29 net48 net36 VSS VSS n w=0.53u l=0.18u
MI5 net46 net63 net48 VSS n w=0.53u l=0.18u
M_u2-M_u4 X_u2-net6 net46 VSS VSS n w=0.715u l=0.18u
M_u2-M_u3 net36 SDN X_u2-net6 VSS n w=0.715u l=0.18u
MI4-M_u2 net062 net63 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net61 net36 VSS VSS n w=0.5u l=0.18u
MI12-M_u2 QN net36 VSS VSS n w=1u l=0.18u
MI11-M_u2 Q net61 VSS VSS n w=1u l=0.18u
MI14-M_u2 net63 E VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net36 net46 VDD VDD p w=1u l=0.18u
M_u2-M_u1 net36 SDN VDD VDD p w=1u l=0.18u
MI21 net46 net63 net70 VDD p w=0.42u l=0.18u
MI17 VDD net36 net73 VDD p w=0.42u l=0.18u
MI24 net70 D VDD VDD p w=1.37u l=0.18u
MI18 net46 net062 net73 VDD p w=0.42u l=0.18u
MI4-M_u3 net062 net63 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net61 net36 VDD VDD p w=0.685u l=0.18u
MI12-M_u3 QN net36 VDD VDD p w=1.37u l=0.18u
MI11-M_u3 Q net61 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net63 E VDD VDD p w=0.685u l=0.18u
.ends
.subckt LHSND2BWP7T D E SDN Q QN VDD VSS 
MI6 net46 net062 net45 VSS n w=0.5u l=0.18u
MI8 net45 D VSS VSS n w=0.5u l=0.18u
MI29 net48 net36 VSS VSS n w=0.42u l=0.18u
MI5 net46 net63 net48 VSS n w=0.42u l=0.18u
M_u2-M_u4 X_u2-net6 net46 VSS VSS n w=0.685u l=0.18u
M_u2-M_u3 net36 SDN X_u2-net6 VSS n w=0.685u l=0.18u
MI4-M_u2 net062 net63 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net64 net36 VSS VSS n w=1u l=0.18u
MI12_0-M_u2 QN net36 VSS VSS n w=1u l=0.18u
MI12_1-M_u2 QN net36 VSS VSS n w=1u l=0.18u
MI11_0-M_u2 Q net64 VSS VSS n w=1u l=0.18u
MI11_1-M_u2 Q net64 VSS VSS n w=1u l=0.18u
MI14-M_u2 net63 E VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net36 net46 VDD VDD p w=0.975u l=0.18u
M_u2-M_u1 net36 SDN VDD VDD p w=0.975u l=0.18u
MI21 net46 net63 net70 VDD p w=0.42u l=0.18u
MI17 VDD net36 net73 VDD p w=0.42u l=0.18u
MI24 net70 D VDD VDD p w=1.345u l=0.18u
MI18 net46 net062 net73 VDD p w=0.42u l=0.18u
MI4-M_u3 net062 net63 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net64 net36 VDD VDD p w=1.37u l=0.18u
MI12_0-M_u3 QN net36 VDD VDD p w=1.37u l=0.18u
MI12_1-M_u3 QN net36 VDD VDD p w=1.37u l=0.18u
MI11_0-M_u3 Q net64 VDD VDD p w=1.37u l=0.18u
MI11_1-M_u3 Q net64 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net63 E VDD VDD p w=0.685u l=0.18u
.ends
.subckt LHSNQD1BWP7T D E SDN Q VDD VSS 
MI6 net46 net060 net45 VSS n w=0.5u l=0.18u
MI8 net45 D VSS VSS n w=0.5u l=0.18u
MI29 net48 net36 VSS VSS n w=0.42u l=0.18u
MI5 net46 net63 net48 VSS n w=0.42u l=0.18u
M_u2-M_u4 X_u2-net6 net46 VSS VSS n w=0.685u l=0.18u
M_u2-M_u3 net36 SDN X_u2-net6 VSS n w=0.685u l=0.18u
MI4-M_u2 net060 net63 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net61 net36 VSS VSS n w=0.5u l=0.18u
MI11-M_u2 Q net61 VSS VSS n w=1u l=0.18u
MI14-M_u2 net63 E VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net36 net46 VDD VDD p w=1u l=0.18u
M_u2-M_u1 net36 SDN VDD VDD p w=1u l=0.18u
MI21 net46 net63 net70 VDD p w=0.42u l=0.18u
MI17 VDD net36 net73 VDD p w=0.42u l=0.18u
MI24 net70 D VDD VDD p w=1u l=0.18u
MI18 net46 net060 net73 VDD p w=0.42u l=0.18u
MI4-M_u3 net060 net63 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net61 net36 VDD VDD p w=0.88u l=0.18u
MI11-M_u3 Q net61 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net63 E VDD VDD p w=0.685u l=0.18u
.ends
.subckt LHSNQD2BWP7T D E SDN Q VDD VSS 
MI6 net46 net062 net45 VSS n w=0.5u l=0.18u
MI8 net45 D VSS VSS n w=0.5u l=0.18u
MI29 net48 net36 VSS VSS n w=0.42u l=0.18u
MI5 net46 net63 net48 VSS n w=0.42u l=0.18u
M_u2-M_u4 X_u2-net6 net46 VSS VSS n w=0.685u l=0.18u
M_u2-M_u3 net36 SDN X_u2-net6 VSS n w=0.685u l=0.18u
MI4-M_u2 net062 net63 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net64 net36 VSS VSS n w=1u l=0.18u
MI11_0-M_u2 Q net64 VSS VSS n w=1u l=0.18u
MI11_1-M_u2 Q net64 VSS VSS n w=1u l=0.18u
MI14-M_u2 net63 E VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net36 net46 VDD VDD p w=0.975u l=0.18u
M_u2-M_u1 net36 SDN VDD VDD p w=0.975u l=0.18u
MI21 net46 net63 net70 VDD p w=0.7u l=0.18u
MI17 VDD net36 net73 VDD p w=0.42u l=0.18u
MI24 net70 D VDD VDD p w=1u l=0.18u
MI18 net46 net062 net73 VDD p w=0.42u l=0.18u
MI4-M_u3 net062 net63 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net64 net36 VDD VDD p w=1.37u l=0.18u
MI11_0-M_u3 Q net64 VDD VDD p w=1.37u l=0.18u
MI11_1-M_u3 Q net64 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net63 E VDD VDD p w=0.685u l=0.18u
.ends
.subckt LNCND1BWP7T D EN CDN Q QN VDD VSS 
MI29 net45 net169 net40 VSS n w=0.42u l=0.18u
MI5 net166 net069 net45 VSS n w=0.42u l=0.18u
MI6 net166 net167 net171 VSS n w=0.57u l=0.18u
MI8 net171 D net51 VSS n w=0.57u l=0.18u
MI9 net51 CDN VSS VSS n w=0.815u l=0.18u
MI10 net40 CDN VSS VSS n w=0.42u l=0.18u
MI33-M_u2 net069 net167 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net170 net169 VSS VSS n w=1u l=0.18u
MI11-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI12-M_u2 QN net169 VSS VSS n w=1u l=0.18u
MI14-M_u2 net167 EN VSS VSS n w=0.5u l=0.18u
MI32-M_u2 net169 net166 VSS VSS n w=1u l=0.18u
MI30 net166 CDN VDD VDD p w=0.685u l=0.18u
MI17 VDD net169 net106 VDD p w=0.42u l=0.18u
MI18 net166 net167 net106 VDD p w=0.42u l=0.18u
MI21 net166 net069 net110 VDD p w=1.12u l=0.18u
MI24 net110 D VDD VDD p w=1.12u l=0.18u
MI33-M_u3 net069 net167 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net170 net169 VDD VDD p w=1.37u l=0.18u
MI11-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI12-M_u3 QN net169 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net167 EN VDD VDD p w=0.685u l=0.18u
MI32-M_u3 net169 net166 VDD VDD p w=1.37u l=0.18u
.ends
.subckt LNCND2BWP7T D EN CDN Q QN VDD VSS 
MI29 net45 net169 net40 VSS n w=0.42u l=0.18u
MI5 net166 net069 net45 VSS n w=0.42u l=0.18u
MI6 net166 net167 net171 VSS n w=0.57u l=0.18u
MI8 net171 D net51 VSS n w=0.57u l=0.18u
MI9 net51 CDN VSS VSS n w=0.815u l=0.18u
MI10 net40 CDN VSS VSS n w=0.42u l=0.18u
MI33-M_u2 net069 net167 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net170 net169 VSS VSS n w=1u l=0.18u
MI11_0-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI11_1-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI12_0-M_u2 QN net169 VSS VSS n w=1u l=0.18u
MI12_1-M_u2 QN net169 VSS VSS n w=1u l=0.18u
MI14-M_u2 net167 EN VSS VSS n w=0.5u l=0.18u
MI32-M_u2 net169 net166 VSS VSS n w=1u l=0.18u
MI30 net166 CDN VDD VDD p w=0.685u l=0.18u
MI17 VDD net169 net106 VDD p w=0.42u l=0.18u
MI18 net166 net167 net106 VDD p w=0.42u l=0.18u
MI21 net166 net069 net110 VDD p w=1.12u l=0.18u
MI24 net110 D VDD VDD p w=1.12u l=0.18u
MI33-M_u3 net069 net167 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net170 net169 VDD VDD p w=1.37u l=0.18u
MI11_0-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI11_1-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI12_0-M_u3 QN net169 VDD VDD p w=1.37u l=0.18u
MI12_1-M_u3 QN net169 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net167 EN VDD VDD p w=0.685u l=0.18u
MI32-M_u3 net169 net166 VDD VDD p w=1.37u l=0.18u
.ends
.subckt LNCNQD1BWP7T D EN CDN Q VDD VSS 
MI29 net45 net169 net40 VSS n w=0.42u l=0.18u
MI5 net166 net069 net45 VSS n w=0.42u l=0.18u
MI6 net166 net167 net171 VSS n w=0.57u l=0.18u
MI8 net171 D net51 VSS n w=0.57u l=0.18u
MI9 net51 CDN VSS VSS n w=0.815u l=0.18u
MI10 net40 CDN VSS VSS n w=0.42u l=0.18u
MI33-M_u2 net069 net167 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net170 net169 VSS VSS n w=1u l=0.18u
MI11-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI14-M_u2 net167 EN VSS VSS n w=0.5u l=0.18u
MI32-M_u2 net169 net166 VSS VSS n w=1u l=0.18u
MI30 net166 CDN VDD VDD p w=0.685u l=0.18u
MI17 VDD net169 net106 VDD p w=0.42u l=0.18u
MI18 net166 net167 net106 VDD p w=0.42u l=0.18u
MI21 net166 net069 net110 VDD p w=1.12u l=0.18u
MI24 net110 D VDD VDD p w=1.12u l=0.18u
MI33-M_u3 net069 net167 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net170 net169 VDD VDD p w=1.37u l=0.18u
MI11-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net167 EN VDD VDD p w=0.685u l=0.18u
MI32-M_u3 net169 net166 VDD VDD p w=1.37u l=0.18u
.ends
.subckt LNCNQD2BWP7T D EN CDN Q VDD VSS 
MI29 net45 net169 net40 VSS n w=0.42u l=0.18u
MI5 net166 net069 net45 VSS n w=0.42u l=0.18u
MI6 net166 net167 net171 VSS n w=0.57u l=0.18u
MI8 net171 D net51 VSS n w=0.57u l=0.18u
MI9 net51 CDN VSS VSS n w=0.815u l=0.18u
MI10 net40 CDN VSS VSS n w=0.42u l=0.18u
MI33-M_u2 net069 net167 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net170 net169 VSS VSS n w=1u l=0.18u
MI11_0-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI11_1-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI14-M_u2 net167 EN VSS VSS n w=0.5u l=0.18u
MI32-M_u2 net169 net166 VSS VSS n w=1u l=0.18u
MI30 net166 CDN VDD VDD p w=0.685u l=0.18u
MI17 VDD net169 net106 VDD p w=0.42u l=0.18u
MI18 net166 net167 net106 VDD p w=0.42u l=0.18u
MI21 net166 net069 net110 VDD p w=1.12u l=0.18u
MI24 net110 D VDD VDD p w=1.12u l=0.18u
MI33-M_u3 net069 net167 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net170 net169 VDD VDD p w=1.37u l=0.18u
MI11_0-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI11_1-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net167 EN VDD VDD p w=0.685u l=0.18u
MI32-M_u3 net169 net166 VDD VDD p w=1.37u l=0.18u
.ends
.subckt LND1BWP7T D EN Q QN VDD VSS 
MI2-M_u2 net9 EN VSS VSS n w=0.5u l=0.18u
MU23-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU24-M_u2 QN net20 VSS VSS n w=1u l=0.18u
MU29-M_u2 net30 net9 VSS VSS n w=0.5u l=0.18u
MU30-M_u2 net20 net15 VSS VSS n w=1u l=0.18u
MU32-MU3 net15 net9 XU32-net16 VSS n w=0.68u l=0.18u
MU32-MU4 XU32-net16 D VSS VSS n w=0.78u l=0.18u
MU22-MU3 net15 net30 XU22-net16 VSS n w=0.42u l=0.18u
MU22-MU4 XU22-net16 net20 VSS VSS n w=0.42u l=0.18u
MI2-M_u3 net9 EN VDD VDD p w=0.685u l=0.18u
MU23-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU24-M_u3 QN net20 VDD VDD p w=1.37u l=0.18u
MU29-M_u3 net30 net9 VDD VDD p w=0.685u l=0.18u
MU30-M_u3 net20 net15 VDD VDD p w=1.37u l=0.18u
MU32-MU2 net15 net30 XU32-net6 VDD p w=1.12u l=0.18u
MU32-MU1 XU32-net6 D VDD VDD p w=1.12u l=0.18u
MU22-MU2 net15 net9 XU22-net6 VDD p w=0.42u l=0.18u
MU22-MU1 XU22-net6 net20 VDD VDD p w=0.42u l=0.18u
.ends
.subckt LND2BWP7T D EN Q QN VDD VSS 
MI2-M_u2 net9 EN VSS VSS n w=0.5u l=0.18u
MU23_0-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU23_1-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU24_0-M_u2 QN net20 VSS VSS n w=1u l=0.18u
MU24_1-M_u2 QN net20 VSS VSS n w=1u l=0.18u
MU29-M_u2 net30 net9 VSS VSS n w=0.5u l=0.18u
MU30-M_u2 net20 net15 VSS VSS n w=1u l=0.18u
MU32-MU3 net15 net9 XU32-net16 VSS n w=0.68u l=0.18u
MU32-MU4 XU32-net16 D VSS VSS n w=0.78u l=0.18u
MU22-MU3 net15 net30 XU22-net16 VSS n w=0.42u l=0.18u
MU22-MU4 XU22-net16 net20 VSS VSS n w=0.42u l=0.18u
MI2-M_u3 net9 EN VDD VDD p w=0.685u l=0.18u
MU23_0-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU23_1-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU24_0-M_u3 QN net20 VDD VDD p w=1.37u l=0.18u
MU24_1-M_u3 QN net20 VDD VDD p w=1.37u l=0.18u
MU29-M_u3 net30 net9 VDD VDD p w=0.685u l=0.18u
MU30-M_u3 net20 net15 VDD VDD p w=1.37u l=0.18u
MU32-MU2 net15 net30 XU32-net6 VDD p w=1.12u l=0.18u
MU32-MU1 XU32-net6 D VDD VDD p w=1.12u l=0.18u
MU22-MU2 net15 net9 XU22-net6 VDD p w=0.42u l=0.18u
MU22-MU1 XU22-net6 net20 VDD VDD p w=0.42u l=0.18u
.ends
.subckt LNQD1BWP7T D EN Q VDD VSS 
MI2-M_u2 net9 EN VSS VSS n w=0.5u l=0.18u
MU23-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU29-M_u2 net30 net9 VSS VSS n w=0.5u l=0.18u
MU30-M_u2 net20 net15 VSS VSS n w=1u l=0.18u
MU32-MU3 net15 net9 XU32-net16 VSS n w=0.68u l=0.18u
MU32-MU4 XU32-net16 D VSS VSS n w=0.78u l=0.18u
MU22-MU3 net15 net30 XU22-net16 VSS n w=0.42u l=0.18u
MU22-MU4 XU22-net16 net20 VSS VSS n w=0.42u l=0.18u
MI2-M_u3 net9 EN VDD VDD p w=0.685u l=0.18u
MU23-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU29-M_u3 net30 net9 VDD VDD p w=0.685u l=0.18u
MU30-M_u3 net20 net15 VDD VDD p w=1.37u l=0.18u
MU32-MU2 net15 net30 XU32-net6 VDD p w=1.12u l=0.18u
MU32-MU1 XU32-net6 D VDD VDD p w=1.12u l=0.18u
MU22-MU2 net15 net9 XU22-net6 VDD p w=0.42u l=0.18u
MU22-MU1 XU22-net6 net20 VDD VDD p w=0.42u l=0.18u
.ends
.subckt LNQD2BWP7T D EN Q VDD VSS 
MI2-M_u2 net9 EN VSS VSS n w=0.5u l=0.18u
MU23_0-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU23_1-M_u2 Q net15 VSS VSS n w=1u l=0.18u
MU29-M_u2 net30 net9 VSS VSS n w=0.5u l=0.18u
MU30-M_u2 net20 net15 VSS VSS n w=1u l=0.18u
MU32-MU3 net15 net9 XU32-net16 VSS n w=0.68u l=0.18u
MU32-MU4 XU32-net16 D VSS VSS n w=0.78u l=0.18u
MU22-MU3 net15 net30 XU22-net16 VSS n w=0.42u l=0.18u
MU22-MU4 XU22-net16 net20 VSS VSS n w=0.42u l=0.18u
MI2-M_u3 net9 EN VDD VDD p w=0.685u l=0.18u
MU23_0-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU23_1-M_u3 Q net15 VDD VDD p w=1.37u l=0.18u
MU29-M_u3 net30 net9 VDD VDD p w=0.685u l=0.18u
MU30-M_u3 net20 net15 VDD VDD p w=1.37u l=0.18u
MU32-MU2 net15 net30 XU32-net6 VDD p w=1.12u l=0.18u
MU32-MU1 XU32-net6 D VDD VDD p w=1.12u l=0.18u
MU22-MU2 net15 net9 XU22-net6 VDD p w=0.42u l=0.18u
MU22-MU1 XU22-net6 net20 VDD VDD p w=0.42u l=0.18u
.ends
.subckt LNSND1BWP7T D EN SDN Q QN VDD VSS 
MI29 net45 net169 VSS VSS n w=0.5u l=0.18u
MI5 net166 net056 net45 VSS n w=0.5u l=0.18u
MI6 net166 net167 net171 VSS n w=0.5u l=0.18u
MI8 net171 D VSS VSS n w=0.5u l=0.18u
M_u2-M_u4 X_u2-net6 net166 VSS VSS n w=0.685u l=0.18u
M_u2-M_u3 net169 SDN X_u2-net6 VSS n w=0.685u l=0.18u
MI32-M_u2 net056 net167 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net170 net169 VSS VSS n w=0.5u l=0.18u
MI11-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI12-M_u2 QN net169 VSS VSS n w=1u l=0.18u
MI14-M_u2 net167 EN VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net169 net166 VDD VDD p w=1u l=0.18u
M_u2-M_u1 net169 SDN VDD VDD p w=1u l=0.18u
MI17 VDD net169 net106 VDD p w=0.42u l=0.18u
MI18 net166 net167 net106 VDD p w=0.42u l=0.18u
MI21 net166 net056 net110 VDD p w=0.42u l=0.18u
MI24 net110 D VDD VDD p w=1u l=0.18u
MI32-M_u3 net056 net167 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net170 net169 VDD VDD p w=0.685u l=0.18u
MI11-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI12-M_u3 QN net169 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net167 EN VDD VDD p w=0.685u l=0.18u
.ends
.subckt LNSND2BWP7T D EN SDN Q QN VDD VSS 
MI29 net45 net169 VSS VSS n w=0.5u l=0.18u
MI5 net166 net056 net45 VSS n w=0.5u l=0.18u
MI6 net166 net167 net171 VSS n w=0.5u l=0.18u
MI8 net171 D VSS VSS n w=0.5u l=0.18u
M_u2-M_u4 X_u2-net6 net166 VSS VSS n w=0.685u l=0.18u
M_u2-M_u3 net169 SDN X_u2-net6 VSS n w=0.685u l=0.18u
MI32-M_u2 net056 net167 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net170 net169 VSS VSS n w=1u l=0.18u
MI11_0-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI11_1-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI12_0-M_u2 QN net169 VSS VSS n w=1u l=0.18u
MI12_1-M_u2 QN net169 VSS VSS n w=1u l=0.18u
MI14-M_u2 net167 EN VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net169 net166 VDD VDD p w=0.975u l=0.18u
M_u2-M_u1 net169 SDN VDD VDD p w=0.975u l=0.18u
MI17 VDD net169 net106 VDD p w=0.42u l=0.18u
MI18 net166 net167 net106 VDD p w=0.42u l=0.18u
MI21 net166 net056 net110 VDD p w=0.42u l=0.18u
MI24 net110 D VDD VDD p w=1u l=0.18u
MI32-M_u3 net056 net167 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net170 net169 VDD VDD p w=1.37u l=0.18u
MI11_0-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI11_1-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI12_0-M_u3 QN net169 VDD VDD p w=1.37u l=0.18u
MI12_1-M_u3 QN net169 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net167 EN VDD VDD p w=0.685u l=0.18u
.ends
.subckt LNSNQD1BWP7T D EN SDN Q VDD VSS 
MI29 net45 net169 VSS VSS n w=0.42u l=0.18u
MI5 net166 net054 net45 VSS n w=0.42u l=0.18u
MI6 net166 net167 net171 VSS n w=0.5u l=0.18u
MI8 net171 D VSS VSS n w=0.5u l=0.18u
M_u2-M_u4 X_u2-net6 net166 VSS VSS n w=0.685u l=0.18u
M_u2-M_u3 net169 SDN X_u2-net6 VSS n w=0.685u l=0.18u
MI32-M_u2 net054 net167 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net170 net169 VSS VSS n w=0.5u l=0.18u
MI11-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI14-M_u2 net167 EN VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net169 net166 VDD VDD p w=1u l=0.18u
M_u2-M_u1 net169 SDN VDD VDD p w=1u l=0.18u
MI17 VDD net169 net106 VDD p w=0.42u l=0.18u
MI18 net166 net167 net106 VDD p w=0.42u l=0.18u
MI21 net166 net054 net110 VDD p w=0.42u l=0.18u
MI24 net110 D VDD VDD p w=1u l=0.18u
MI32-M_u3 net054 net167 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net170 net169 VDD VDD p w=0.685u l=0.18u
MI11-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net167 EN VDD VDD p w=0.685u l=0.18u
.ends
.subckt LNSNQD2BWP7T D EN SDN Q VDD VSS 
MI29 net45 net169 VSS VSS n w=0.5u l=0.18u
MI5 net166 net059 net45 VSS n w=0.5u l=0.18u
MI6 net166 net167 net171 VSS n w=0.5u l=0.18u
MI8 net171 D VSS VSS n w=0.5u l=0.18u
M_u2-M_u4 X_u2-net6 net166 VSS VSS n w=0.685u l=0.18u
M_u2-M_u3 net169 SDN X_u2-net6 VSS n w=0.685u l=0.18u
MI32-M_u2 net059 net167 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net170 net169 VSS VSS n w=1u l=0.18u
MI11_0-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI11_1-M_u2 Q net170 VSS VSS n w=1u l=0.18u
MI14-M_u2 net167 EN VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net169 net166 VDD VDD p w=0.975u l=0.18u
M_u2-M_u1 net169 SDN VDD VDD p w=0.975u l=0.18u
MI17 VDD net169 net106 VDD p w=0.42u l=0.18u
MI18 net166 net167 net106 VDD p w=0.42u l=0.18u
MI21 net166 net059 net110 VDD p w=0.42u l=0.18u
MI24 net110 D VDD VDD p w=1u l=0.18u
MI32-M_u3 net059 net167 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net170 net169 VDD VDD p w=1.37u l=0.18u
MI11_0-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI11_1-M_u3 Q net170 VDD VDD p w=1.37u l=0.18u
MI14-M_u3 net167 EN VDD VDD p w=0.685u l=0.18u
.ends
.subckt MAOI222D0BWP7T A B C ZN VDD VSS 
MU10 net26 C VSS VSS n w=0.5u l=0.18u
MU9 net26 A ZN VSS n w=0.5u l=0.18u
MU8 net26 B ZN VSS n w=0.5u l=0.18u
MU6 ZN A net38 VSS n w=0.5u l=0.18u
MU7 net38 B VSS VSS n w=0.5u l=0.18u
MU2 net16 B VDD VDD p w=0.685u l=0.18u
MU5 net20 A ZN VDD p w=0.685u l=0.18u
MU3 ZN A net16 VDD p w=0.685u l=0.18u
MU4 net20 B ZN VDD p w=0.685u l=0.18u
MU1 net20 C VDD VDD p w=0.685u l=0.18u
.ends
.subckt MAOI222D1BWP7T A B C ZN VDD VSS 
MU10 net26 C VSS VSS n w=1u l=0.18u
MU9 net26 A ZN VSS n w=1u l=0.18u
MI1 net26 B ZN VSS n w=1u l=0.18u
MU6 ZN A net38 VSS n w=1u l=0.18u
MU7 net38 B VSS VSS n w=1u l=0.18u
MU2 net16 B VDD VDD p w=1.37u l=0.18u
MU5 net20 A ZN VDD p w=1.37u l=0.18u
MU3 ZN A net16 VDD p w=1.37u l=0.18u
MU4 net20 B ZN VDD p w=1.37u l=0.18u
MU1 net20 C VDD VDD p w=1.37u l=0.18u
.ends
.subckt MAOI222D2BWP7T A B C ZN VDD VSS 
MU10 net26 C VSS VSS n w=1u l=0.18u
MU9 net26 A net31 VSS n w=1u l=0.18u
MU8 net26 B net31 VSS n w=1u l=0.18u
MU6 net31 A net38 VSS n w=1u l=0.18u
MU7 net38 B VSS VSS n w=1u l=0.18u
MU20_0-M_u2 ZN net58 VSS VSS n w=1u l=0.18u
MU20_1-M_u2 ZN net58 VSS VSS n w=1u l=0.18u
MU19-M_u2 net58 net31 VSS VSS n w=1u l=0.18u
MU20_0-M_u3 ZN net58 VDD VDD p w=1.37u l=0.18u
MU20_1-M_u3 ZN net58 VDD VDD p w=1.37u l=0.18u
MU19-M_u3 net58 net31 VDD VDD p w=1.37u l=0.18u
MU2 net16 B VDD VDD p w=1.37u l=0.18u
MU5 net20 A net31 VDD p w=1.37u l=0.18u
MU3 net31 A net16 VDD p w=1.37u l=0.18u
MU4 net20 B net31 VDD p w=1.37u l=0.18u
MU1 net20 C VDD VDD p w=1.37u l=0.18u
.ends
.subckt MAOI22D0BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI11 net17 B2 VSS VSS n w=0.5u l=0.18u
MI12 net17 B1 VSS VSS n w=0.5u l=0.18u
MI9 net63 A2 VSS VSS n w=0.5u l=0.18u
MI10 ZN net17 VSS VSS n w=0.5u l=0.18u
MI3 ZN A1 net63 VSS n w=0.5u l=0.18u
MI6 ZN A2 net31 VDD p w=0.685u l=0.18u
MI1 net39 B2 VDD VDD p w=0.685u l=0.18u
MI5 net17 B1 net39 VDD p w=0.685u l=0.18u
MI13 net31 net17 VDD VDD p w=0.685u l=0.18u
MI7 ZN A1 net31 VDD p w=0.685u l=0.18u
.ends
.subckt MAOI22D1BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI11 net17 B2 VSS VSS n w=1u l=0.18u
MI12 net17 B1 VSS VSS n w=1u l=0.18u
MI9 net63 A2 VSS VSS n w=1u l=0.18u
MI10 ZN net17 VSS VSS n w=1u l=0.18u
MI3 ZN A1 net63 VSS n w=1u l=0.18u
MI6 ZN A2 net31 VDD p w=1.37u l=0.18u
MI1 net39 B2 VDD VDD p w=1.37u l=0.18u
MI5 net17 B1 net39 VDD p w=1.37u l=0.18u
MI13 net31 net17 VDD VDD p w=1.37u l=0.18u
MI7 ZN A1 net31 VDD p w=1.37u l=0.18u
.ends
.subckt MAOI22D2BWP7T A1 A2 B1 B2 ZN VDD VSS 
MU16_0-M_u2 ZN net25 VSS VSS n w=1u l=0.18u
MU16_1-M_u2 ZN net25 VSS VSS n w=1u l=0.18u
MI1 net37 A1 net67 VSS n w=1u l=0.18u
MI2 net67 A2 VSS VSS n w=1u l=0.18u
MU10 net22 B2 net25 VSS n w=1u l=0.18u
MU9 net22 B1 net25 VSS n w=1u l=0.18u
MU8 net22 net37 VSS VSS n w=1u l=0.18u
MU16_0-M_u3 ZN net25 VDD VDD p w=1.37u l=0.18u
MU16_1-M_u3 ZN net25 VDD VDD p w=1.37u l=0.18u
MI5 net50 B1 net25 VDD p w=1.37u l=0.18u
MI4 VDD B2 net50 VDD p w=1.37u l=0.18u
MU5 net25 net37 VDD VDD p w=1.37u l=0.18u
MU4 net37 A1 VDD VDD p w=1.37u l=0.18u
MU3 net37 A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt MOAI22D0BWP7T A1 A2 B1 B2 ZN VDD VSS 
MU1 net8 B1 net26 VSS n w=0.5u l=0.18u
MI5 net26 B2 VSS VSS n w=0.5u l=0.18u
MI6 net29 net8 VSS VSS n w=0.5u l=0.18u
MU9 net29 A1 ZN VSS n w=0.5u l=0.18u
MU10 net29 A2 ZN VSS n w=0.5u l=0.18u
MU3 net8 B2 VDD VDD p w=0.685u l=0.18u
MI1 net8 B1 VDD VDD p w=0.685u l=0.18u
MI2 ZN net8 VDD VDD p w=0.685u l=0.18u
MI4 ZN A1 net20 VDD p w=0.685u l=0.18u
MI3 net20 A2 VDD VDD p w=0.685u l=0.18u
.ends
.subckt MOAI22D1BWP7T A1 A2 B1 B2 ZN VDD VSS 
MU1 net8 B1 net26 VSS n w=1u l=0.18u
MI5 net26 B2 VSS VSS n w=1u l=0.18u
MI6 net29 net8 VSS VSS n w=1u l=0.18u
MU9 net29 A1 ZN VSS n w=1u l=0.18u
MU10 net29 A2 ZN VSS n w=1u l=0.18u
MU3 net8 B2 VDD VDD p w=1.37u l=0.18u
MI1 net8 B1 VDD VDD p w=1.37u l=0.18u
MI2 ZN net8 VDD VDD p w=1.37u l=0.18u
MI4 ZN A1 net20 VDD p w=1.37u l=0.18u
MI3 net20 A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt MOAI22D2BWP7T A1 A2 B1 B2 ZN VDD VSS 
MU18_0-M_u2 ZN net22 VSS VSS n w=1u l=0.18u
MU18_1-M_u2 ZN net22 VSS VSS n w=1u l=0.18u
MU6 net22 B1 net13 VSS n w=1u l=0.18u
MU7 net13 B2 VSS VSS n w=1u l=0.18u
MU8 net16 A1 VSS VSS n w=1u l=0.18u
MU9 net16 A2 VSS VSS n w=1u l=0.18u
MU5 net22 net16 VSS VSS n w=1u l=0.18u
MU18_0-M_u3 ZN net22 VDD VDD p w=1.37u l=0.18u
MU18_1-M_u3 ZN net22 VDD VDD p w=1.37u l=0.18u
MU4 net22 B1 net31 VDD p w=1.37u l=0.18u
MU1 net31 net16 VDD VDD p w=1.37u l=0.18u
MU2 net31 B2 net22 VDD p w=1.37u l=0.18u
MU10 net36 A1 VDD VDD p w=1.37u l=0.18u
MU11 net16 A2 net36 VDD p w=1.37u l=0.18u
.ends
.subckt MUX2D0BWP7T I0 I1 S Z VDD VSS 
MI15-M_u2 net6 S VSS VSS n w=0.5u l=0.18u
MU29-M_u2 Z net28 VSS VSS n w=0.5u l=0.18u
MI19 net026 I0 VSS VSS n w=0.5u l=0.18u
MI20 net023 I1 VSS VSS n w=0.5u l=0.18u
MI12 net28 net6 net026 VSS n w=0.5u l=0.18u
MI21 net28 S net023 VSS n w=0.5u l=0.18u
MI15-M_u3 net6 S VDD VDD p w=0.685u l=0.18u
MU29-M_u3 Z net28 VDD VDD p w=0.685u l=0.18u
MI111 net042 I0 VDD VDD p w=0.685u l=0.18u
MI5 net28 S net042 VDD p w=0.685u l=0.18u
MI25 net28 net6 net033 VDD p w=0.685u l=0.18u
MI24 net033 I1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt MUX2D1BWP7T I0 I1 S Z VDD VSS 
MI15-M_u2 net6 S VSS VSS n w=0.5u l=0.18u
MU29-M_u2 Z net28 VSS VSS n w=1u l=0.18u
M_u2 net026 I0 VSS VSS n w=1u l=0.18u
MI17 net28 net6 net026 VSS n w=0.5u l=0.18u
MI23 net056 I1 VSS VSS n w=1u l=0.18u
MI24 net28 S net056 VSS n w=0.5u l=0.18u
MI15-M_u3 net6 S VDD VDD p w=0.685u l=0.18u
MU29-M_u3 Z net28 VDD VDD p w=1.37u l=0.18u
MI21 net28 net6 net045 VDD p w=0.685u l=0.18u
M_u1 net021 I0 VDD VDD p w=0.94u l=0.18u
MI16 net28 S net021 VDD p w=0.685u l=0.18u
MI22 net045 I1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt MUX2D2BWP7T I0 I1 S Z VDD VSS 
MI15-M_u2 net043 S VSS VSS n w=0.5u l=0.18u
MU29_0-M_u2 Z net026 VSS VSS n w=1u l=0.18u
MU29_1-M_u2 Z net026 VSS VSS n w=1u l=0.18u
MI23 net023 I1 VSS VSS n w=1u l=0.18u
MI24 net026 S net023 VSS n w=0.5u l=0.18u
MI17 net026 net043 net029 VSS n w=0.5u l=0.18u
M_u2 net029 I0 VSS VSS n w=1u l=0.18u
MI15-M_u3 net043 S VDD VDD p w=0.685u l=0.18u
MU29_0-M_u3 Z net026 VDD VDD p w=1.37u l=0.18u
MU29_1-M_u3 Z net026 VDD VDD p w=1.37u l=0.18u
MI21 net026 net043 net042 VDD p w=0.685u l=0.18u
M_u1 net036 I0 VDD VDD p w=0.94u l=0.18u
MI22 net042 I1 VDD VDD p w=1.37u l=0.18u
MI16 net026 S net036 VDD p w=0.685u l=0.18u
.ends
.subckt MUX2ND0BWP7T I0 I1 S ZN VDD VSS 
MI15-M_u2 net19 S VSS VSS n w=0.5u l=0.18u
MI21 ZN S net40 VSS n w=0.5u l=0.18u
MI12 ZN net19 net36 VSS n w=0.5u l=0.18u
MI20 net40 I1 VSS VSS n w=1u l=0.18u
MI19 net36 I0 VSS VSS n w=1u l=0.18u
MI15-M_u3 net19 S VDD VDD p w=0.685u l=0.18u
MI25 ZN net19 net26 VDD p w=0.685u l=0.18u
MI24 net26 I1 VDD VDD p w=1.37u l=0.18u
MI5 ZN S net30 VDD p w=0.685u l=0.18u
MI111 net30 I0 VDD VDD p w=0.94u l=0.18u
.ends
.subckt MUX2ND1BWP7T I0 I1 S ZN VDD VSS 
MI15-M_u2 net045 S VSS VSS n w=0.5u l=0.18u
MI16-M_u2 net48 net28 VSS VSS n w=0.5u l=0.18u
MU29-M_u2 ZN net48 VSS VSS n w=1u l=0.18u
MI25 net28 S net025 VSS n w=0.5u l=0.18u
M_u2 net031 I0 VSS VSS n w=1u l=0.18u
MI24 net025 I1 VSS VSS n w=1u l=0.18u
MI23 net28 net045 net031 VSS n w=0.5u l=0.18u
MI15-M_u3 net045 S VDD VDD p w=0.685u l=0.18u
MI16-M_u3 net48 net28 VDD VDD p w=0.685u l=0.18u
MU29-M_u3 ZN net48 VDD VDD p w=1.37u l=0.18u
M_u1 net038 I0 VDD VDD p w=0.94u l=0.18u
MI17 net28 S net038 VDD p w=0.685u l=0.18u
MI22 net044 I1 VDD VDD p w=1.37u l=0.18u
MI21 net28 net045 net044 VDD p w=0.685u l=0.18u
.ends
.subckt MUX2ND2BWP7T I0 I1 S ZN VDD VSS 
MI15-M_u2 net045 S VSS VSS n w=0.5u l=0.18u
MI16-M_u2 net27 net28 VSS VSS n w=1u l=0.18u
MU29_0-M_u2 ZN net27 VSS VSS n w=1u l=0.18u
MU29_1-M_u2 ZN net27 VSS VSS n w=1u l=0.18u
MI25 net28 S net025 VSS n w=0.5u l=0.18u
M_u2 net031 I0 VSS VSS n w=1u l=0.18u
MI24 net025 I1 VSS VSS n w=1u l=0.18u
MI17 net28 net045 net031 VSS n w=0.5u l=0.18u
MI15-M_u3 net045 S VDD VDD p w=0.685u l=0.18u
MI16-M_u3 net27 net28 VDD VDD p w=1.37u l=0.18u
MU29_0-M_u3 ZN net27 VDD VDD p w=1.37u l=0.18u
MU29_1-M_u3 ZN net27 VDD VDD p w=1.37u l=0.18u
M_u1 net038 I0 VDD VDD p w=0.94u l=0.18u
MI22 net28 S net038 VDD p w=0.685u l=0.18u
MI23 net044 I1 VDD VDD p w=1.37u l=0.18u
MI21 net28 net045 net044 VDD p w=0.685u l=0.18u
.ends
.subckt MUX3D0BWP7T I0 I1 I2 S0 S1 Z VDD VSS 
MI41 net75 I0 VSS VSS n w=0.5u l=0.18u
MI42 net72 I1 VSS VSS n w=0.5u l=0.18u
MI43 PG1 net88 net75 VSS n w=0.5u l=0.18u
MI44 PG1 S0 net72 VSS n w=0.5u l=0.18u
MI45 net70 I2 VSS VSS n w=0.5u l=0.18u
MI46 OUT S1 net70 VSS n w=0.5u l=0.18u
MI50-M_u2 net88 S0 VSS VSS n w=0.5u l=0.18u
MI51-M_u2 Z OUT VSS VSS n w=0.5u l=0.18u
MI52-M_u2 net84 S1 VSS VSS n w=0.5u l=0.18u
MI53-M_u2 PG1 net84 OUT VSS n w=0.5u l=0.18u
MI35 net62 I0 VDD VDD p w=0.685u l=0.18u
MI36 PG1 S0 net62 VDD p w=0.685u l=0.18u
MI37 PG1 net88 net54 VDD p w=0.685u l=0.18u
MI38 net54 I1 VDD VDD p w=0.685u l=0.18u
MI39 net50 I2 VDD VDD p w=0.685u l=0.18u
MI40 OUT net84 net50 VDD p w=0.685u l=0.18u
MI50-M_u3 net88 S0 VDD VDD p w=0.685u l=0.18u
MI51-M_u3 Z OUT VDD VDD p w=0.685u l=0.18u
MI52-M_u3 net84 S1 VDD VDD p w=0.685u l=0.18u
MI53-M_u3 PG1 S1 OUT VDD p w=0.685u l=0.18u
.ends
.subckt MUX3D1BWP7T I0 I1 I2 S0 S1 Z VDD VSS 
MI53-M_u2 PG1 net35 OUT VSS n w=0.5u l=0.18u
MI51-M_u2 Z OUT VSS VSS n w=1u l=0.18u
MI50-M_u2 net39 S0 VSS VSS n w=0.5u l=0.18u
MI52-M_u2 net35 S1 VSS VSS n w=0.5u l=0.18u
MI44 PG1 S0 net54 VSS n w=0.5u l=0.18u
MI45 net45 I2 VSS VSS n w=1u l=0.18u
MI46 OUT S1 net45 VSS n w=0.5u l=0.18u
MI43 PG1 net39 net50 VSS n w=0.665u l=0.18u
MI42 net54 I1 VSS VSS n w=1u l=0.18u
MI41 net50 I0 VSS VSS n w=0.665u l=0.18u
MI53-M_u3 PG1 S1 OUT VDD p w=0.685u l=0.18u
MI51-M_u3 Z OUT VDD VDD p w=1.37u l=0.18u
MI50-M_u3 net39 S0 VDD VDD p w=0.685u l=0.18u
MI52-M_u3 net35 S1 VDD VDD p w=0.685u l=0.18u
MI38 net70 I1 VDD VDD p w=1.37u l=0.18u
MI39 net62 I2 VDD VDD p w=1.37u l=0.18u
MI40 OUT net35 net62 VDD p w=0.685u l=0.18u
MI35 net74 I0 VDD VDD p w=1.27u l=0.18u
MI36 PG1 S0 net74 VDD p w=0.685u l=0.18u
MI37 PG1 net39 net70 VDD p w=0.685u l=0.18u
.ends
.subckt MUX3D2BWP7T I0 I1 I2 S0 S1 Z VDD VSS 
MI51_0-M_u2 Z OUT VSS VSS n w=1u l=0.18u
MI51_1-M_u2 Z OUT VSS VSS n w=1u l=0.18u
MI50-M_u2 net40 S0 VSS VSS n w=0.5u l=0.18u
MI52-M_u2 net38 S1 VSS VSS n w=0.5u l=0.18u
MI53-M_u2 PG1 net38 OUT VSS n w=0.57u l=0.18u
MI44 PG1 S0 net52 VSS n w=0.62u l=0.18u
MI45 net57 I2 VSS VSS n w=0.925u l=0.18u
MI46 OUT S1 net57 VSS n w=0.925u l=0.18u
MI43 PG1 net40 net54 VSS n w=1u l=0.18u
MI42 net52 I1 VSS VSS n w=1u l=0.18u
MI41 net54 I0 VSS VSS n w=1u l=0.18u
MI51_0-M_u3 Z OUT VDD VDD p w=1.37u l=0.18u
MI51_1-M_u3 Z OUT VDD VDD p w=1.37u l=0.18u
MI50-M_u3 net40 S0 VDD VDD p w=0.685u l=0.18u
MI52-M_u3 net38 S1 VDD VDD p w=0.685u l=0.18u
MI53-M_u3 PG1 S1 OUT VDD p w=1.05u l=0.18u
MI38 net81 I1 VDD VDD p w=1.37u l=0.18u
MI39 net78 I2 VDD VDD p w=1.37u l=0.18u
MI40 OUT net38 net78 VDD p w=1.37u l=0.18u
MI35 net71 I0 VDD VDD p w=1.37u l=0.18u
MI36 PG1 S0 net71 VDD p w=0.77u l=0.18u
MI37 PG1 net40 net81 VDD p w=1.37u l=0.18u
.ends
.subckt MUX3ND0BWP7T I0 I1 I2 S0 S1 ZN VDD VSS 
MI41 net40 I0 VSS VSS n w=0.665u l=0.18u
MI42 net37 I1 VSS VSS n w=0.5u l=0.18u
MI43 PG1 net69 net40 VSS n w=0.665u l=0.18u
MI44 PG1 S0 net37 VSS n w=0.5u l=0.18u
MI45 net35 I2 VSS VSS n w=0.5u l=0.18u
MI46 ZN S1 net35 VSS n w=0.5u l=0.18u
MI50-M_u2 net69 S0 VSS VSS n w=0.5u l=0.18u
MI52-M_u2 net67 S1 VSS VSS n w=0.5u l=0.18u
MI53-M_u2 PG1 net67 ZN VSS n w=0.5u l=0.18u
MI35 net64 I0 VDD VDD p w=0.685u l=0.18u
MI36 PG1 S0 net64 VDD p w=0.685u l=0.18u
MI37 PG1 net69 net55 VDD p w=0.685u l=0.18u
MI38 net55 I1 VDD VDD p w=0.685u l=0.18u
MI39 net51 I2 VDD VDD p w=0.685u l=0.18u
MI40 ZN net67 net51 VDD p w=0.685u l=0.18u
MI50-M_u3 net69 S0 VDD VDD p w=0.685u l=0.18u
MI52-M_u3 net67 S1 VDD VDD p w=0.685u l=0.18u
MI53-M_u3 PG1 S1 ZN VDD p w=0.685u l=0.18u
.ends
.subckt MUX3ND1BWP7T I0 I1 I2 S0 S1 ZN VDD VSS 
MI44 PG1 S0 net066 VSS n w=0.5u l=0.18u
MI45 net064 I2 VSS VSS n w=1u l=0.18u
MI46 net59 S1 net064 VSS n w=0.5u l=0.18u
MI43 PG1 net075 net052 VSS n w=0.665u l=0.18u
MI42 net066 I1 VSS VSS n w=1u l=0.18u
MI41 net052 I0 VSS VSS n w=0.665u l=0.18u
MI3-M_u2 net33 net59 VSS VSS n w=1u l=0.18u
MI50-M_u2 net075 S0 VSS VSS n w=0.5u l=0.18u
MI52-M_u2 net073 S1 VSS VSS n w=0.5u l=0.18u
MU18-M_u2 ZN net33 VSS VSS n w=1u l=0.18u
MI53-M_u2 PG1 net073 net59 VSS n w=0.5u l=0.18u
MI38 net048 I1 VDD VDD p w=1.37u l=0.18u
MI39 net044 I2 VDD VDD p w=1.37u l=0.18u
MI40 net59 net073 net044 VDD p w=0.685u l=0.18u
MI35 net038 I0 VDD VDD p w=1.27u l=0.18u
MI36 PG1 S0 net038 VDD p w=0.685u l=0.18u
MI37 PG1 net075 net048 VDD p w=0.685u l=0.18u
MI3-M_u3 net33 net59 VDD VDD p w=1.37u l=0.18u
MI50-M_u3 net075 S0 VDD VDD p w=0.685u l=0.18u
MI52-M_u3 net073 S1 VDD VDD p w=0.685u l=0.18u
MU18-M_u3 ZN net33 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 PG1 S1 net59 VDD p w=0.685u l=0.18u
.ends
.subckt MUX3ND2BWP7T I0 I1 I2 S0 S1 ZN VDD VSS 
MI52-M_u2 net044 S1 VSS VSS n w=0.5u l=0.18u
MI3-M_u2 net33 net079 VSS VSS n w=1u l=0.18u
MI50-M_u2 net046 S0 VSS VSS n w=0.5u l=0.18u
MU18_0-M_u2 ZN net33 VSS VSS n w=1u l=0.18u
MU18_1-M_u2 ZN net33 VSS VSS n w=1u l=0.18u
MI53-M_u2 PG1 net044 net079 VSS n w=0.655u l=0.18u
MI44 PG1 S0 net067 VSS n w=0.89u l=0.18u
MI45 net061 I2 VSS VSS n w=1u l=0.18u
MI46 net079 S1 net061 VSS n w=0.94u l=0.18u
MI43 PG1 net046 net053 VSS n w=0.665u l=0.18u
MI42 net067 I1 VSS VSS n w=1u l=0.18u
MI41 net053 I0 VSS VSS n w=0.665u l=0.18u
MI52-M_u3 net044 S1 VDD VDD p w=0.685u l=0.18u
MI3-M_u3 net33 net079 VDD VDD p w=1.37u l=0.18u
MI50-M_u3 net046 S0 VDD VDD p w=0.685u l=0.18u
MU18_0-M_u3 ZN net33 VDD VDD p w=1.37u l=0.18u
MU18_1-M_u3 ZN net33 VDD VDD p w=1.37u l=0.18u
MI53-M_u3 PG1 S1 net079 VDD p w=0.95u l=0.18u
MI38 net072 I1 VDD VDD p w=1.37u l=0.18u
MI39 net082 I2 VDD VDD p w=1.37u l=0.18u
MI40 net079 net044 net082 VDD p w=1.285u l=0.18u
MI35 net075 I0 VDD VDD p w=1.27u l=0.18u
MI36 PG1 S0 net075 VDD p w=0.84u l=0.18u
MI37 PG1 net046 net072 VDD p w=0.84u l=0.18u
.ends
.subckt MUX4D0BWP7T I0 I1 I2 I3 S0 S1 Z VDD VSS 
MI19 net91 I0 VSS VSS n w=0.5u l=0.18u
MI20 net88 I1 VSS VSS n w=0.5u l=0.18u
MI12 PG1 net97 net91 VSS n w=0.5u l=0.18u
MI21 PG1 S0 net88 VSS n w=0.5u l=0.18u
MI52 PG2 S0 net73 VSS n w=0.5u l=0.18u
MI53 PG2 net97 net75 VSS n w=0.5u l=0.18u
MI54 net73 I3 VSS VSS n w=0.5u l=0.18u
MI55 net75 I2 VSS VSS n w=0.5u l=0.18u
MI15-M_u2 net97 S0 VSS VSS n w=0.5u l=0.18u
MI59-M_u2 net95 S1 VSS VSS n w=0.5u l=0.18u
MI60-M_u2 Z net101 VSS VSS n w=0.5u l=0.18u
MI61-M_u2 PG2 S1 net101 VSS n w=0.5u l=0.18u
MI62-M_u2 PG1 net95 net101 VSS n w=0.5u l=0.18u
MI111 net65 I0 VDD VDD p w=0.685u l=0.18u
MI5 PG1 S0 net65 VDD p w=0.685u l=0.18u
MI25 PG1 net97 net62 VDD p w=0.685u l=0.18u
MI24 net62 I1 VDD VDD p w=0.685u l=0.18u
MI48 net53 I3 VDD VDD p w=0.685u l=0.18u
MI49 PG2 net97 net53 VDD p w=0.685u l=0.18u
MI50 PG2 S0 net45 VDD p w=0.685u l=0.18u
MI51 net45 I2 VDD VDD p w=0.685u l=0.18u
MI15-M_u3 net97 S0 VDD VDD p w=0.685u l=0.18u
MI59-M_u3 net95 S1 VDD VDD p w=0.685u l=0.18u
MI60-M_u3 Z net101 VDD VDD p w=0.685u l=0.18u
MI61-M_u3 PG2 net95 net101 VDD p w=0.685u l=0.18u
MI62-M_u3 PG1 S1 net101 VDD p w=0.685u l=0.18u
.ends
.subckt MUX4D1BWP7T I0 I1 I2 I3 S0 S1 Z VDD VSS 
MI64 net81 I1 VSS VSS n w=0.79u l=0.18u
MI65 PG1 S0 net81 VSS n w=0.5u l=0.18u
MI68 net73 I3 VSS VSS n w=1u l=0.18u
MI63 net84 I0 VSS VSS n w=0.5u l=0.18u
MI66 PG2 S0 net73 VSS n w=0.5u l=0.18u
MI12 PG1 net97 net84 VSS n w=0.5u l=0.18u
MI67 PG2 net97 net70 VSS n w=0.5u l=0.18u
MI69 net70 I2 VSS VSS n w=0.5u l=0.18u
MI73-M_u2 net97 S0 VSS VSS n w=0.5u l=0.18u
MI74-M_u2 net95 S1 VSS VSS n w=0.5u l=0.18u
MI75-M_u2 Z net105 VSS VSS n w=1u l=0.18u
MI76-M_u2 PG2 S1 net105 VSS n w=0.5u l=0.18u
MI77-M_u2 PG1 net95 net105 VSS n w=0.5u l=0.18u
MI5 PG1 S0 net65 VDD p w=0.685u l=0.18u
MI62 net45 I2 VDD VDD p w=0.685u l=0.18u
MI111 net65 I0 VDD VDD p w=0.7u l=0.18u
MI61 PG2 S0 net45 VDD p w=0.685u l=0.18u
MI60 PG2 net97 net53 VDD p w=0.685u l=0.18u
MI59 net53 I3 VDD VDD p w=1.13u l=0.18u
MI58 net62 I1 VDD VDD p w=1.13u l=0.18u
MI25 PG1 net97 net62 VDD p w=0.685u l=0.18u
MI73-M_u3 net97 S0 VDD VDD p w=0.635u l=0.18u
MI74-M_u3 net95 S1 VDD VDD p w=0.685u l=0.18u
MI75-M_u3 Z net105 VDD VDD p w=1.37u l=0.18u
MI76-M_u3 PG2 net95 net105 VDD p w=0.685u l=0.18u
MI77-M_u3 PG1 S1 net105 VDD p w=0.685u l=0.18u
.ends
.subckt MUX4D2BWP7T I0 I1 I2 I3 S0 S1 Z VDD VSS 
MI64 net63 I1 VSS VSS n w=2u l=0.18u
MI65 PG1 S0 net63 VSS n w=0.5u l=0.18u
MI68 net54 I3 VSS VSS n w=2u l=0.18u
MI63 net51 I0 VSS VSS n w=2u l=0.18u
MI66 PG2 S0 net54 VSS n w=0.5u l=0.18u
MI12 PG1 net97 net51 VSS n w=0.5u l=0.18u
MI67 PG2 net97 net48 VSS n w=0.5u l=0.18u
MI69 net48 I2 VSS VSS n w=2u l=0.18u
MI73-M_u2 net97 S0 VSS VSS n w=0.5u l=0.18u
MI74-M_u2 net95 S1 VSS VSS n w=0.5u l=0.18u
MI75_0-M_u2 Z net105 VSS VSS n w=1u l=0.18u
MI75_1-M_u2 Z net105 VSS VSS n w=1u l=0.18u
MI76-M_u2 PG2 S1 net105 VSS n w=0.5u l=0.18u
MI77-M_u2 PG1 net95 net105 VSS n w=0.5u l=0.18u
MI5 PG1 S0 net84 VDD p w=0.685u l=0.18u
MI62 net83 I2 VDD VDD p w=2.715u l=0.18u
MI111 net84 I0 VDD VDD p w=2.74u l=0.18u
MI61 PG2 S0 net83 VDD p w=0.685u l=0.18u
MI60 PG2 net97 net75 VDD p w=0.685u l=0.18u
MI59 net75 I3 VDD VDD p w=2.74u l=0.18u
MI58 net72 I1 VDD VDD p w=2.74u l=0.18u
MI25 PG1 net97 net72 VDD p w=0.685u l=0.18u
MI73-M_u3 net97 S0 VDD VDD p w=0.635u l=0.18u
MI74-M_u3 net95 S1 VDD VDD p w=0.685u l=0.18u
MI75_0-M_u3 Z net105 VDD VDD p w=1.37u l=0.18u
MI75_1-M_u3 Z net105 VDD VDD p w=1.37u l=0.18u
MI76-M_u3 PG2 net95 net105 VDD p w=0.685u l=0.18u
MI77-M_u3 PG1 S1 net105 VDD p w=0.685u l=0.18u
.ends
.subckt MUX4ND0BWP7T I0 I1 I2 I3 S0 S1 ZN VDD VSS 
MI64 net62 I1 VSS VSS n w=0.79u l=0.18u
MI65 PG1 S0 net62 VSS n w=0.5u l=0.18u
MI68 net53 I3 VSS VSS n w=0.705u l=0.18u
MI63 net57 I0 VSS VSS n w=0.5u l=0.18u
MI66 PG2 S0 net53 VSS n w=0.5u l=0.18u
MI12 PG1 net94 net57 VSS n w=0.5u l=0.18u
MI67 PG2 net94 net45 VSS n w=0.5u l=0.18u
MI69 net45 I2 VSS VSS n w=0.8u l=0.18u
MI73-M_u2 net94 S0 VSS VSS n w=0.5u l=0.18u
MI74-M_u2 net92 S1 VSS VSS n w=0.5u l=0.18u
MI76-M_u2 PG2 S1 ZN VSS n w=0.5u l=0.18u
MI77-M_u2 PG1 net92 ZN VSS n w=0.5u l=0.18u
MI5 PG1 S0 net83 VDD p w=0.685u l=0.18u
MI62 net82 I2 VDD VDD p w=0.685u l=0.18u
MI111 net83 I0 VDD VDD p w=0.685u l=0.18u
MI61 PG2 S0 net82 VDD p w=0.685u l=0.18u
MI60 PG2 net94 net74 VDD p w=0.685u l=0.18u
MI59 net74 I3 VDD VDD p w=1.13u l=0.18u
MI58 net70 I1 VDD VDD p w=0.685u l=0.18u
MI25 PG1 net94 net70 VDD p w=0.685u l=0.18u
MI73-M_u3 net94 S0 VDD VDD p w=0.685u l=0.18u
MI74-M_u3 net92 S1 VDD VDD p w=0.685u l=0.18u
MI76-M_u3 PG2 net92 ZN VDD p w=0.685u l=0.18u
MI77-M_u3 PG1 S1 ZN VDD p w=0.685u l=0.18u
.ends
.subckt MUX4ND1BWP7T I0 I1 I2 I3 S0 S1 ZN VDD VSS 
MI64 net060 I1 VSS VSS n w=0.79u l=0.18u
MI65 net063 S0 net060 VSS n w=0.5u l=0.18u
MI68 net071 I3 VSS VSS n w=1u l=0.18u
MI63 net074 I0 VSS VSS n w=0.5u l=0.18u
MI66 net0107 S0 net071 VSS n w=0.5u l=0.18u
MI12 net063 net0123 net074 VSS n w=0.5u l=0.18u
MI67 net0107 net0123 net081 VSS n w=0.5u l=0.18u
MI69 net081 I2 VSS VSS n w=0.5u l=0.18u
MI41 net085 net0107 VSS VSS n w=1u l=0.18u
MI44 net59 net0121 net089 VSS n w=0.5u l=0.18u
MI43 net089 net063 VSS VSS n w=1u l=0.18u
MI42 net59 S1 net085 VSS n w=0.5u l=0.18u
MI73-M_u2 net0123 S0 VSS VSS n w=0.5u l=0.18u
MI51-M_u2 net0121 S1 VSS VSS n w=0.5u l=0.18u
MI36-M_u2 ZN net59 VSS VSS n w=1u l=0.18u
MI46 net089 net063 VDD VDD p w=1.22u l=0.18u
MI5 net063 S0 net0101 VDD p w=0.685u l=0.18u
MI62 net0106 I2 VDD VDD p w=0.685u l=0.18u
MI111 net0101 I0 VDD VDD p w=0.685u l=0.18u
MI61 net0107 S0 net0106 VDD p w=0.685u l=0.18u
MI60 net0107 net0123 net0110 VDD p w=0.685u l=0.18u
MI59 net0110 I3 VDD VDD p w=1.13u l=0.18u
MI58 net0118 I1 VDD VDD p w=1.13u l=0.18u
MI25 net063 net0123 net0118 VDD p w=0.685u l=0.18u
MI47 net085 net0107 VDD VDD p w=1.22u l=0.18u
MI48 net59 net0121 net085 VDD p w=0.685u l=0.18u
MI45 net59 S1 net089 VDD p w=0.685u l=0.18u
MI73-M_u3 net0123 S0 VDD VDD p w=0.635u l=0.18u
MI51-M_u3 net0121 S1 VDD VDD p w=0.685u l=0.18u
MI36-M_u3 ZN net59 VDD VDD p w=1.37u l=0.18u
.ends
.subckt MUX4ND2BWP7T I0 I1 I2 I3 S0 S1 ZN VDD VSS 
MI41 net052 net0105 VSS VSS n w=1u l=0.18u
MI44 net77 net0121 net087 VSS n w=0.5u l=0.18u
MI43 net087 net056 VSS VSS n w=1u l=0.18u
MI68 net0111 I3 VSS VSS n w=1u l=0.18u
MI63 net0108 I0 VSS VSS n w=0.5u l=0.18u
MI66 net0105 S0 net0111 VSS n w=0.5u l=0.18u
MI12 net056 net0123 net0108 VSS n w=0.5u l=0.18u
MI42 net77 S1 net052 VSS n w=0.5u l=0.18u
MI64 net0113 I1 VSS VSS n w=0.79u l=0.18u
MI65 net056 S0 net0113 VSS n w=0.5u l=0.18u
MI67 net0105 net0123 net098 VSS n w=0.5u l=0.18u
MI69 net098 I2 VSS VSS n w=0.5u l=0.18u
MI73-M_u2 net0123 S0 VSS VSS n w=0.5u l=0.18u
MI51-M_u2 net0121 S1 VSS VSS n w=0.5u l=0.18u
MU18_0-M_u2 ZN net77 VSS VSS n w=1u l=0.18u
MU18_1-M_u2 ZN net77 VSS VSS n w=1u l=0.18u
MI58 net058 I1 VDD VDD p w=1.13u l=0.18u
MI47 net052 net0105 VDD VDD p w=1.235u l=0.18u
MI45 net77 S1 net087 VDD p w=0.685u l=0.18u
MI46 net087 net056 VDD VDD p w=1.235u l=0.18u
MI62 net074 I2 VDD VDD p w=0.685u l=0.18u
MI61 net0105 S0 net074 VDD p w=0.685u l=0.18u
MI59 net062 I3 VDD VDD p w=1.13u l=0.18u
MI48 net77 net0121 net052 VDD p w=0.685u l=0.18u
MI25 net056 net0123 net058 VDD p w=0.685u l=0.18u
MI5 net056 S0 net079 VDD p w=0.685u l=0.18u
MI111 net079 I0 VDD VDD p w=0.685u l=0.18u
MI60 net0105 net0123 net062 VDD p w=0.685u l=0.18u
MI73-M_u3 net0123 S0 VDD VDD p w=0.635u l=0.18u
MI51-M_u3 net0121 S1 VDD VDD p w=0.635u l=0.18u
MU18_0-M_u3 ZN net77 VDD VDD p w=1.37u l=0.18u
MU18_1-M_u3 ZN net77 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND2D0BWP7T A1 A2 ZN VDD VSS 
MI0-M_u4 XI0-net6 A2 VSS VSS n w=0.5u l=0.18u
MI0-M_u3 ZN A1 XI0-net6 VSS n w=0.5u l=0.18u
MI0-M_u2 ZN A2 VDD VDD p w=0.685u l=0.18u
MI0-M_u1 ZN A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt ND2D1BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 XI1-net6 A2 VSS VSS n w=1u l=0.18u
MI1-M_u3 ZN A1 XI1-net6 VSS n w=1u l=0.18u
MI1-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
MI1-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND2D1P5BWP7T A1 A2 ZN VDD VSS 
MI8 ZN A1 net018 VSS n w=0.75u l=0.18u
MI7 net018 A2 VSS VSS n w=0.75u l=0.18u
MI6 net8 A2 VSS VSS n w=0.75u l=0.18u
MI5 ZN A1 net8 VSS n w=0.75u l=0.18u
MI3 ZN A1 VDD VDD p w=2.055u l=0.18u
MU19 ZN A2 VDD VDD p w=2.055u l=0.18u
.ends
.subckt ND2D2BWP7T A1 A2 ZN VDD VSS 
MU3_0-M_u4 XU3_0-net6 A2 VSS VSS n w=1u l=0.18u
MU3_0-M_u3 ZN A1 XU3_0-net6 VSS n w=1u l=0.18u
MU3_1-M_u4 XU3_1-net6 A2 VSS VSS n w=1u l=0.18u
MU3_1-M_u3 ZN A1 XU3_1-net6 VSS n w=1u l=0.18u
MU3_0-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
MU3_0-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
MU3_1-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
MU3_1-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND2D2P5BWP7T A1 A2 ZN VDD VSS 
MI8 net26 A2 VSS VSS n w=0.835u l=0.18u
MI7 ZN A1 net26 VSS n w=0.835u l=0.18u
MU14 net41 A2 VSS VSS n w=0.835u l=0.18u
MI6 net38 A2 VSS VSS n w=0.835u l=0.18u
MI5 ZN A1 net38 VSS n w=0.835u l=0.18u
MI4 ZN A1 net41 VSS n w=0.835u l=0.18u
MI11 ZN A1 VDD VDD p w=3.425u l=0.18u
MI9 ZN A2 VDD VDD p w=3.425u l=0.18u
.ends
.subckt ND2D3BWP7T A1 A2 ZN VDD VSS 
MI2_0 net19 A2 VSS VSS n w=1u l=0.18u
MI2_1 net19 A2 VSS VSS n w=1u l=0.18u
MI2_2 net19 A2 VSS VSS n w=1u l=0.18u
MI3_0 ZN A1 net19 VSS n w=1u l=0.18u
MI3_1 ZN A1 net19 VSS n w=1u l=0.18u
MI3_2 ZN A1 net19 VSS n w=1u l=0.18u
MI4_0 ZN A2 VDD VDD p w=1.37u l=0.18u
MI4_1 ZN A2 VDD VDD p w=1.37u l=0.18u
MI4_2 ZN A2 VDD VDD p w=1.37u l=0.18u
MI5_0 ZN A1 VDD VDD p w=1.37u l=0.18u
MI5_1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI5_2 ZN A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND2D4BWP7T A1 A2 ZN VDD VSS 
MI2_0 net19 A2 VSS VSS n w=1u l=0.18u
MI2_1 net19 A2 VSS VSS n w=1u l=0.18u
MI2_2 net19 A2 VSS VSS n w=1u l=0.18u
MI2_3 net19 A2 VSS VSS n w=1u l=0.18u
MI3_0 ZN A1 net19 VSS n w=1u l=0.18u
MI3_1 ZN A1 net19 VSS n w=1u l=0.18u
MI3_2 ZN A1 net19 VSS n w=1u l=0.18u
MI3_3 ZN A1 net19 VSS n w=1u l=0.18u
MI4_0 ZN A2 VDD VDD p w=1.37u l=0.18u
MI4_1 ZN A2 VDD VDD p w=1.37u l=0.18u
MI4_2 ZN A2 VDD VDD p w=1.37u l=0.18u
MI4_3 ZN A2 VDD VDD p w=1.37u l=0.18u
MI5_0 ZN A1 VDD VDD p w=1.37u l=0.18u
MI5_1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI5_2 ZN A1 VDD VDD p w=1.37u l=0.18u
MI5_3 ZN A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND2D5BWP7T A1 A2 ZN VDD VSS 
MI5 ZN A1 net11 VSS n w=5u l=0.18u
MI6 net11 A2 VSS VSS n w=5u l=0.18u
MU19 ZN A2 VDD VDD p w=6.85u l=0.18u
MI11 ZN A1 VDD VDD p w=6.85u l=0.18u
.ends
.subckt ND2D6BWP7T A1 A2 ZN VDD VSS 
MI2 ZN A1 net20 VSS n w=6u l=0.18u
MI3 net20 A2 VSS VSS n w=6u l=0.18u
MI11 ZN A1 VDD VDD p w=8.22u l=0.18u
MU19 ZN A2 VDD VDD p w=8.22u l=0.18u
.ends
.subckt ND2D8BWP7T A1 A2 ZN VDD VSS 
MI13_0 ZN A1 net66 VSS n w=1u l=0.18u
MI13_1 ZN A1 net66 VSS n w=1u l=0.18u
MI13_2 ZN A1 net66 VSS n w=1u l=0.18u
MI13_3 ZN A1 net66 VSS n w=1u l=0.18u
MI13_4 ZN A1 net66 VSS n w=1u l=0.18u
MI13_5 ZN A1 net66 VSS n w=1u l=0.18u
MI13_6 ZN A1 net66 VSS n w=1u l=0.18u
MI13_7 ZN A1 net66 VSS n w=1u l=0.18u
MI14_0 net66 A2 VSS VSS n w=1u l=0.18u
MI14_1 net66 A2 VSS VSS n w=1u l=0.18u
MI14_2 net66 A2 VSS VSS n w=1u l=0.18u
MI14_3 net66 A2 VSS VSS n w=1u l=0.18u
MI14_4 net66 A2 VSS VSS n w=1u l=0.18u
MI14_5 net66 A2 VSS VSS n w=1u l=0.18u
MI14_6 net66 A2 VSS VSS n w=1u l=0.18u
MI14_7 net66 A2 VSS VSS n w=1u l=0.18u
M_u2_0 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_1 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_2 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_3 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_4 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_5 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_6 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_7 ZN A2 VDD VDD p w=1.37u l=0.18u
MI6_0 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_2 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_3 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_4 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_5 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_6 ZN A1 VDD VDD p w=1.37u l=0.18u
MI6_7 ZN A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND3D0BWP7T A1 A2 A3 ZN VDD VSS 
MI0-M_u4 ZN A1 XI0-net10 VSS n w=0.5u l=0.18u
MI0-M_u5 XI0-net10 A2 XI0-net13 VSS n w=0.5u l=0.18u
MI0-M_u6 XI0-net13 A3 VSS VSS n w=0.5u l=0.18u
MI0-M_u3 ZN A3 VDD VDD p w=0.685u l=0.18u
MI0-M_u1 ZN A1 VDD VDD p w=0.685u l=0.18u
MI0-M_u2 ZN A2 VDD VDD p w=0.685u l=0.18u
.ends
.subckt ND3D1BWP7T A1 A2 A3 ZN VDD VSS 
MI1-M_u4 ZN A1 XI1-net10 VSS n w=1u l=0.18u
MI1-M_u5 XI1-net10 A2 XI1-net13 VSS n w=1u l=0.18u
MI1-M_u6 XI1-net13 A3 VSS VSS n w=1u l=0.18u
MI1-M_u3 ZN A3 VDD VDD p w=1.37u l=0.18u
MI1-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND3D2BWP7T A1 A2 A3 ZN VDD VSS 
MI0_0-M_u4 ZN A1 XI0_0-net10 VSS n w=1u l=0.18u
MI0_0-M_u5 XI0_0-net10 A2 XI0_0-net13 VSS n w=1u l=0.18u
MI0_0-M_u6 XI0_0-net13 A3 VSS VSS n w=1u l=0.18u
MI0_1-M_u4 ZN A1 XI0_1-net10 VSS n w=1u l=0.18u
MI0_1-M_u5 XI0_1-net10 A2 XI0_1-net13 VSS n w=1u l=0.18u
MI0_1-M_u6 XI0_1-net13 A3 VSS VSS n w=1u l=0.18u
MI0_0-M_u3 ZN A3 VDD VDD p w=1.37u l=0.18u
MI0_0-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI0_0-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
MI0_1-M_u3 ZN A3 VDD VDD p w=1.37u l=0.18u
MI0_1-M_u1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI0_1-M_u2 ZN A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND3D3BWP7T A1 A2 A3 ZN VDD VSS 
M_u6_0 net051 A3 VSS VSS n w=1u l=0.18u
M_u6_1 net051 A3 VSS VSS n w=1u l=0.18u
M_u6_2 net051 A3 VSS VSS n w=1u l=0.18u
M_u4_0 ZN A1 net054 VSS n w=1u l=0.18u
M_u4_1 ZN A1 net054 VSS n w=1u l=0.18u
M_u4_2 ZN A1 net054 VSS n w=1u l=0.18u
M_u5_0 net054 A2 net051 VSS n w=1u l=0.18u
M_u5_1 net054 A2 net051 VSS n w=1u l=0.18u
M_u5_2 net054 A2 net051 VSS n w=1u l=0.18u
M_u1_0 ZN A1 VDD VDD p w=1.37u l=0.18u
M_u1_1 ZN A1 VDD VDD p w=1.37u l=0.18u
M_u1_2 ZN A1 VDD VDD p w=1.37u l=0.18u
M_u2_0 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_1 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_2 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u3_0 ZN A3 VDD VDD p w=1.37u l=0.18u
M_u3_1 ZN A3 VDD VDD p w=1.37u l=0.18u
M_u3_2 ZN A3 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND3D4BWP7T A1 A2 A3 ZN VDD VSS 
M_u6_0 net051 A3 VSS VSS n w=1u l=0.18u
M_u6_1 net051 A3 VSS VSS n w=1u l=0.18u
M_u6_2 net051 A3 VSS VSS n w=1u l=0.18u
M_u6_3 net051 A3 VSS VSS n w=1u l=0.18u
M_u4_0 ZN A1 net054 VSS n w=1u l=0.18u
M_u4_1 ZN A1 net054 VSS n w=1u l=0.18u
M_u4_2 ZN A1 net054 VSS n w=1u l=0.18u
M_u4_3 ZN A1 net054 VSS n w=1u l=0.18u
M_u5_0 net054 A2 net051 VSS n w=1u l=0.18u
M_u5_1 net054 A2 net051 VSS n w=1u l=0.18u
M_u5_2 net054 A2 net051 VSS n w=1u l=0.18u
M_u5_3 net054 A2 net051 VSS n w=1u l=0.18u
M_u1_0 ZN A1 VDD VDD p w=1.37u l=0.18u
M_u1_1 ZN A1 VDD VDD p w=1.37u l=0.18u
M_u1_2 ZN A1 VDD VDD p w=1.37u l=0.18u
M_u1_3 ZN A1 VDD VDD p w=1.37u l=0.18u
M_u2_0 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_1 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_2 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u2_3 ZN A2 VDD VDD p w=1.37u l=0.18u
M_u3_0 ZN A3 VDD VDD p w=1.37u l=0.18u
M_u3_1 ZN A3 VDD VDD p w=1.37u l=0.18u
M_u3_2 ZN A3 VDD VDD p w=1.37u l=0.18u
M_u3_3 ZN A3 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND4D0BWP7T A1 A2 A3 A4 ZN VDD VSS 
MI13 p2 A4 VSS VSS n w=0.5u l=0.18u
MI11 p0 A2 p1 VSS n w=0.5u l=0.18u
MI12 p1 A3 p2 VSS n w=0.5u l=0.18u
MU53 ZN A1 p0 VSS n w=0.5u l=0.18u
MI7 ZN A1 VDD VDD p w=0.685u l=0.18u
MI6 ZN A2 VDD VDD p w=0.685u l=0.18u
MI8 ZN A3 VDD VDD p w=0.685u l=0.18u
MI9 ZN A4 VDD VDD p w=0.685u l=0.18u
.ends
.subckt ND4D1BWP7T A1 A2 A3 A4 ZN VDD VSS 
MI5 p2 A4 VSS VSS n w=1u l=0.18u
MI3 p0 A2 p1 VSS n w=1u l=0.18u
MI4 p1 A3 p2 VSS n w=1u l=0.18u
MU53 ZN A1 p0 VSS n w=1u l=0.18u
MI7 ZN A1 VDD VDD p w=1.37u l=0.18u
MI2 ZN A4 VDD VDD p w=1.37u l=0.18u
MI1 ZN A3 VDD VDD p w=1.37u l=0.18u
MI0 ZN A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND4D2BWP7T A1 A2 A3 A4 ZN VDD VSS 
MI5 p2 A4 VSS VSS n w=2u l=0.18u
MI3 p0 A2 p1 VSS n w=2u l=0.18u
MI4 p1 A3 p2 VSS n w=2u l=0.18u
MU53 ZN A1 p0 VSS n w=2u l=0.18u
MI7 ZN A1 VDD VDD p w=2.74u l=0.18u
MI2 ZN A4 VDD VDD p w=2.74u l=0.18u
MI1 ZN A3 VDD VDD p w=2.74u l=0.18u
MI0 ZN A2 VDD VDD p w=2.74u l=0.18u
.ends
.subckt ND4D3BWP7T A1 A2 A3 A4 ZN VDD VSS 
MI16 net032 A4 VSS VSS n w=3u l=0.18u
MI17 net037 A3 net032 VSS n w=3u l=0.18u
MI18 net67 A2 net037 VSS n w=3u l=0.18u
MI19 ZN A1 net67 VSS n w=3u l=0.18u
MI8_0 ZN A1 VDD VDD p w=1.37u l=0.18u
MI8_1 ZN A1 VDD VDD p w=1.37u l=0.18u
MI8_2 ZN A1 VDD VDD p w=1.37u l=0.18u
MI2_0 ZN A4 VDD VDD p w=1.37u l=0.18u
MI2_1 ZN A4 VDD VDD p w=1.37u l=0.18u
MI2_2 ZN A4 VDD VDD p w=1.37u l=0.18u
MI6_0 ZN A3 VDD VDD p w=1.37u l=0.18u
MI6_1 ZN A3 VDD VDD p w=1.37u l=0.18u
MI6_2 ZN A3 VDD VDD p w=1.37u l=0.18u
MI7_0 ZN A2 VDD VDD p w=1.37u l=0.18u
MI7_1 ZN A2 VDD VDD p w=1.37u l=0.18u
MI7_2 ZN A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt ND4D4BWP7T A1 A2 A3 A4 ZN VDD VSS 
MU3-M_u5 ZN A1 XU3-net23 VSS n w=4u l=0.18u
MU3-M_u6 XU3-net23 A2 XU3-net26 VSS n w=4u l=0.18u
MU3-M_u7 XU3-net26 A3 XU3-net29 VSS n w=4u l=0.18u
MU3-M_u8 XU3-net29 A4 VSS VSS n w=4u l=0.18u
MU3-M_u4 ZN A4 VDD VDD p w=5.48u l=0.18u
MU3-M_u3 ZN A3 VDD VDD p w=5.48u l=0.18u
MU3-M_u2 ZN A2 VDD VDD p w=5.47u l=0.18u
MU3-M_u1 ZN A1 VDD VDD p w=5.48u l=0.18u
.ends
.subckt NR2D0BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=0.5u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=0.5u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=0.685u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=0.685u l=0.18u
.ends
.subckt NR2D1BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=1u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=1u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=1.37u l=0.18u
.ends
.subckt NR2D1P5BWP7T A1 A2 ZN VDD VSS 
MI5 ZN A2 VSS VSS n w=1.5u l=0.18u
MU14 ZN A1 VSS VSS n w=1.5u l=0.18u
MI6 net023 A2 VDD VDD p w=1.03u l=0.18u
MI7 ZN A1 net023 VDD p w=1.03u l=0.18u
MI3 net15 A2 VDD VDD p w=1.03u l=0.18u
MU19 ZN A1 net15 VDD p w=1.03u l=0.18u
.ends
.subckt NR2D2BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=2u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=2u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=2.74u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=2.74u l=0.18u
.ends
.subckt NR2D2P5BWP7T A1 A2 ZN VDD VSS 
MI8 ZN A2 VSS VSS n w=2.5u l=0.18u
MI7 ZN A1 VSS VSS n w=2.5u l=0.18u
MI9 ZN A1 net072 VDD p w=1.14u l=0.18u
MI3 net32 A2 VDD VDD p w=1.14u l=0.18u
MI2 net29 A2 VDD VDD p w=1.14u l=0.18u
MU19 ZN A1 net32 VDD p w=1.14u l=0.18u
MU20 ZN A1 net29 VDD p w=1.14u l=0.18u
MI11 net072 A2 VDD VDD p w=1.14u l=0.18u
.ends
.subckt NR2D3BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=3u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=3u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=4.11u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=4.11u l=0.18u
.ends
.subckt NR2D4BWP7T A1 A2 ZN VDD VSS 
MI13 ZN A1 VSS VSS n w=4u l=0.18u
MI6 ZN A2 VSS VSS n w=4u l=0.18u
MI27 net20 A2 VDD VDD p w=5.48u l=0.18u
MI28 ZN A1 net20 VDD p w=5.48u l=0.18u
.ends
.subckt NR2D5BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=5u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=5u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=6.85u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=6.85u l=0.18u
.ends
.subckt NR2D6BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=6u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=6u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=8.22u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=8.22u l=0.18u
.ends
.subckt NR2D8BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=8u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=8u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=10.96u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=10.96u l=0.18u
.ends
.subckt NR2XD0BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=0.5u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=0.5u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=1.37u l=0.18u
.ends
.subckt NR2XD1BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=1u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=1u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=2.74u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=2.74u l=0.18u
.ends
.subckt NR2XD2BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=2u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=2u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=5.48u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=5.48u l=0.18u
.ends
.subckt NR2XD3BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=3u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=3u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=8.22u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=8.22u l=0.18u
.ends
.subckt NR2XD4BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=3.99u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=3.99u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=10.96u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=10.96u l=0.18u
.ends
.subckt NR2XD8BWP7T A1 A2 ZN VDD VSS 
MI1-M_u4 ZN A1 VSS VSS n w=8u l=0.18u
MI1-M_u3 ZN A2 VSS VSS n w=8u l=0.18u
MI1-M_u1 XI1-net8 A2 VDD VDD p w=21.92u l=0.18u
MI1-M_u2 ZN A1 XI1-net8 VDD p w=21.92u l=0.18u
.ends
.subckt NR3D0BWP7T A1 A2 A3 ZN VDD VSS 
M_u4 ZN A3 VSS VSS n w=0.5u l=0.18u
MI2 ZN A2 VSS VSS n w=0.5u l=0.18u
MI3 ZN A1 VSS VSS n w=0.5u l=0.18u
M_u1 net25 A3 VDD VDD p w=1.37u l=0.18u
MI0 net28 A2 net25 VDD p w=1.37u l=0.18u
MI1 ZN A1 net28 VDD p w=1.37u l=0.18u
.ends
.subckt NR3D1BWP7T A1 A2 A3 ZN VDD VSS 
M_u4 ZN A3 VSS VSS n w=1u l=0.18u
MI2 ZN A2 VSS VSS n w=1u l=0.18u
MI3 ZN A1 VSS VSS n w=1u l=0.18u
M_u1_0 net023[0] A3 VDD VDD p w=1.37u l=0.18u
M_u1_1 net023[1] A3 VDD VDD p w=1.37u l=0.18u
MI0_0 net026[0] A2 net023[0] VDD p w=1.37u l=0.18u
MI0_1 net026[1] A2 net023[1] VDD p w=1.37u l=0.18u
MI1_0 ZN A1 net026[0] VDD p w=1.37u l=0.18u
MI1_1 ZN A1 net026[1] VDD p w=1.37u l=0.18u
.ends
.subckt NR3D2BWP7T A1 A2 A3 ZN VDD VSS 
M_u4_0 ZN A3 VSS VSS n w=1u l=0.18u
M_u4_1 ZN A3 VSS VSS n w=1u l=0.18u
MI7_0 ZN A1 VSS VSS n w=1u l=0.18u
MI7_1 ZN A1 VSS VSS n w=1u l=0.18u
MI6_0 ZN A2 VSS VSS n w=1u l=0.18u
MI6_1 ZN A2 VSS VSS n w=1u l=0.18u
M_u1 net70 A3 VDD VDD p w=5.48u l=0.18u
MI20 net67 A2 net70 VDD p w=5.48u l=0.18u
MI21 ZN A1 net67 VDD p w=5.48u l=0.18u
.ends
.subckt NR3D3BWP7T A1 A2 A3 ZN VDD VSS 
MI0-M_u6 ZN A1 VSS VSS n w=3u l=0.18u
MI0-M_u5 ZN A2 VSS VSS n w=3u l=0.18u
MI0-M_u4 ZN A3 VSS VSS n w=3u l=0.18u
MI0-M_u1 XI0-net9 A3 VDD VDD p w=8.22u l=0.18u
MI0-M_u2 XI0-net12 A2 XI0-net9 VDD p w=8.225u l=0.18u
MI0-M_u3 ZN A1 XI0-net12 VDD p w=8.22u l=0.18u
.ends
.subckt NR3D4BWP7T A1 A2 A3 ZN VDD VSS 
MI0-M_u6 ZN A1 VSS VSS n w=3.99u l=0.18u
MI0-M_u5 ZN A2 VSS VSS n w=3.99u l=0.18u
MI0-M_u4 ZN A3 VSS VSS n w=3.99u l=0.18u
MI0-M_u1 XI0-net9 A3 VDD VDD p w=10.96u l=0.18u
MI0-M_u2 XI0-net12 A2 XI0-net9 VDD p w=11.2u l=0.18u
MI0-M_u3 ZN A1 XI0-net12 VDD p w=10.96u l=0.18u
.ends
.subckt NR4D0BWP7T A1 A2 A3 A4 ZN VDD VSS 
MI36 ZN A4 VSS VSS n w=0.5u l=0.18u
MI35 ZN A3 VSS VSS n w=0.5u l=0.18u
MI34 ZN A2 VSS VSS n w=0.5u l=0.18u
MI5 ZN A1 VSS VSS n w=0.5u l=0.18u
MI26 net49 A3 net52 VDD p w=1.37u l=0.18u
MI7 net52 A4 VDD VDD p w=1.37u l=0.18u
MI27 net46 A2 net49 VDD p w=1.37u l=0.18u
MI28 ZN A1 net46 VDD p w=1.37u l=0.18u
.ends
.subckt NR4D1BWP7T A1 A2 A3 A4 ZN VDD VSS 
MI36 ZN A4 VSS VSS n w=1u l=0.18u
MI35 ZN A3 VSS VSS n w=1u l=0.18u
MI34 ZN A2 VSS VSS n w=1u l=0.18u
MI5 ZN A1 VSS VSS n w=1u l=0.18u
MI26 net49 A3 net52 VDD p w=1.37u l=0.18u
MI30 net43 A2 net40 VDD p w=1.37u l=0.18u
MI31 net40 A3 net37 VDD p w=1.37u l=0.18u
MI32 net37 A4 VDD VDD p w=1.37u l=0.18u
MI29 ZN A1 net43 VDD p w=1.37u l=0.18u
MI7 net52 A4 VDD VDD p w=1.37u l=0.18u
MI27 net46 A2 net49 VDD p w=1.37u l=0.18u
MI28 ZN A1 net46 VDD p w=1.37u l=0.18u
.ends
.subckt NR4D2BWP7T A1 A2 A3 A4 ZN VDD VSS 
MI45_0 ZN A4 VSS VSS n w=1u l=0.18u
MI45_1 ZN A4 VSS VSS n w=1u l=0.18u
MI44_0 ZN A3 VSS VSS n w=1u l=0.18u
MI44_1 ZN A3 VSS VSS n w=1u l=0.18u
MI43_0 ZN A2 VSS VSS n w=1u l=0.18u
MI43_1 ZN A2 VSS VSS n w=1u l=0.18u
MI5_0 ZN A1 VSS VSS n w=1u l=0.18u
MI5_1 ZN A1 VSS VSS n w=1u l=0.18u
MI46_0 p1 A3 p0 VDD p w=1.37u l=0.18u
MI46_1 p1 A3 p0 VDD p w=1.37u l=0.18u
MI46_2 p1 A3 p0 VDD p w=1.37u l=0.18u
MI46_3 p1 A3 p0 VDD p w=1.37u l=0.18u
MI7_0 p0 A4 VDD VDD p w=1.37u l=0.18u
MI7_1 p0 A4 VDD VDD p w=1.37u l=0.18u
MI7_2 p0 A4 VDD VDD p w=1.37u l=0.18u
MI7_3 p0 A4 VDD VDD p w=1.37u l=0.18u
MI47_0 p2 A2 p1 VDD p w=1.37u l=0.18u
MI47_1 p2 A2 p1 VDD p w=1.37u l=0.18u
MI47_2 p2 A2 p1 VDD p w=1.37u l=0.18u
MI47_3 p2 A2 p1 VDD p w=1.37u l=0.18u
MI48_0 ZN A1 p2 VDD p w=1.37u l=0.18u
MI48_1 ZN A1 p2 VDD p w=1.37u l=0.18u
MI48_2 ZN A1 p2 VDD p w=1.37u l=0.18u
MI48_3 ZN A1 p2 VDD p w=1.37u l=0.18u
.ends
.subckt NR4D3BWP7T A1 A2 A3 A4 ZN VDD VSS 
MI48_0 ZN A4 VSS VSS n w=1u l=0.18u
MI48_1 ZN A4 VSS VSS n w=1u l=0.18u
MI48_2 ZN A4 VSS VSS n w=1u l=0.18u
MI47_0 ZN A3 VSS VSS n w=1u l=0.18u
MI47_1 ZN A3 VSS VSS n w=1u l=0.18u
MI47_2 ZN A3 VSS VSS n w=1u l=0.18u
MI46_0 ZN A2 VSS VSS n w=1u l=0.18u
MI46_1 ZN A2 VSS VSS n w=1u l=0.18u
MI46_2 ZN A2 VSS VSS n w=1u l=0.18u
MI42_0 ZN A1 VSS VSS n w=1u l=0.18u
MI42_1 ZN A1 VSS VSS n w=1u l=0.18u
MI42_2 ZN A1 VSS VSS n w=1u l=0.18u
MI43 net39 A3 net42 VDD p w=8.225u l=0.18u
MI7 net42 A4 VDD VDD p w=8.22u l=0.18u
MI44 net36 A2 net39 VDD p w=8.225u l=0.18u
MI45 ZN A1 net36 VDD p w=8.22u l=0.18u
.ends
.subckt NR4D4BWP7T A1 A2 A3 A4 ZN VDD VSS 
MI46-M_u4 ZN A4 VSS VSS n w=3.99u l=0.18u
MI46-M_u3 ZN A3 VSS VSS n w=3.99u l=0.18u
MI46-M_u5 ZN A2 VSS VSS n w=3.99u l=0.18u
MI46-M_u8 ZN A1 VSS VSS n w=3.99u l=0.18u
MI46-M_u7 ZN A1 XI46-net7 VDD p w=10.96u l=0.18u
MI46-M_u6 XI46-net7 A2 XI46-net10 VDD p w=11.2u l=0.18u
MI46-M_u2 XI46-net10 A3 XI46-net13 VDD p w=11.2u l=0.18u
MI46-M_u1 XI46-net13 A4 VDD VDD p w=10.96u l=0.18u
.ends
.subckt OA211D0BWP7T A1 A2 B C Z VDD VSS 
MI8 net36 B net24 VSS n w=0.5u l=0.18u
MI9 net24 C VSS VSS n w=0.5u l=0.18u
M_u2 net33 A1 net36 VSS n w=0.5u l=0.18u
MI7 net33 A2 net36 VSS n w=0.5u l=0.18u
MI11-M_u2 Z net33 VSS VSS n w=0.5u l=0.18u
MI11-M_u3 Z net33 VDD VDD p w=0.685u l=0.18u
MI6 net33 A2 net35 VDD p w=0.685u l=0.18u
MI5 net35 A1 VDD VDD p w=0.685u l=0.18u
MI4 net33 C VDD VDD p w=0.685u l=0.18u
M_u12 net33 B VDD VDD p w=0.685u l=0.18u
.ends
.subckt OA211D1BWP7T A1 A2 B C Z VDD VSS 
MI16 net36 B net24 VSS n w=1u l=0.18u
MI17 net24 C VSS VSS n w=1u l=0.18u
MI15 net33 A1 net36 VSS n w=1u l=0.18u
MI7 net33 A2 net36 VSS n w=1u l=0.18u
MI11-M_u2 Z net33 VSS VSS n w=1u l=0.18u
MI11-M_u3 Z net33 VDD VDD p w=1.37u l=0.18u
MI14 net33 A2 net35 VDD p w=1.37u l=0.18u
MI13 net35 A1 VDD VDD p w=1.37u l=0.18u
MI12 net33 C VDD VDD p w=1.37u l=0.18u
M_u12 net33 B VDD VDD p w=1.37u l=0.18u
.ends
.subckt OA211D2BWP7T A1 A2 B C Z VDD VSS 
MI16 net36 B net24 VSS n w=1u l=0.18u
MI17 net24 C VSS VSS n w=1u l=0.18u
MI15 net33 A1 net36 VSS n w=1u l=0.18u
MI7 net33 A2 net36 VSS n w=1u l=0.18u
MI11_0-M_u2 Z net33 VSS VSS n w=1u l=0.18u
MI11_1-M_u2 Z net33 VSS VSS n w=1u l=0.18u
MI11_0-M_u3 Z net33 VDD VDD p w=1.37u l=0.18u
MI11_1-M_u3 Z net33 VDD VDD p w=1.37u l=0.18u
MI14 net33 A2 net35 VDD p w=1.37u l=0.18u
MI13 net35 A1 VDD VDD p w=1.37u l=0.18u
MI12 net33 C VDD VDD p w=1.37u l=0.18u
M_u12 net33 B VDD VDD p w=1.37u l=0.18u
.ends
.subckt OA21D0BWP7T A1 A2 B Z VDD VSS 
MI15 net14 A2 net20 VSS n w=0.5u l=0.18u
MI11 net14 A1 net20 VSS n w=0.5u l=0.18u
MI16 net20 B VSS VSS n w=0.5u l=0.18u
MI8-M_u2 Z net14 VSS VSS n w=0.5u l=0.18u
MI8-M_u3 Z net14 VDD VDD p w=0.685u l=0.18u
M_u2 net14 B VDD VDD p w=0.685u l=0.18u
MI13 net24 A2 VDD VDD p w=0.685u l=0.18u
MI14 net14 A1 net24 VDD p w=0.685u l=0.18u
.ends
.subckt OA21D1BWP7T A1 A2 B Z VDD VSS 
MI12 net14 A2 net20 VSS n w=1u l=0.18u
MI11 net14 A1 net20 VSS n w=1u l=0.18u
MI6 net20 B VSS VSS n w=1u l=0.18u
MI8-M_u2 Z net14 VSS VSS n w=1u l=0.18u
MI8-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
M_u2 net14 B VDD VDD p w=1.37u l=0.18u
MI7 net24 A2 VDD VDD p w=1.37u l=0.18u
MI9 net14 A1 net24 VDD p w=1.37u l=0.18u
.ends
.subckt OA21D2BWP7T A1 A2 B Z VDD VSS 
MI12 net14 A2 net20 VSS n w=1u l=0.18u
MI11 net14 A1 net20 VSS n w=1u l=0.18u
MI6 net20 B VSS VSS n w=1u l=0.18u
MI8_0-M_u2 Z net14 VSS VSS n w=1u l=0.18u
MI8_1-M_u2 Z net14 VSS VSS n w=1u l=0.18u
MI8_0-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
MI8_1-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
M_u2 net14 B VDD VDD p w=1.37u l=0.18u
MI7 net24 A2 VDD VDD p w=1.37u l=0.18u
MI9 net14 A1 net24 VDD p w=1.37u l=0.18u
.ends
.subckt OA221D0BWP7T A1 A2 B1 B2 C Z VDD VSS 
MI14 net32 A2 net26 VSS n w=0.5u l=0.18u
MI7 net32 A1 net26 VSS n w=0.5u l=0.18u
MI6 net29 C VSS VSS n w=0.5u l=0.18u
M_u4 net26 B1 net29 VSS n w=0.5u l=0.18u
MI5 net26 B2 net29 VSS n w=0.5u l=0.18u
MI15-M_u2 Z net32 VSS VSS n w=0.5u l=0.18u
MI15-M_u3 Z net32 VDD VDD p w=0.685u l=0.18u
MI13 net32 A1 net43 VDD p w=0.685u l=0.18u
MI11 net32 B2 net49 VDD p w=0.685u l=0.18u
MI9 net49 B1 VDD VDD p w=0.685u l=0.18u
MI12 net43 A2 VDD VDD p w=0.685u l=0.18u
MU24 net32 C VDD VDD p w=0.685u l=0.18u
.ends
.subckt OA221D1BWP7T A1 A2 B1 B2 C Z VDD VSS 
MI14 net32 A2 net26 VSS n w=1u l=0.18u
MI7 net32 A1 net26 VSS n w=1u l=0.18u
MI6 net29 C VSS VSS n w=1u l=0.18u
M_u4 net26 B1 net29 VSS n w=1u l=0.18u
MI5 net26 B2 net29 VSS n w=1u l=0.18u
MI15-M_u2 Z net32 VSS VSS n w=1u l=0.18u
MI15-M_u3 Z net32 VDD VDD p w=1.37u l=0.18u
MI13 net32 A1 net43 VDD p w=1.37u l=0.18u
MI11 net32 B2 net49 VDD p w=1.37u l=0.18u
MI9 net49 B1 VDD VDD p w=1.225u l=0.18u
MI12 net43 A2 VDD VDD p w=1.37u l=0.18u
MU24 net32 C VDD VDD p w=1.225u l=0.18u
.ends
.subckt OA221D2BWP7T A1 A2 B1 B2 C Z VDD VSS 
MI14 net32 A2 net26 VSS n w=1u l=0.18u
MI7 net32 A1 net26 VSS n w=1u l=0.18u
MI6 net29 C VSS VSS n w=1u l=0.18u
M_u4 net26 B1 net29 VSS n w=1u l=0.18u
MI5 net26 B2 net29 VSS n w=1u l=0.18u
MI15_0-M_u2 Z net32 VSS VSS n w=1u l=0.18u
MI15_1-M_u2 Z net32 VSS VSS n w=1u l=0.18u
MI15_0-M_u3 Z net32 VDD VDD p w=1.37u l=0.18u
MI15_1-M_u3 Z net32 VDD VDD p w=1.37u l=0.18u
MI13 net32 A1 net43 VDD p w=1.37u l=0.18u
MI11 net32 B2 net49 VDD p w=1.37u l=0.18u
MI9 net49 B1 VDD VDD p w=1.37u l=0.18u
MI12 net43 A2 VDD VDD p w=1.37u l=0.18u
MU24 net32 C VDD VDD p w=1.37u l=0.18u
.ends
.subckt OA222D0BWP7T A1 A2 B1 B2 C1 C2 Z VDD VSS 
MI18 net36 A2 net27 VSS n w=0.5u l=0.18u
MI14 net39 C2 VSS VSS n w=0.5u l=0.18u
MI15 net27 B1 net39 VSS n w=0.5u l=0.18u
MI16 net27 B2 net39 VSS n w=0.5u l=0.18u
MI17 net36 A1 net27 VSS n w=0.5u l=0.18u
MU25 net39 C1 VSS VSS n w=0.5u l=0.18u
MI19-M_u2 Z net36 VSS VSS n w=0.5u l=0.18u
MI19-M_u3 Z net36 VDD VDD p w=0.685u l=0.18u
MI8 net36 C2 net46 VDD p w=0.685u l=0.18u
MI2 net46 C1 VDD VDD p w=0.685u l=0.18u
MI13 net36 A1 net34 VDD p w=0.685u l=0.18u
MI12 net34 A2 VDD VDD p w=0.685u l=0.18u
MI9 net36 B2 net37 VDD p w=0.685u l=0.18u
MI11 net37 B1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt OA222D1BWP7T A1 A2 B1 B2 C1 C2 Z VDD VSS 
MI18 net36 A2 net27 VSS n w=1u l=0.18u
MI14 net39 C2 VSS VSS n w=1u l=0.18u
MI15 net27 B1 net39 VSS n w=1u l=0.18u
MI16 net27 B2 net39 VSS n w=1u l=0.18u
MI17 net36 A1 net27 VSS n w=1u l=0.18u
MU25 net39 C1 VSS VSS n w=1u l=0.18u
MI19-M_u2 Z net36 VSS VSS n w=1u l=0.18u
MI19-M_u3 Z net36 VDD VDD p w=1.37u l=0.18u
MI8 net36 C2 net46 VDD p w=1.37u l=0.18u
MI2 net46 C1 VDD VDD p w=1.37u l=0.18u
MI13 net36 A1 net34 VDD p w=1.37u l=0.18u
MI12 net34 A2 VDD VDD p w=1.37u l=0.18u
MI9 net36 B2 net37 VDD p w=1.37u l=0.18u
MI11 net37 B1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OA222D2BWP7T A1 A2 B1 B2 C1 C2 Z VDD VSS 
MI18 net36 A2 net27 VSS n w=1u l=0.18u
MI14 net39 C2 VSS VSS n w=1u l=0.18u
MI15 net27 B1 net39 VSS n w=1u l=0.18u
MI16 net27 B2 net39 VSS n w=1u l=0.18u
MI17 net36 A1 net27 VSS n w=1u l=0.18u
MU25 net39 C1 VSS VSS n w=1u l=0.18u
MI19_0-M_u2 Z net36 VSS VSS n w=1u l=0.18u
MI19_1-M_u2 Z net36 VSS VSS n w=1u l=0.18u
MI19_0-M_u3 Z net36 VDD VDD p w=1.37u l=0.18u
MI19_1-M_u3 Z net36 VDD VDD p w=1.37u l=0.18u
MI8 net36 C2 net46 VDD p w=1.37u l=0.18u
MI2 net46 C1 VDD VDD p w=1.37u l=0.18u
MI13 net36 A1 net34 VDD p w=1.37u l=0.18u
MI12 net34 A2 VDD VDD p w=1.37u l=0.18u
MI9 net36 B2 net37 VDD p w=1.37u l=0.18u
MI11 net37 B1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OA22D0BWP7T A1 A2 B1 B2 Z VDD VSS 
M_u4 net29 B2 VSS VSS n w=0.5u l=0.18u
MI13 net30 A2 net29 VSS n w=0.5u l=0.18u
MI14 net30 A1 net29 VSS n w=0.5u l=0.18u
MI12 net29 B1 VSS VSS n w=0.5u l=0.18u
MU1-M_u2 Z net30 VSS VSS n w=0.5u l=0.18u
MU1-M_u3 Z net30 VDD VDD p w=0.685u l=0.18u
MU24 net25 B2 VDD VDD p w=0.685u l=0.18u
MI11 net22 A2 VDD VDD p w=0.685u l=0.18u
MI8 net30 B1 net25 VDD p w=0.685u l=0.18u
MI9 net30 A1 net22 VDD p w=0.685u l=0.18u
.ends
.subckt OA22D1BWP7T A1 A2 B1 B2 Z VDD VSS 
M_u4 net29 B2 VSS VSS n w=1u l=0.18u
MI13 net30 A2 net29 VSS n w=1u l=0.18u
MI14 net30 A1 net29 VSS n w=1u l=0.18u
MI12 net29 B1 VSS VSS n w=1u l=0.18u
MU1-M_u2 Z net30 VSS VSS n w=1u l=0.18u
MU1-M_u3 Z net30 VDD VDD p w=1.37u l=0.18u
MU24 net25 B2 VDD VDD p w=1.37u l=0.18u
MI11 net22 A2 VDD VDD p w=1.37u l=0.18u
MI8 net30 B1 net25 VDD p w=1.37u l=0.18u
MI9 net30 A1 net22 VDD p w=1.37u l=0.18u
.ends
.subckt OA22D2BWP7T A1 A2 B1 B2 Z VDD VSS 
M_u4 net29 B2 VSS VSS n w=1u l=0.18u
MI13 net30 A2 net29 VSS n w=1u l=0.18u
MI14 net30 A1 net29 VSS n w=1u l=0.18u
MI12 net29 B1 VSS VSS n w=1u l=0.18u
MU1_0-M_u2 Z net30 VSS VSS n w=1u l=0.18u
MU1_1-M_u2 Z net30 VSS VSS n w=1u l=0.18u
MU1_0-M_u3 Z net30 VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 Z net30 VDD VDD p w=1.37u l=0.18u
MU24 net25 B2 VDD VDD p w=1.37u l=0.18u
MI11 net22 A2 VDD VDD p w=1.37u l=0.18u
MI8 net30 B1 net25 VDD p w=1.37u l=0.18u
MI9 net30 A1 net22 VDD p w=1.37u l=0.18u
.ends
.subckt OA31D0BWP7T A1 A2 A3 B Z VDD VSS 
M_u5 VSS B net22 VSS n w=0.5u l=0.18u
MI8 net22 A3 net30 VSS n w=0.5u l=0.18u
MI7 net22 A2 net30 VSS n w=0.5u l=0.18u
MI6 net22 A1 net30 VSS n w=0.5u l=0.18u
MU1-M_u2 Z net30 VSS VSS n w=0.5u l=0.18u
MU1-M_u3 Z net30 VDD VDD p w=0.685u l=0.18u
MI3 net38 A1 VDD VDD p w=0.685u l=0.18u
MI4 net35 A2 net38 VDD p w=0.685u l=0.18u
MI5 net30 A3 net35 VDD p w=0.685u l=0.18u
M_u11 net30 B VDD VDD p w=0.685u l=0.18u
.ends
.subckt OA31D1BWP7T A1 A2 A3 B Z VDD VSS 
M_u5 VSS B net22 VSS n w=1u l=0.18u
MI8 net22 A3 net30 VSS n w=1u l=0.18u
MI7 net22 A2 net30 VSS n w=1u l=0.18u
MI6 net22 A1 net30 VSS n w=1u l=0.18u
MU1-M_u2 Z net30 VSS VSS n w=1u l=0.18u
MU1-M_u3 Z net30 VDD VDD p w=1.37u l=0.18u
MI3 net38 A1 VDD VDD p w=1.37u l=0.18u
MI4 net35 A2 net38 VDD p w=1.37u l=0.18u
MI5 net30 A3 net35 VDD p w=1.37u l=0.18u
M_u11 net30 B VDD VDD p w=1.37u l=0.18u
.ends
.subckt OA31D2BWP7T A1 A2 A3 B Z VDD VSS 
M_u5 VSS B net22 VSS n w=1u l=0.18u
MI8 net22 A3 net30 VSS n w=1u l=0.18u
MI7 net22 A2 net30 VSS n w=1u l=0.18u
MI6 net22 A1 net30 VSS n w=1u l=0.18u
MU1_0-M_u2 Z net30 VSS VSS n w=1u l=0.18u
MU1_1-M_u2 Z net30 VSS VSS n w=1u l=0.18u
MU1_0-M_u3 Z net30 VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 Z net30 VDD VDD p w=1.37u l=0.18u
MI3 net38 A1 VDD VDD p w=1.37u l=0.18u
MI4 net35 A2 net38 VDD p w=1.37u l=0.18u
MI5 net30 A3 net35 VDD p w=1.37u l=0.18u
M_u11 net30 B VDD VDD p w=1.37u l=0.18u
.ends
.subckt OA32D0BWP7T A1 A2 A3 B1 B2 Z VDD VSS 
MI12 net14 B1 VSS VSS n w=0.5u l=0.18u
MI11 net14 B2 VSS VSS n w=0.5u l=0.18u
MI3 net35 A3 net14 VSS n w=0.5u l=0.18u
MI8 net35 A2 net14 VSS n w=0.5u l=0.18u
MI9 net35 A1 net14 VSS n w=0.5u l=0.18u
MU1-M_u2 Z net35 VSS VSS n w=0.465u l=0.18u
MU1-M_u3 Z net35 VDD VDD p w=0.685u l=0.18u
MI16-MI12 net35 B2 XI16-net11 VDD p w=0.685u l=0.18u
MI16-MI13 XI16-net11 B1 VDD VDD p w=0.685u l=0.18u
MI15-MI12 net35 A3 XI15-net11 VDD p w=0.685u l=0.18u
MI15-MI13 XI15-net11 A2 XI15-net18 VDD p w=0.685u l=0.18u
MI15-MI15 XI15-net18 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt OA32D1BWP7T A1 A2 A3 B1 B2 Z VDD VSS 
MI7 net14 B1 VSS VSS n w=1u l=0.18u
MI6 net14 B2 VSS VSS n w=1u l=0.18u
MI3 net35 A3 net14 VSS n w=1u l=0.18u
MI4 net35 A2 net14 VSS n w=1u l=0.18u
MI5 net35 A1 net14 VSS n w=1u l=0.18u
MU1-M_u2 Z net35 VSS VSS n w=1u l=0.18u
MU1-M_u3 Z net35 VDD VDD p w=1.37u l=0.18u
MI16-MI12 net35 B2 XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 B1 VDD VDD p w=1.37u l=0.18u
MI15-MI12 net35 A3 XI15-net11 VDD p w=1.37u l=0.18u
MI15-MI13 XI15-net11 A2 XI15-net18 VDD p w=1.37u l=0.18u
MI15-MI15 XI15-net18 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OA32D2BWP7T A1 A2 A3 B1 B2 Z VDD VSS 
MI7 net14 B1 VSS VSS n w=1u l=0.18u
MI6 net14 B2 VSS VSS n w=1u l=0.18u
MI3 net35 A3 net14 VSS n w=1u l=0.18u
MI4 net35 A2 net14 VSS n w=1u l=0.18u
MI5 net35 A1 net14 VSS n w=1u l=0.18u
MU1_0-M_u2 Z net35 VSS VSS n w=1u l=0.18u
MU1_1-M_u2 Z net35 VSS VSS n w=1u l=0.18u
MU1_0-M_u3 Z net35 VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 Z net35 VDD VDD p w=1.37u l=0.18u
MI16-MI12 net35 B2 XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 B1 VDD VDD p w=1.37u l=0.18u
MI15-MI12 net35 A3 XI15-net11 VDD p w=1.37u l=0.18u
MI15-MI13 XI15-net11 A2 XI15-net18 VDD p w=1.37u l=0.18u
MI15-MI15 XI15-net18 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OA33D0BWP7T A1 A2 A3 B1 B2 B3 Z VDD VSS 
MI5 net15 B2 VSS VSS n w=0.5u l=0.18u
MI6 net15 B1 VSS VSS n w=0.5u l=0.18u
M_u3 net37 A3 net15 VSS n w=0.5u l=0.18u
MI2 net37 A2 net15 VSS n w=0.5u l=0.18u
MI4 net15 B3 VSS VSS n w=0.5u l=0.18u
MI3 net37 A1 net15 VSS n w=0.5u l=0.18u
MU1-M_u2 Z net37 VSS VSS n w=0.5u l=0.18u
MU1-M_u3 Z net37 VDD VDD p w=0.685u l=0.18u
MI1-MI12 net37 B3 XI1-net11 VDD p w=0.685u l=0.18u
MI1-MI13 XI1-net11 B2 XI1-net18 VDD p w=0.685u l=0.18u
MI1-MI15 XI1-net18 B1 VDD VDD p w=0.685u l=0.18u
MI0-MI12 net37 A3 XI0-net11 VDD p w=0.685u l=0.18u
MI0-MI13 XI0-net11 A2 XI0-net18 VDD p w=0.685u l=0.18u
MI0-MI15 XI0-net18 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt OA33D1BWP7T A1 A2 A3 B1 B2 B3 Z VDD VSS 
MI5 net15 B2 VSS VSS n w=1u l=0.18u
MI6 net15 B1 VSS VSS n w=1u l=0.18u
M_u3 net37 A3 net15 VSS n w=1u l=0.18u
MI2 net37 A2 net15 VSS n w=1u l=0.18u
MI4 net15 B3 VSS VSS n w=1u l=0.18u
MI3 net37 A1 net15 VSS n w=1u l=0.18u
MU1-M_u2 Z net37 VSS VSS n w=1u l=0.18u
MU1-M_u3 Z net37 VDD VDD p w=1.37u l=0.18u
MI1-MI12 net37 B3 XI1-net11 VDD p w=1.37u l=0.18u
MI1-MI13 XI1-net11 B2 XI1-net18 VDD p w=1.37u l=0.18u
MI1-MI15 XI1-net18 B1 VDD VDD p w=1.37u l=0.18u
MI0-MI12 net37 A3 XI0-net11 VDD p w=1.37u l=0.18u
MI0-MI13 XI0-net11 A2 XI0-net18 VDD p w=1.37u l=0.18u
MI0-MI15 XI0-net18 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OA33D2BWP7T A1 A2 A3 B1 B2 B3 Z VDD VSS 
MI5 net15 B2 VSS VSS n w=1u l=0.18u
MI6 net15 B1 VSS VSS n w=1u l=0.18u
M_u3 net37 A3 net15 VSS n w=1u l=0.18u
MI2 net37 A2 net15 VSS n w=1u l=0.18u
MI4 net15 B3 VSS VSS n w=1u l=0.18u
MI3 net37 A1 net15 VSS n w=1u l=0.18u
MU1_0-M_u2 Z net37 VSS VSS n w=1u l=0.18u
MU1_1-M_u2 Z net37 VSS VSS n w=1u l=0.18u
MU1_0-M_u3 Z net37 VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 Z net37 VDD VDD p w=1.37u l=0.18u
MI1-MI12 net37 B3 XI1-net11 VDD p w=1.37u l=0.18u
MI1-MI13 XI1-net11 B2 XI1-net18 VDD p w=1.37u l=0.18u
MI1-MI15 XI1-net18 B1 VDD VDD p w=1.37u l=0.18u
MI0-MI12 net37 A3 XI0-net11 VDD p w=1.37u l=0.18u
MI0-MI13 XI0-net11 A2 XI0-net18 VDD p w=1.37u l=0.18u
MI0-MI15 XI0-net18 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OAI211D0BWP7T A1 A2 B C ZN VDD VSS 
MI8 net36 B net24 VSS n w=0.5u l=0.18u
MI9 net24 C VSS VSS n w=0.5u l=0.18u
M_u2 ZN A1 net36 VSS n w=0.5u l=0.18u
MI7 ZN A2 net36 VSS n w=0.5u l=0.18u
MI6 ZN A2 net35 VDD p w=0.685u l=0.18u
MI5 net35 A1 VDD VDD p w=0.685u l=0.18u
MI4 ZN C VDD VDD p w=0.685u l=0.18u
M_u12 ZN B VDD VDD p w=0.685u l=0.18u
.ends
.subckt OAI211D1BWP7T A1 A2 B C ZN VDD VSS 
MI2 net36 B net24 VSS n w=1u l=0.18u
MI3 net24 C VSS VSS n w=1u l=0.18u
M_u2 ZN A1 net36 VSS n w=1u l=0.18u
M_u3 ZN A2 net36 VSS n w=1u l=0.18u
MI1 ZN A2 net35 VDD p w=1.37u l=0.18u
MI0 net35 A1 VDD VDD p w=1.37u l=0.18u
M_u11 ZN C VDD VDD p w=1.37u l=0.18u
M_u12 ZN B VDD VDD p w=1.37u l=0.18u
.ends
.subckt OAI211D2BWP7T A1 A2 B C ZN VDD VSS 
MI8_0 net36 B net_026[0] VSS n w=1u l=0.18u
MI8_1 net36 B net_026[1] VSS n w=1u l=0.18u
MI11_0 net_026[0] C VSS VSS n w=1u l=0.18u
MI11_1 net_026[1] C VSS VSS n w=1u l=0.18u
M_u2 ZN A1 net36 VSS n w=2u l=0.18u
MI7 ZN A2 net36 VSS n w=2u l=0.18u
MI12 ZN A2 net38 VDD p w=1.37u l=0.18u
MI5 net38 A1 VDD VDD p w=1.37u l=0.18u
MI13 ZN A2 net040 VDD p w=1.37u l=0.18u
MI14 net040 A1 VDD VDD p w=1.37u l=0.18u
MI4 ZN C VDD VDD p w=2.74u l=0.18u
M_u12 ZN B VDD VDD p w=2.74u l=0.18u
.ends
.subckt OAI21D0BWP7T A1 A2 B ZN VDD VSS 
MI0 net15 B VSS VSS n w=0.465u l=0.18u
M_u2 ZN A1 net15 VSS n w=0.5u l=0.18u
M_u3 ZN A2 net15 VSS n w=0.5u l=0.18u
M_u9 ZN B VDD VDD p w=0.685u l=0.18u
MI16-MI12 ZN A1 XI16-net11 VDD p w=0.685u l=0.18u
MI16-MI13 XI16-net11 A2 VDD VDD p w=0.685u l=0.18u
.ends
.subckt OAI21D1BWP7T A1 A2 B ZN VDD VSS 
M_u2 ZN A1 net15 VSS n w=1u l=0.18u
M_u3 ZN A2 net15 VSS n w=1u l=0.18u
M_u4 net15 B VSS VSS n w=1u l=0.18u
M_u9 ZN B VDD VDD p w=1.37u l=0.18u
MI16-MI12 ZN A1 XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OAI21D2BWP7T A1 A2 B ZN VDD VSS 
M_u2 ZN A1 net15 VSS n w=2u l=0.18u
M_u3 ZN A2 net15 VSS n w=2u l=0.18u
M_u4 net15 B VSS VSS n w=2u l=0.18u
M_u9 ZN B VDD VDD p w=2.74u l=0.18u
MI16_0-MI12 ZN A1 XI16_0-net11 VDD p w=1.37u l=0.18u
MI16_0-MI13 XI16_0-net11 A2 VDD VDD p w=1.37u l=0.18u
MI16_1-MI12 ZN A1 XI16_1-net11 VDD p w=1.37u l=0.18u
MI16_1-MI13 XI16_1-net11 A2 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OAI221D0BWP7T A1 A2 B1 B2 C ZN VDD VSS 
MI14 ZN A2 net26 VSS n w=0.5u l=0.18u
MI7 ZN A1 net26 VSS n w=0.5u l=0.18u
MI6 net29 C VSS VSS n w=0.5u l=0.18u
M_u4 net26 B1 net29 VSS n w=0.5u l=0.18u
MI5 net26 B2 net29 VSS n w=0.5u l=0.18u
MI13 ZN A1 net43 VDD p w=0.685u l=0.18u
MI11 ZN B2 net49 VDD p w=0.685u l=0.18u
MI9 net49 B1 VDD VDD p w=0.685u l=0.18u
MI12 net43 A2 VDD VDD p w=0.685u l=0.18u
MU24 ZN C VDD VDD p w=0.685u l=0.18u
.ends
.subckt OAI221D1BWP7T A1 A2 B1 B2 C ZN VDD VSS 
M_u2 ZN A1 net26 VSS n w=1u l=0.18u
M_u3 ZN A2 net26 VSS n w=1u l=0.18u
M_u5 net26 B2 net29 VSS n w=1u l=0.18u
M_u4 net26 B1 net29 VSS n w=1u l=0.18u
MU23 net29 C VSS VSS n w=1u l=0.18u
MI2 ZN B2 net49 VDD p w=1.37u l=0.18u
MI3 net43 A2 VDD VDD p w=1.37u l=0.18u
MI4 ZN A1 net43 VDD p w=1.37u l=0.18u
MI1 net49 B1 VDD VDD p w=1.37u l=0.18u
MU24 ZN C VDD VDD p w=1.37u l=0.18u
.ends
.subckt OAI221D2BWP7T A1 A2 B1 B2 C ZN VDD VSS 
MI14 ZN A2 net26 VSS n w=2u l=0.18u
MI7 ZN A1 net26 VSS n w=2u l=0.18u
MI6 net29 C VSS VSS n w=2u l=0.18u
M_u4 net26 B1 net29 VSS n w=2u l=0.18u
MI5 net26 B2 net29 VSS n w=2u l=0.18u
MI17_0 net49[0] A2 VDD VDD p w=1.37u l=0.18u
MI17_1 net49[1] A2 VDD VDD p w=1.37u l=0.18u
MI15_0 ZN B2 net52[0] VDD p w=1.37u l=0.18u
MI15_1 ZN B2 net52[1] VDD p w=1.37u l=0.18u
MI9_0 net52[0] B1 VDD VDD p w=1.37u l=0.18u
MI9_1 net52[1] B1 VDD VDD p w=1.37u l=0.18u
MI16_0 ZN A1 net49[0] VDD p w=1.37u l=0.18u
MI16_1 ZN A1 net49[1] VDD p w=1.37u l=0.18u
MU24 ZN C VDD VDD p w=2.74u l=0.18u
.ends
.subckt OAI222D0BWP7T A1 A2 B1 B2 C1 C2 ZN VDD VSS 
MI18 ZN A2 net27 VSS n w=0.5u l=0.18u
MI14 net39 C2 VSS VSS n w=0.5u l=0.18u
MI15 net27 B1 net39 VSS n w=0.5u l=0.18u
MI16 net27 B2 net39 VSS n w=0.5u l=0.18u
MI17 ZN A1 net27 VSS n w=0.5u l=0.18u
MU25 net39 C1 VSS VSS n w=0.5u l=0.18u
MI8 ZN C2 net46 VDD p w=0.685u l=0.18u
MI2 net46 C1 VDD VDD p w=0.685u l=0.18u
MI13 ZN A1 net34 VDD p w=0.685u l=0.18u
MI12 net34 A2 VDD VDD p w=0.685u l=0.18u
MI9 ZN B2 net37 VDD p w=0.685u l=0.18u
MI11 net37 B1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt OAI222D1BWP7T A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_u3 ZN A2 net27 VSS n w=1u l=0.18u
M_u2 ZN A1 net27 VSS n w=1u l=0.18u
MU25 net39 C1 VSS VSS n w=1u l=0.18u
MU23 net39 C2 VSS VSS n w=1u l=0.18u
M_u5 net27 B2 net39 VSS n w=1u l=0.18u
M_u4 net27 B1 net39 VSS n w=1u l=0.18u
MI4 net37 B1 VDD VDD p w=1.25u l=0.18u
MI5 ZN B2 net37 VDD p w=1.37u l=0.18u
MI6 ZN A1 net34 VDD p w=1.295u l=0.18u
MI7 net34 A2 VDD VDD p w=1.25u l=0.18u
MI2 net46 C1 VDD VDD p w=1.37u l=0.18u
MI3 ZN C2 net46 VDD p w=1.37u l=0.18u
.ends
.subckt OAI222D2BWP7T A1 A2 B1 B2 C1 C2 ZN VDD VSS 
MI18 ZN A2 net27 VSS n w=2u l=0.18u
MI14 net39 C2 VSS VSS n w=2u l=0.18u
MI15 net27 B1 net39 VSS n w=2u l=0.18u
MI16 net27 B2 net39 VSS n w=2u l=0.18u
MI17 ZN A1 net27 VSS n w=2u l=0.18u
MU25 net39 C1 VSS VSS n w=2u l=0.18u
MI23_0 ZN A1 net53[0] VDD p w=1.37u l=0.18u
MI23_1 ZN A1 net53[1] VDD p w=1.37u l=0.18u
MI2_0 net65[0] C1 VDD VDD p w=1.37u l=0.18u
MI2_1 net65[1] C1 VDD VDD p w=1.37u l=0.18u
MI22_0 net53[0] A2 VDD VDD p w=1.37u l=0.18u
MI22_1 net53[1] A2 VDD VDD p w=1.37u l=0.18u
MI21_0 ZN B2 net59[0] VDD p w=1.37u l=0.18u
MI21_1 ZN B2 net59[1] VDD p w=1.37u l=0.18u
MI19_0 ZN C2 net65[0] VDD p w=1.37u l=0.18u
MI19_1 ZN C2 net65[1] VDD p w=1.37u l=0.18u
MI20_0 net59[0] B1 VDD VDD p w=1.37u l=0.18u
MI20_1 net59[1] B1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OAI22D0BWP7T A1 A2 B1 B2 ZN VDD VSS 
MI9 ZN A1 net10 VSS n w=0.5u l=0.18u
M_u4 net10 B2 VSS VSS n w=0.5u l=0.18u
MI8 ZN A2 net10 VSS n w=0.5u l=0.18u
MI7 net10 B1 VSS VSS n w=0.5u l=0.18u
MU24 net30 B2 VDD VDD p w=0.685u l=0.18u
MI6 ZN A1 net24 VDD p w=0.685u l=0.18u
MI5 net24 A2 VDD VDD p w=0.685u l=0.18u
MI4 ZN B1 net30 VDD p w=0.685u l=0.18u
.ends
.subckt OAI22D1BWP7T A1 A2 B1 B2 ZN VDD VSS 
M_u4 net10 B2 VSS VSS n w=1u l=0.18u
M_u3 ZN A1 net10 VSS n w=1u l=0.18u
M_u2 ZN A2 net10 VSS n w=1u l=0.18u
M_u5 net10 B1 VSS VSS n w=1u l=0.18u
MU24 net30 B2 VDD VDD p w=1.37u l=0.18u
MI3 ZN A1 net24 VDD p w=1.37u l=0.18u
MI2 net24 A2 VDD VDD p w=1.37u l=0.18u
MI1 ZN B1 net30 VDD p w=1.37u l=0.18u
.ends
.subckt OAI22D2BWP7T A1 A2 B1 B2 ZN VDD VSS 
M_u4 net10 B2 VSS VSS n w=2u l=0.18u
M_u3 ZN A1 net10 VSS n w=2u l=0.18u
M_u2 ZN A2 net10 VSS n w=2u l=0.18u
M_u5 net10 B1 VSS VSS n w=2u l=0.18u
MU24_0 net45[0] B2 VDD VDD p w=1.37u l=0.18u
MU24_1 net45[1] B2 VDD VDD p w=1.37u l=0.18u
MI6_0 net42[0] A2 VDD VDD p w=1.37u l=0.18u
MI6_1 net42[1] A2 VDD VDD p w=1.37u l=0.18u
MI5_0 ZN A1 net42[0] VDD p w=1.37u l=0.18u
MI5_1 ZN A1 net42[1] VDD p w=1.37u l=0.18u
MI4_0 ZN B1 net45[0] VDD p w=1.37u l=0.18u
MI4_1 ZN B1 net45[1] VDD p w=1.37u l=0.18u
.ends
.subckt OAI31D0BWP7T A1 A2 A3 B ZN VDD VSS 
M_u5 VSS B net22 VSS n w=0.5u l=0.18u
MI8 net22 A3 ZN VSS n w=0.5u l=0.18u
MI7 net22 A2 ZN VSS n w=0.5u l=0.18u
MI6 net22 A1 ZN VSS n w=0.5u l=0.18u
MI3 net38 A1 VDD VDD p w=0.685u l=0.18u
MI4 net35 A2 net38 VDD p w=0.685u l=0.18u
MI5 ZN A3 net35 VDD p w=0.685u l=0.18u
M_u11 ZN B VDD VDD p w=0.685u l=0.18u
.ends
.subckt OAI31D1BWP7T A1 A2 A3 B ZN VDD VSS 
M_u5 VSS B net22 VSS n w=1u l=0.18u
M_u3 ZN A3 net22 VSS n w=1u l=0.18u
M_u2 ZN A2 net22 VSS n w=1u l=0.18u
MU21 ZN A1 net22 VSS n w=1u l=0.18u
MI0 net38 A1 VDD VDD p w=1.37u l=0.18u
MI1 net35 A2 net38 VDD p w=1.37u l=0.18u
MI2 ZN A3 net35 VDD p w=1.37u l=0.18u
M_u11 ZN B VDD VDD p w=1.37u l=0.18u
.ends
.subckt OAI31D2BWP7T A1 A2 A3 B ZN VDD VSS 
M_u5 VSS B net22 VSS n w=1.86u l=0.18u
MI8 net22 A3 ZN VSS n w=1.86u l=0.18u
MI7 net22 A2 ZN VSS n w=1.86u l=0.18u
MI6 net22 A1 ZN VSS n w=1.86u l=0.18u
MI3 net041 A1 VDD VDD p w=1.37u l=0.18u
MI9 net044 A2 net041 VDD p w=1.25u l=0.18u
MI11 ZN A3 net044 VDD p w=1.305u l=0.18u
MI12 net023 A1 VDD VDD p w=1.25u l=0.18u
MI13 net038 A2 net023 VDD p w=1.25u l=0.18u
MI14 ZN A3 net038 VDD p w=1.305u l=0.18u
M_u11 ZN B VDD VDD p w=2.74u l=0.18u
.ends
.subckt OAI32D0BWP7T A1 A2 A3 B1 B2 ZN VDD VSS 
MI7 net14 B1 VSS VSS n w=0.5u l=0.18u
MI6 net14 B2 VSS VSS n w=0.5u l=0.18u
MI3 ZN A3 net14 VSS n w=0.5u l=0.18u
MI4 ZN A2 net14 VSS n w=0.5u l=0.18u
MI5 ZN A1 net14 VSS n w=0.5u l=0.18u
MI16-MI12 ZN B2 XI16-net11 VDD p w=0.685u l=0.18u
MI16-MI13 XI16-net11 B1 VDD VDD p w=0.685u l=0.18u
MI15-MI12 ZN A3 XI15-net11 VDD p w=0.685u l=0.18u
MI15-MI13 XI15-net11 A2 XI15-net18 VDD p w=0.685u l=0.18u
MI15-MI15 XI15-net18 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt OAI32D1BWP7T A1 A2 A3 B1 B2 ZN VDD VSS 
MI0 net14 B2 VSS VSS n w=1u l=0.18u
MI3 ZN A3 net14 VSS n w=1u l=0.18u
MI2 ZN A2 net14 VSS n w=1u l=0.18u
M_u4 net14 B1 VSS VSS n w=1u l=0.18u
MI1 ZN A1 net14 VSS n w=1u l=0.18u
MI16-MI12 ZN B2 XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 B1 VDD VDD p w=1.37u l=0.18u
MI15-MI12 ZN A3 XI15-net11 VDD p w=1.37u l=0.18u
MI15-MI13 XI15-net11 A2 XI15-net18 VDD p w=1.37u l=0.18u
MI15-MI15 XI15-net18 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OAI32D2BWP7T A1 A2 A3 B1 B2 ZN VDD VSS 
MI0 net14 B2 VSS VSS n w=2u l=0.18u
MI3 ZN A3 net14 VSS n w=2u l=0.18u
MI2 ZN A2 net14 VSS n w=2u l=0.18u
M_u4 net14 B1 VSS VSS n w=2u l=0.18u
MI1 ZN A1 net14 VSS n w=2u l=0.18u
MI16-MI12 ZN B2 XI16-net11 VDD p w=1.37u l=0.18u
MI16-MI13 XI16-net11 B1 VDD VDD p w=1.37u l=0.18u
MI4-MI12 ZN B2 XI4-net11 VDD p w=1.37u l=0.18u
MI4-MI13 XI4-net11 B1 VDD VDD p w=1.37u l=0.18u
MI5 ZN A3 net028 VDD p w=1.37u l=0.18u
MI6 net028 A2 net031 VDD p w=1.37u l=0.18u
MI7 net031 A1 VDD VDD p w=1.37u l=0.18u
MI12 ZN A3 net028 VDD p w=1.37u l=0.18u
MI13 net028 A2 net031 VDD p w=1.37u l=0.18u
MI15 net031 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OAI33D0BWP7T A1 A2 A3 B1 B2 B3 ZN VDD VSS 
MI5 net15 B2 VSS VSS n w=0.5u l=0.18u
MI6 net15 B1 VSS VSS n w=0.5u l=0.18u
M_u3 ZN A3 net15 VSS n w=0.5u l=0.18u
MI2 ZN A2 net15 VSS n w=0.5u l=0.18u
MI4 net15 B3 VSS VSS n w=0.5u l=0.18u
MI3 ZN A1 net15 VSS n w=0.5u l=0.18u
MI1-MI12 ZN B3 XI1-net11 VDD p w=0.685u l=0.18u
MI1-MI13 XI1-net11 B2 XI1-net18 VDD p w=0.685u l=0.18u
MI1-MI15 XI1-net18 B1 VDD VDD p w=0.685u l=0.18u
MI0-MI12 ZN A3 XI0-net11 VDD p w=0.685u l=0.18u
MI0-MI13 XI0-net11 A2 XI0-net18 VDD p w=0.685u l=0.18u
MI0-MI15 XI0-net18 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt OAI33D1BWP7T A1 A2 A3 B1 B2 B3 ZN VDD VSS 
MI7 net15 B2 VSS VSS n w=1u l=0.18u
MI8 net15 B1 VSS VSS n w=1u l=0.18u
MI4 ZN A2 net15 VSS n w=1u l=0.18u
MI5 ZN A3 net15 VSS n w=1u l=0.18u
MI6 net15 B3 VSS VSS n w=1u l=0.18u
MU21 ZN A1 net15 VSS n w=1u l=0.18u
MI2-MI12 ZN B3 XI2-net11 VDD p w=1.37u l=0.18u
MI2-MI13 XI2-net11 B2 XI2-net18 VDD p w=1.37u l=0.18u
MI2-MI15 XI2-net18 B1 VDD VDD p w=1.37u l=0.18u
MI3-MI12 ZN A3 XI3-net11 VDD p w=1.37u l=0.18u
MI3-MI13 XI3-net11 A2 XI3-net18 VDD p w=1.37u l=0.18u
MI3-MI15 XI3-net18 A1 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OAI33D2BWP7T A1 A2 A3 B1 B2 B3 ZN VDD VSS 
MI7 net15 B2 VSS VSS n w=1.9u l=0.18u
MI8 net15 B1 VSS VSS n w=1.9u l=0.18u
MI4 ZN A2 net15 VSS n w=1.9u l=0.18u
MI5 ZN A3 net15 VSS n w=1.9u l=0.18u
MI6 net15 B3 VSS VSS n w=1.9u l=0.18u
MU21 ZN A1 net15 VSS n w=1.9u l=0.18u
MI11-MI12 ZN B3 XI11-net11 VDD p w=1.23u l=0.18u
MI11-MI13 XI11-net11 B2 XI11-net18 VDD p w=1.23u l=0.18u
MI11-MI15 XI11-net18 B1 VDD VDD p w=1.23u l=0.18u
MI12-MI12 ZN A3 XI12-net11 VDD p w=1.23u l=0.18u
MI12-MI13 XI12-net11 A2 XI12-net18 VDD p w=1.23u l=0.18u
MI12-MI15 XI12-net18 A1 VDD VDD p w=1.23u l=0.18u
MI13-MI12 ZN B3 XI13-net11 VDD p w=1.23u l=0.18u
MI13-MI13 XI13-net11 B2 XI13-net18 VDD p w=1.23u l=0.18u
MI13-MI15 XI13-net18 B1 VDD VDD p w=1.23u l=0.18u
MI3-MI12 ZN A3 XI3-net11 VDD p w=1.23u l=0.18u
MI3-MI13 XI3-net11 A2 XI3-net18 VDD p w=1.23u l=0.18u
MI3-MI15 XI3-net18 A1 VDD VDD p w=1.23u l=0.18u
.ends
.subckt OR2D0BWP7T A1 A2 Z VDD VSS 
MU1-M_u2 Z net7 VSS VSS n w=0.5u l=0.18u
M_u7-M_u4 net7 A1 VSS VSS n w=0.5u l=0.18u
M_u7-M_u3 net7 A2 VSS VSS n w=0.5u l=0.18u
MU1-M_u3 Z net7 VDD VDD p w=0.685u l=0.18u
M_u7-M_u1 X_u7-net8 A2 VDD VDD p w=0.685u l=0.18u
M_u7-M_u2 net7 A1 X_u7-net8 VDD p w=0.685u l=0.18u
.ends
.subckt OR2D1BWP7T A1 A2 Z VDD VSS 
MU1-M_u2 Z net7 VSS VSS n w=1u l=0.18u
M_u7-M_u4 net7 A1 VSS VSS n w=0.5u l=0.18u
M_u7-M_u3 net7 A2 VSS VSS n w=0.5u l=0.18u
MU1-M_u3 Z net7 VDD VDD p w=1.37u l=0.18u
M_u7-M_u1 X_u7-net8 A2 VDD VDD p w=1.37u l=0.18u
M_u7-M_u2 net7 A1 X_u7-net8 VDD p w=1.37u l=0.18u
.ends
.subckt OR2D2BWP7T A1 A2 Z VDD VSS 
MU1_0-M_u2 Z net9 VSS VSS n w=1u l=0.18u
MU1_1-M_u2 Z net9 VSS VSS n w=1u l=0.18u
M_u7-M_u4 net9 A1 VSS VSS n w=0.5u l=0.18u
M_u7-M_u3 net9 A2 VSS VSS n w=0.5u l=0.18u
MU1_0-M_u3 Z net9 VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 Z net9 VDD VDD p w=1.37u l=0.18u
M_u7-M_u1 X_u7-net8 A2 VDD VDD p w=1.37u l=0.18u
M_u7-M_u2 net9 A1 X_u7-net8 VDD p w=1.37u l=0.18u
.ends
.subckt OR2D4BWP7T A1 A2 Z VDD VSS 
MU1_0-M_u2 Z p0 VSS VSS n w=1u l=0.18u
MU1_1-M_u2 Z p0 VSS VSS n w=1u l=0.18u
MU1_2-M_u2 Z p0 VSS VSS n w=1u l=0.18u
MU1_3-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u7_0-M_u4 p0 A1 VSS VSS n w=0.5u l=0.18u
M_u7_0-M_u3 p0 A2 VSS VSS n w=0.5u l=0.18u
M_u7_1-M_u4 p0 A1 VSS VSS n w=0.5u l=0.18u
M_u7_1-M_u3 p0 A2 VSS VSS n w=0.5u l=0.18u
MU1_0-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
MU1_2-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
MU1_3-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u7_0-M_u1 X_u7_0-net8 A2 VDD VDD p w=1.37u l=0.18u
M_u7_0-M_u2 p0 A1 X_u7_0-net8 VDD p w=1.37u l=0.18u
M_u7_1-M_u1 X_u7_1-net8 A2 VDD VDD p w=1.37u l=0.18u
M_u7_1-M_u2 p0 A1 X_u7_1-net8 VDD p w=1.37u l=0.18u
.ends
.subckt OR2D8BWP7T A1 A2 Z VDD VSS 
MU1_0-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU1_1-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU1_2-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU1_3-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU1_4-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU1_5-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU1_6-M_u2 Z n0 VSS VSS n w=1u l=0.18u
MU1_7-M_u2 Z n0 VSS VSS n w=1u l=0.18u
M_u7_0-M_u4 n0 A1 VSS VSS n w=0.5u l=0.18u
M_u7_0-M_u3 n0 A2 VSS VSS n w=0.5u l=0.18u
M_u7_1-M_u4 n0 A1 VSS VSS n w=0.5u l=0.18u
M_u7_1-M_u3 n0 A2 VSS VSS n w=0.5u l=0.18u
M_u7_2-M_u4 n0 A1 VSS VSS n w=0.5u l=0.18u
M_u7_2-M_u3 n0 A2 VSS VSS n w=0.5u l=0.18u
MU1_0-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU1_1-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU1_2-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU1_3-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU1_4-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU1_5-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU1_6-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
MU1_7-M_u3 Z n0 VDD VDD p w=1.37u l=0.18u
M_u7_0-M_u1 X_u7_0-net8 A2 VDD VDD p w=1.37u l=0.18u
M_u7_0-M_u2 n0 A1 X_u7_0-net8 VDD p w=1.37u l=0.18u
M_u7_1-M_u1 X_u7_1-net8 A2 VDD VDD p w=1.37u l=0.18u
M_u7_1-M_u2 n0 A1 X_u7_1-net8 VDD p w=1.37u l=0.18u
M_u7_2-M_u1 X_u7_2-net8 A2 VDD VDD p w=1.37u l=0.18u
M_u7_2-M_u2 n0 A1 X_u7_2-net8 VDD p w=1.37u l=0.18u
.ends
.subckt OR2XD1BWP7T A1 A2 Z VDD VSS 
MU1-M_u2 Z net7 VSS VSS n w=1u l=0.18u
M_u7-M_u4 net7 A1 VSS VSS n w=1u l=0.18u
M_u7-M_u3 net7 A2 VSS VSS n w=1u l=0.18u
MU1-M_u3 Z net7 VDD VDD p w=1.37u l=0.18u
M_u7-M_u1 X_u7-net8 A2 VDD VDD p w=1.37u l=0.18u
M_u7-M_u2 net7 A1 X_u7-net8 VDD p w=1.37u l=0.18u
.ends
.subckt OR3D0BWP7T A1 A2 A3 Z VDD VSS 
MU42-M_u6 net7 A3 VSS VSS n w=0.5u l=0.18u
MU42-M_u5 net7 A2 VSS VSS n w=0.5u l=0.18u
MU42-M_u4 net7 A1 VSS VSS n w=0.5u l=0.18u
M_u4-M_u2 Z net7 VSS VSS n w=0.5u l=0.18u
MU42-M_u1 XU42-net9 A1 VDD VDD p w=0.685u l=0.18u
MU42-M_u2 XU42-net12 A2 XU42-net9 VDD p w=0.685u l=0.18u
MU42-M_u3 net7 A3 XU42-net12 VDD p w=0.685u l=0.18u
M_u4-M_u3 Z net7 VDD VDD p w=0.685u l=0.18u
.ends
.subckt OR3D1BWP7T A1 A2 A3 Z VDD VSS 
MU42-M_u6 net7 A3 VSS VSS n w=0.5u l=0.18u
MU42-M_u5 net7 A2 VSS VSS n w=0.5u l=0.18u
MU42-M_u4 net7 A1 VSS VSS n w=0.5u l=0.18u
M_u4-M_u2 Z net7 VSS VSS n w=1u l=0.18u
MU42-M_u1 XU42-net9 A1 VDD VDD p w=1.37u l=0.18u
MU42-M_u2 XU42-net12 A2 XU42-net9 VDD p w=1.37u l=0.18u
MU42-M_u3 net7 A3 XU42-net12 VDD p w=1.37u l=0.18u
M_u4-M_u3 Z net7 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OR3D2BWP7T A1 A2 A3 Z VDD VSS 
MU42-M_u6 net12 A3 VSS VSS n w=0.5u l=0.18u
MU42-M_u5 net12 A2 VSS VSS n w=0.5u l=0.18u
MU42-M_u4 net12 A1 VSS VSS n w=0.5u l=0.18u
M_u4_0-M_u2 Z net12 VSS VSS n w=1u l=0.18u
M_u4_1-M_u2 Z net12 VSS VSS n w=1u l=0.18u
MU42-M_u1 XU42-net9 A1 VDD VDD p w=1.37u l=0.18u
MU42-M_u2 XU42-net12 A2 XU42-net9 VDD p w=1.37u l=0.18u
MU42-M_u3 net12 A3 XU42-net12 VDD p w=1.37u l=0.18u
M_u4_0-M_u3 Z net12 VDD VDD p w=1.37u l=0.18u
M_u4_1-M_u3 Z net12 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OR3D4BWP7T A1 A2 A3 Z VDD VSS 
MI1-M_u6 p0 A3 VSS VSS n w=0.5u l=0.18u
MI1-M_u5 p0 A2 VSS VSS n w=0.5u l=0.18u
MI1-M_u4 p0 A1 VSS VSS n w=0.5u l=0.18u
MU42-M_u6 p0 A3 VSS VSS n w=0.5u l=0.18u
MU42-M_u5 p0 A2 VSS VSS n w=0.5u l=0.18u
MU42-M_u4 p0 A1 VSS VSS n w=0.5u l=0.18u
M_u4_0-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u4_1-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u4_2-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u4_3-M_u2 Z p0 VSS VSS n w=1u l=0.18u
MI1-M_u1 XI1-net9 A1 VDD VDD p w=1.37u l=0.18u
MI1-M_u2 XI1-net12 A2 XI1-net9 VDD p w=1.37u l=0.18u
MI1-M_u3 p0 A3 XI1-net12 VDD p w=1.37u l=0.18u
MU42-M_u1 XU42-net9 A1 VDD VDD p w=1.37u l=0.18u
MU42-M_u2 XU42-net12 A2 XU42-net9 VDD p w=1.37u l=0.18u
MU42-M_u3 p0 A3 XU42-net12 VDD p w=1.37u l=0.18u
M_u4_0-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u4_1-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u4_2-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u4_3-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OR3XD1BWP7T A1 A2 A3 Z VDD VSS 
MU42-M_u6 net7 A3 VSS VSS n w=1u l=0.18u
MU42-M_u5 net7 A2 VSS VSS n w=1u l=0.18u
MU42-M_u4 net7 A1 VSS VSS n w=1u l=0.18u
M_u4-M_u2 Z net7 VSS VSS n w=1u l=0.18u
MU42-M_u1 XU42-net9 A1 VDD VDD p w=1.37u l=0.18u
MU42-M_u2 XU42-net12 A2 XU42-net9 VDD p w=1.37u l=0.18u
MU42-M_u3 net7 A3 XU42-net12 VDD p w=1.37u l=0.18u
M_u4-M_u3 Z net7 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OR4D0BWP7T A1 A2 A3 A4 Z VDD VSS 
MU8-M_u4 net14 A1 VSS VSS n w=0.5u l=0.18u
MU8-M_u3 net14 A2 VSS VSS n w=0.5u l=0.18u
MU8-M_u5 net14 A3 VSS VSS n w=0.5u l=0.18u
MU8-M_u8 net14 A4 VSS VSS n w=0.5u l=0.18u
M_u3-M_u2 Z net14 VSS VSS n w=0.5u l=0.18u
MU8-M_u7 net14 A4 XU8-net7 VDD p w=0.685u l=0.18u
MU8-M_u6 XU8-net7 A3 XU8-net10 VDD p w=0.685u l=0.18u
MU8-M_u2 XU8-net10 A2 XU8-net13 VDD p w=0.685u l=0.18u
MU8-M_u1 XU8-net13 A1 VDD VDD p w=0.685u l=0.18u
M_u3-M_u3 Z net14 VDD VDD p w=0.685u l=0.18u
.ends
.subckt OR4D1BWP7T A1 A2 A3 A4 Z VDD VSS 
MU8-M_u4 net14 A1 VSS VSS n w=0.5u l=0.18u
MU8-M_u3 net14 A2 VSS VSS n w=0.5u l=0.18u
MU8-M_u5 net14 A3 VSS VSS n w=0.5u l=0.18u
MU8-M_u8 net14 A4 VSS VSS n w=0.5u l=0.18u
M_u3-M_u2 Z net14 VSS VSS n w=1u l=0.18u
MU8-M_u7 net14 A4 XU8-net7 VDD p w=1.37u l=0.18u
MU8-M_u6 XU8-net7 A3 XU8-net10 VDD p w=1.37u l=0.18u
MU8-M_u2 XU8-net10 A2 XU8-net13 VDD p w=1.37u l=0.18u
MU8-M_u1 XU8-net13 A1 VDD VDD p w=1.37u l=0.18u
M_u3-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OR4D2BWP7T A1 A2 A3 A4 Z VDD VSS 
MU8-M_u4 net14 A1 VSS VSS n w=0.5u l=0.18u
MU8-M_u3 net14 A2 VSS VSS n w=0.5u l=0.18u
MU8-M_u5 net14 A3 VSS VSS n w=0.5u l=0.18u
MU8-M_u8 net14 A4 VSS VSS n w=0.5u l=0.18u
M_u3_0-M_u2 Z net14 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z net14 VSS VSS n w=1u l=0.18u
MU8-M_u7 net14 A4 XU8-net7 VDD p w=1.37u l=0.18u
MU8-M_u6 XU8-net7 A3 XU8-net10 VDD p w=1.37u l=0.18u
MU8-M_u2 XU8-net10 A2 XU8-net13 VDD p w=1.37u l=0.18u
MU8-M_u1 XU8-net13 A1 VDD VDD p w=1.37u l=0.18u
M_u3_0-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OR4D4BWP7T A1 A2 A3 A4 Z VDD VSS 
MU8_0-M_u4 p0 A1 VSS VSS n w=0.5u l=0.18u
MU8_0-M_u3 p0 A2 VSS VSS n w=0.5u l=0.18u
MU8_0-M_u5 p0 A3 VSS VSS n w=0.5u l=0.18u
MU8_0-M_u8 p0 A4 VSS VSS n w=0.5u l=0.18u
MU8_1-M_u4 p0 A1 VSS VSS n w=0.5u l=0.18u
MU8_1-M_u3 p0 A2 VSS VSS n w=0.5u l=0.18u
MU8_1-M_u5 p0 A3 VSS VSS n w=0.5u l=0.18u
MU8_1-M_u8 p0 A4 VSS VSS n w=0.5u l=0.18u
M_u3_0-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_1-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_2-M_u2 Z p0 VSS VSS n w=1u l=0.18u
M_u3_3-M_u2 Z p0 VSS VSS n w=1u l=0.18u
MU8_0-M_u7 p0 A4 XU8_0-net7 VDD p w=1.37u l=0.18u
MU8_0-M_u6 XU8_0-net7 A3 XU8_0-net10 VDD p w=1.37u l=0.18u
MU8_0-M_u2 XU8_0-net10 A2 XU8_0-net13 VDD p w=1.37u l=0.18u
MU8_0-M_u1 XU8_0-net13 A1 VDD VDD p w=1.37u l=0.18u
MU8_1-M_u7 p0 A4 XU8_1-net7 VDD p w=1.37u l=0.18u
MU8_1-M_u6 XU8_1-net7 A3 XU8_1-net10 VDD p w=1.37u l=0.18u
MU8_1-M_u2 XU8_1-net10 A2 XU8_1-net13 VDD p w=1.37u l=0.18u
MU8_1-M_u1 XU8_1-net13 A1 VDD VDD p w=1.37u l=0.18u
M_u3_0-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_1-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_2-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
M_u3_3-M_u3 Z p0 VDD VDD p w=1.37u l=0.18u
.ends
.subckt OR4XD1BWP7T A1 A2 A3 A4 Z VDD VSS 
MU8-M_u4 net14 A1 VSS VSS n w=1u l=0.18u
MU8-M_u3 net14 A2 VSS VSS n w=1u l=0.18u
MU8-M_u5 net14 A3 VSS VSS n w=1u l=0.18u
MU8-M_u8 net14 A4 VSS VSS n w=1u l=0.18u
M_u3-M_u2 Z net14 VSS VSS n w=1u l=0.18u
MU8-M_u7 net14 A4 XU8-net7 VDD p w=1.37u l=0.18u
MU8-M_u6 XU8-net7 A3 XU8-net10 VDD p w=1.37u l=0.18u
MU8-M_u2 XU8-net10 A2 XU8-net13 VDD p w=1.37u l=0.18u
MU8-M_u1 XU8-net13 A1 VDD VDD p w=1.37u l=0.18u
M_u3-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
.ends
.subckt SDFCND0BWP7T SI D SE CP CDN Q QN VDD VSS 
MI150 net62 INCPB net163 VSS n w=0.42u l=0.18u
MI149 d1 INCP net163 VSS n w=0.91u l=0.18u
MI165 net63 d1 VSS VSS n w=0.42u l=0.18u
MI164 net82 CDN net63 VSS n w=0.42u l=0.18u
MI47 d0 INCP net82 VSS n w=0.42u l=0.18u
MI169 net177 net120 net69 VSS n w=1u l=0.18u
MI77 d0 INCPB net177 VSS n w=0.8u l=0.18u
MI161 net67 SI VSS VSS n w=0.42u l=0.18u
MI160 net177 SE net67 VSS n w=0.42u l=0.18u
MI158-M_u4 XI158-net6 CDN VSS VSS n w=0.97u l=0.18u
MI158-M_u3 d3 net163 XI158-net6 VSS n w=0.97u l=0.18u
MI166-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI151-M_u2 QN net62 VSS VSS n w=0.5u l=0.18u
MI152-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI153-M_u2 net62 d3 VSS VSS n w=0.42u l=0.18u
MI85-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI173-M_u2 net69 D VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI158-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI158-M_u1 d3 net163 VDD VDD p w=1.31u l=0.18u
MI166-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI151-M_u3 QN net62 VDD VDD p w=0.685u l=0.18u
MI152-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI153-M_u3 net62 d3 VDD VDD p w=0.685u l=0.18u
MI85-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI173-M_u3 net69 D VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI155 net62 INCP net163 VDD p w=0.42u l=0.18u
MI170 net177 SE net69 VDD p w=1.095u l=0.18u
MI163 d0 INCPB net166 VDD p w=0.42u l=0.18u
MI162 net166 CDN VDD VDD p w=0.42u l=0.18u
MI71 net177 net120 net142 VDD p w=0.42u l=0.18u
MI74 d0 INCP net177 VDD p w=0.92u l=0.18u
MI75 net142 SI VDD VDD p w=0.42u l=0.18u
MI44 net166 d1 VDD VDD p w=0.42u l=0.18u
MI154 d1 INCPB net163 VDD p w=0.62u l=0.18u
.ends
.subckt SDFCND1BWP7T SI D SE CP CDN Q QN VDD VSS 
MI150 net62 INCPB net163 VSS n w=0.42u l=0.18u
MI149 d1 INCP net163 VSS n w=0.91u l=0.18u
MI165 net63 d1 VSS VSS n w=0.42u l=0.18u
MI164 net82 CDN net63 VSS n w=0.42u l=0.18u
MI47 d0 INCP net82 VSS n w=0.42u l=0.18u
MI169 net177 net120 net69 VSS n w=1u l=0.18u
MI77 d0 INCPB net177 VSS n w=0.8u l=0.18u
MI161 net67 SI VSS VSS n w=0.42u l=0.18u
MI160 net177 SE net67 VSS n w=0.42u l=0.18u
MI158-M_u4 XI158-net6 CDN VSS VSS n w=0.97u l=0.18u
MI158-M_u3 d3 net163 XI158-net6 VSS n w=1u l=0.18u
MI166-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI151-M_u2 QN net62 VSS VSS n w=0.94u l=0.18u
MI152-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI153-M_u2 net62 d3 VSS VSS n w=0.42u l=0.18u
MI85-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI173-M_u2 net69 D VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI158-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI158-M_u1 d3 net163 VDD VDD p w=1.37u l=0.18u
MI166-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI151-M_u3 QN net62 VDD VDD p w=1.37u l=0.18u
MI152-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI153-M_u3 net62 d3 VDD VDD p w=0.685u l=0.18u
MI85-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI173-M_u3 net69 D VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI155 net62 INCP net163 VDD p w=0.42u l=0.18u
MI170 net177 SE net69 VDD p w=1.095u l=0.18u
MI163 d0 INCPB net166 VDD p w=0.42u l=0.18u
MI162 net166 CDN VDD VDD p w=0.42u l=0.18u
MI71 net177 net120 net142 VDD p w=0.42u l=0.18u
MI74 d0 INCP net177 VDD p w=0.92u l=0.18u
MI75 net142 SI VDD VDD p w=0.42u l=0.18u
MI44 net166 d1 VDD VDD p w=0.42u l=0.18u
MI154 d1 INCPB net163 VDD p w=0.62u l=0.18u
.ends
.subckt SDFCND2BWP7T SI D SE CP CDN Q QN VDD VSS 
MI150 net62 INCPB net163 VSS n w=0.42u l=0.18u
MI149 d1 INCP net163 VSS n w=0.91u l=0.18u
MI165 net63 d1 VSS VSS n w=0.42u l=0.18u
MI164 net82 CDN net63 VSS n w=0.42u l=0.18u
MI47 d0 INCP net82 VSS n w=0.42u l=0.18u
MI169 net177 net120 net69 VSS n w=1u l=0.18u
MI77 d0 INCPB net177 VSS n w=0.8u l=0.18u
MI161 net67 SI VSS VSS n w=0.42u l=0.18u
MI160 net177 SE net67 VSS n w=0.42u l=0.18u
MI158-M_u4 XI158-net6 CDN VSS VSS n w=0.97u l=0.18u
MI158-M_u3 d3 net163 XI158-net6 VSS n w=0.97u l=0.18u
MI166-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI151_0-M_u2 QN net62 VSS VSS n w=1u l=0.18u
MI151_1-M_u2 QN net62 VSS VSS n w=1u l=0.18u
MI152_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI152_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI153-M_u2 net62 d3 VSS VSS n w=0.97u l=0.18u
MI85-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI173-M_u2 net69 D VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI158-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI158-M_u1 d3 net163 VDD VDD p w=1.23u l=0.18u
MI166-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI151_0-M_u3 QN net62 VDD VDD p w=1.3u l=0.18u
MI151_1-M_u3 QN net62 VDD VDD p w=1.3u l=0.18u
MI152_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI152_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI153-M_u3 net62 d3 VDD VDD p w=0.97u l=0.18u
MI85-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI173-M_u3 net69 D VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI155 net62 INCP net163 VDD p w=0.42u l=0.18u
MI170 net177 SE net69 VDD p w=1.095u l=0.18u
MI163 d0 INCPB net166 VDD p w=0.42u l=0.18u
MI162 net166 CDN VDD VDD p w=0.42u l=0.18u
MI71 net177 net120 net142 VDD p w=0.42u l=0.18u
MI74 d0 INCP net177 VDD p w=0.92u l=0.18u
MI75 net142 SI VDD VDD p w=0.42u l=0.18u
MI44 net166 d1 VDD VDD p w=0.42u l=0.18u
MI154 d1 INCPB net163 VDD p w=0.62u l=0.18u
.ends
.subckt SDFCNQD0BWP7T SI D SE CP CDN Q VDD VSS 
MI150 net62 INCPB net163 VSS n w=0.42u l=0.18u
MI149 d1 INCP net163 VSS n w=0.91u l=0.18u
MI165 net63 d1 VSS VSS n w=0.42u l=0.18u
MI164 net82 CDN net63 VSS n w=0.42u l=0.18u
MI47 d0 INCP net82 VSS n w=0.42u l=0.18u
MI169 net177 net120 net69 VSS n w=1u l=0.18u
MI77 d0 INCPB net177 VSS n w=0.91u l=0.18u
MI161 net67 SI VSS VSS n w=0.42u l=0.18u
MI160 net177 SE net67 VSS n w=0.42u l=0.18u
MI158-M_u4 XI158-net6 CDN VSS VSS n w=0.97u l=0.18u
MI158-M_u3 d3 net163 XI158-net6 VSS n w=0.97u l=0.18u
MI166-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI152-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI153-M_u2 net62 d3 VSS VSS n w=0.42u l=0.18u
MI85-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI173-M_u2 net69 D VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI158-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI158-M_u1 d3 net163 VDD VDD p w=1.37u l=0.18u
MI166-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI152-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI153-M_u3 net62 d3 VDD VDD p w=0.42u l=0.18u
MI85-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI173-M_u3 net69 D VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI155 net62 INCP net163 VDD p w=0.42u l=0.18u
MI170 net177 SE net69 VDD p w=1.095u l=0.18u
MI163 d0 INCPB net166 VDD p w=0.42u l=0.18u
MI162 net166 CDN VDD VDD p w=0.42u l=0.18u
MI71 net177 net120 net142 VDD p w=0.42u l=0.18u
MI74 d0 INCP net177 VDD p w=0.92u l=0.18u
MI75 net142 SI VDD VDD p w=0.42u l=0.18u
MI44 net166 d1 VDD VDD p w=0.42u l=0.18u
MI154 d1 INCPB net163 VDD p w=0.62u l=0.18u
.ends
.subckt SDFCNQD1BWP7T SI D SE CP CDN Q VDD VSS 
MI150 net62 INCPB net163 VSS n w=0.42u l=0.18u
MI149 d1 INCP net163 VSS n w=0.91u l=0.18u
MI165 net63 d1 VSS VSS n w=0.42u l=0.18u
MI164 net82 CDN net63 VSS n w=0.42u l=0.18u
MI47 d0 INCP net82 VSS n w=0.42u l=0.18u
MI169 net177 net120 net69 VSS n w=1u l=0.18u
MI77 d0 INCPB net177 VSS n w=0.91u l=0.18u
MI161 net67 SI VSS VSS n w=0.42u l=0.18u
MI160 net177 SE net67 VSS n w=0.42u l=0.18u
MI158-M_u4 XI158-net6 CDN VSS VSS n w=0.97u l=0.18u
MI158-M_u3 d3 net163 XI158-net6 VSS n w=0.97u l=0.18u
MI166-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI152-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI153-M_u2 net62 d3 VSS VSS n w=0.42u l=0.18u
MI85-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI173-M_u2 net69 D VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI158-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI158-M_u1 d3 net163 VDD VDD p w=1.37u l=0.18u
MI166-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI152-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI153-M_u3 net62 d3 VDD VDD p w=0.42u l=0.18u
MI85-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI173-M_u3 net69 D VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI155 net62 INCP net163 VDD p w=0.42u l=0.18u
MI170 net177 SE net69 VDD p w=1.095u l=0.18u
MI163 d0 INCPB net166 VDD p w=0.42u l=0.18u
MI162 net166 CDN VDD VDD p w=0.42u l=0.18u
MI71 net177 net120 net142 VDD p w=0.42u l=0.18u
MI74 d0 INCP net177 VDD p w=0.92u l=0.18u
MI75 net142 SI VDD VDD p w=0.42u l=0.18u
MI44 net166 d1 VDD VDD p w=0.42u l=0.18u
MI154 d1 INCPB net163 VDD p w=0.62u l=0.18u
.ends
.subckt SDFCNQD2BWP7T SI D SE CP CDN Q VDD VSS 
MI150 net62 INCPB net163 VSS n w=0.42u l=0.18u
MI149 d1 INCP net163 VSS n w=0.91u l=0.18u
MI165 net63 d1 VSS VSS n w=0.42u l=0.18u
MI164 net82 CDN net63 VSS n w=0.42u l=0.18u
MI47 d0 INCP net82 VSS n w=0.42u l=0.18u
MI169 net177 net120 net69 VSS n w=1u l=0.18u
MI77 d0 INCPB net177 VSS n w=0.91u l=0.18u
MI161 net67 SI VSS VSS n w=0.42u l=0.18u
MI160 net177 SE net67 VSS n w=0.42u l=0.18u
MI158-M_u4 XI158-net6 CDN VSS VSS n w=0.97u l=0.18u
MI158-M_u3 d3 net163 XI158-net6 VSS n w=0.97u l=0.18u
MI166-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI152_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI152_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI153-M_u2 net62 d3 VSS VSS n w=0.42u l=0.18u
MI85-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI173-M_u2 net69 D VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI158-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI158-M_u1 d3 net163 VDD VDD p w=1.37u l=0.18u
MI166-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI152_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI152_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI153-M_u3 net62 d3 VDD VDD p w=0.42u l=0.18u
MI85-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI173-M_u3 net69 D VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI155 net62 INCP net163 VDD p w=0.42u l=0.18u
MI170 net177 SE net69 VDD p w=1.095u l=0.18u
MI163 d0 INCPB net166 VDD p w=0.42u l=0.18u
MI162 net166 CDN VDD VDD p w=0.42u l=0.18u
MI71 net177 net120 net142 VDD p w=0.42u l=0.18u
MI74 d0 INCP net177 VDD p w=0.92u l=0.18u
MI75 net142 SI VDD VDD p w=0.42u l=0.18u
MI44 net166 d1 VDD VDD p w=0.42u l=0.18u
MI154 d1 INCPB net163 VDD p w=0.62u l=0.18u
.ends
.subckt SDFD0BWP7T SI D SE CP Q QN VDD VSS 
MI39 net13 net57 net64 VSS n w=1u l=0.18u
MI25 net65 INCP d2 VSS n w=0.91u l=0.18u
MI13 net28 INCP net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net55 INCPB d2 VSS n w=0.42u l=0.18u
MU65 net28 INCPB net13 VSS n w=0.5u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net64 D VSS VSS n w=1u l=0.18u
MI28-M_u2 net55 d3 VSS VSS n w=0.42u l=0.18u
MI30-M_u2 d3 d2 VSS VSS n w=0.5u l=0.18u
MI33-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI34-M_u2 QN net55 VSS VSS n w=0.5u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MU84-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net55 d3 VDD VDD p w=0.685u l=0.18u
MI30-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI33-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI34-M_u3 QN net55 VDD VDD p w=0.685u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MU84-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net55 INCP d2 VDD p w=0.42u l=0.18u
MI36 net65 INCPB d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net0126 D VDD VDD p w=1.18u l=0.18u
MU62 net28 INCP net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 INCPB net137 VDD p w=0.42u l=0.18u
MI40 net13 SE net0126 VDD p w=1.18u l=0.18u
.ends
.subckt SDFD1BWP7T SI D SE CP Q QN VDD VSS 
MI39 net13 net57 net64 VSS n w=1u l=0.18u
MI25 net65 INCP d2 VSS n w=0.91u l=0.18u
MI13 net28 INCP net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net55 INCPB d2 VSS n w=0.42u l=0.18u
MU65 net28 INCPB net13 VSS n w=0.5u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net64 D VSS VSS n w=1u l=0.18u
MI28-M_u2 net55 d3 VSS VSS n w=0.42u l=0.18u
MI30-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI33-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI34-M_u2 QN net55 VSS VSS n w=0.94u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MU84-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net55 d3 VDD VDD p w=0.685u l=0.18u
MI30-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI33-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI34-M_u3 QN net55 VDD VDD p w=1.37u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MU84-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net55 INCP d2 VDD p w=0.42u l=0.18u
MI36 net65 INCPB d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net0126 D VDD VDD p w=1.18u l=0.18u
MU62 net28 INCP net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 INCPB net137 VDD p w=0.42u l=0.18u
MI40 net13 SE net0126 VDD p w=1.18u l=0.18u
.ends
.subckt SDFD2BWP7T SI D SE CP Q QN VDD VSS 
MI39 net13 net57 net64 VSS n w=1u l=0.18u
MI25 net65 INCP d2 VSS n w=0.91u l=0.18u
MI13 net28 INCP net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net068 INCPB d2 VSS n w=0.42u l=0.18u
MU65 net28 INCPB net13 VSS n w=0.5u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net64 D VSS VSS n w=1u l=0.18u
MI28-M_u2 net068 d3 VSS VSS n w=1u l=0.18u
MI30_0-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI30_1-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI33_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI33_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI34_0-M_u2 QN net068 VSS VSS n w=1u l=0.18u
MI34_1-M_u2 QN net068 VSS VSS n w=1u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MU84-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net068 d3 VDD VDD p w=1.37u l=0.18u
MI30_0-M_u3 d3 d2 VDD VDD p w=1.23u l=0.18u
MI30_1-M_u3 d3 d2 VDD VDD p w=1.23u l=0.18u
MI33_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI33_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI34_0-M_u3 QN net068 VDD VDD p w=1.3u l=0.18u
MI34_1-M_u3 QN net068 VDD VDD p w=1.3u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MU84-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net068 INCP d2 VDD p w=0.42u l=0.18u
MI36 net65 INCPB d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net0126 D VDD VDD p w=1.18u l=0.18u
MU62 net28 INCP net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 INCPB net137 VDD p w=0.42u l=0.18u
MI40 net13 SE net0126 VDD p w=1.18u l=0.18u
.ends
.subckt SDFKCND0BWP7T SI D SE CP CN Q QN VDD VSS 
MI138-M_u2 QN net69 VSS VSS n w=0.5u l=0.18u
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI136-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net69 net105 VSS VSS n w=0.5u l=0.18u
MI116-M_u2 Q net105 VSS VSS n w=0.5u l=0.18u
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net69 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI79 net132 D net135 VSS n w=1u l=0.18u
MI80 net135 CN VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI138-M_u3 QN net69 VDD VDD p w=0.685u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI136-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net69 net105 VDD VDD p w=0.685u l=0.18u
MI116-M_u3 Q net105 VDD VDD p w=0.685u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net69 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI74 VDD CN net132 VDD p w=0.42u l=0.18u
MI77 VDD D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKCND1BWP7T SI D SE CP CN Q QN VDD VSS 
MI138-M_u2 QN net69 VSS VSS n w=1u l=0.18u
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI136-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net69 net105 VSS VSS n w=0.5u l=0.18u
MI116-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net69 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI79 net132 D net135 VSS n w=1u l=0.18u
MI80 net135 CN VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI138-M_u3 QN net69 VDD VDD p w=1.37u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI136-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net69 net105 VDD VDD p w=0.685u l=0.18u
MI116-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net69 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI74 VDD CN net132 VDD p w=0.42u l=0.18u
MI77 VDD D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKCND2BWP7T SI D SE CP CN Q QN VDD VSS 
MI138_0-M_u2 QN net089 VSS VSS n w=1u l=0.18u
MI138_1-M_u2 QN net089 VSS VSS n w=1u l=0.18u
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI136-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net089 net105 VSS VSS n w=0.97u l=0.18u
MI116_0-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI116_1-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net089 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI79 net132 D net135 VSS n w=1u l=0.18u
MI80 net135 CN VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI138_0-M_u3 QN net089 VDD VDD p w=1.37u l=0.18u
MI138_1-M_u3 QN net089 VDD VDD p w=1.37u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI136-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net089 net105 VDD VDD p w=1.37u l=0.18u
MI116_0-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI116_1-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net089 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI74 VDD CN net132 VDD p w=0.42u l=0.18u
MI77 VDD D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKCNQD0BWP7T SI D SE CP CN Q VDD VSS 
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI136-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net69 net105 VSS VSS n w=0.5u l=0.18u
MI116-M_u2 Q net105 VSS VSS n w=0.5u l=0.18u
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net69 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI79 net132 D net135 VSS n w=1u l=0.18u
MI80 net135 CN VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI136-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net69 net105 VDD VDD p w=0.685u l=0.18u
MI116-M_u3 Q net105 VDD VDD p w=0.685u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net69 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI74 VDD CN net132 VDD p w=0.42u l=0.18u
MI77 VDD D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKCNQD1BWP7T SI D SE CP CN Q VDD VSS 
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI136-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net69 net105 VSS VSS n w=0.5u l=0.18u
MI116-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net69 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI79 net132 D net135 VSS n w=1u l=0.18u
MI80 net135 CN VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI136-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net69 net105 VDD VDD p w=0.685u l=0.18u
MI116-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net69 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI74 VDD CN net132 VDD p w=0.42u l=0.18u
MI77 VDD D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKCNQD2BWP7T SI D SE CP CN Q VDD VSS 
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI136-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net69 net105 VSS VSS n w=0.5u l=0.18u
MI116_0-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI116_1-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net69 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI79 net132 D net135 VSS n w=1u l=0.18u
MI80 net135 CN VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI136-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net69 net105 VDD VDD p w=0.685u l=0.18u
MI116_0-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI116_1-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net69 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI74 VDD CN net132 VDD p w=0.42u l=0.18u
MI77 VDD D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKSND0BWP7T SI D SE CP SN Q QN VDD VSS 
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net69 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI78 net132 net116 VSS VSS n w=0.42u l=0.18u
MI79 net132 D VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI138-M_u2 QN net69 VSS VSS n w=0.5u l=0.18u
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI139-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net69 net105 VSS VSS n w=0.5u l=0.18u
MI116-M_u2 Q net105 VSS VSS n w=0.5u l=0.18u
MI72-M_u2 net116 SN VSS VSS n w=0.5u l=0.18u
MI138-M_u3 QN net69 VDD VDD p w=0.685u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI139-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net69 net105 VDD VDD p w=0.685u l=0.18u
MI116-M_u3 Q net105 VDD VDD p w=0.685u l=0.18u
MI72-M_u3 net116 SN VDD VDD p w=0.685u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net69 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI75 VDD net116 net139 VDD p w=1.37u l=0.18u
MI77 net139 D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKSND1BWP7T SI D SE CP SN Q QN VDD VSS 
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net69 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI78 net132 net116 VSS VSS n w=0.42u l=0.18u
MI79 net132 D VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI138-M_u2 QN net69 VSS VSS n w=1u l=0.18u
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI139-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net69 net105 VSS VSS n w=0.5u l=0.18u
MI116-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI72-M_u2 net116 SN VSS VSS n w=0.5u l=0.18u
MI138-M_u3 QN net69 VDD VDD p w=1.37u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI139-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net69 net105 VDD VDD p w=0.685u l=0.18u
MI116-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI72-M_u3 net116 SN VDD VDD p w=0.685u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net69 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI75 VDD net116 net139 VDD p w=1.37u l=0.18u
MI77 net139 D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKSND2BWP7T SI D SE CP SN Q QN VDD VSS 
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net0120 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI78 net132 net116 VSS VSS n w=0.42u l=0.18u
MI79 net132 D VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI138_0-M_u2 QN net0120 VSS VSS n w=1u l=0.18u
MI138_1-M_u2 QN net0120 VSS VSS n w=1u l=0.18u
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI139-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net0120 net105 VSS VSS n w=0.97u l=0.18u
MI116_0-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI116_1-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI72-M_u2 net116 SN VSS VSS n w=0.5u l=0.18u
MI138_0-M_u3 QN net0120 VDD VDD p w=1.37u l=0.18u
MI138_1-M_u3 QN net0120 VDD VDD p w=1.37u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI139-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net0120 net105 VDD VDD p w=1.37u l=0.18u
MI116_0-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI116_1-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI72-M_u3 net116 SN VDD VDD p w=0.685u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net0120 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI75 VDD net116 net139 VDD p w=1.37u l=0.18u
MI77 net139 D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKSNQD0BWP7T SI D SE CP SN Q VDD VSS 
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net69 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI78 net132 net116 VSS VSS n w=0.42u l=0.18u
MI79 net132 D VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI139-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net69 net105 VSS VSS n w=0.5u l=0.18u
MI116-M_u2 Q net105 VSS VSS n w=0.5u l=0.18u
MI72-M_u2 net116 SN VSS VSS n w=0.5u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI139-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net69 net105 VDD VDD p w=0.685u l=0.18u
MI116-M_u3 Q net105 VDD VDD p w=0.685u l=0.18u
MI72-M_u3 net116 SN VDD VDD p w=0.685u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net69 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI75 VDD net116 net139 VDD p w=1.37u l=0.18u
MI77 net139 D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKSNQD1BWP7T SI D SE CP SN Q VDD VSS 
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net69 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI78 net132 net116 VSS VSS n w=0.42u l=0.18u
MI79 net132 D VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI139-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net69 net105 VSS VSS n w=0.5u l=0.18u
MI116-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI72-M_u2 net116 SN VSS VSS n w=0.5u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI139-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net69 net105 VDD VDD p w=0.685u l=0.18u
MI116-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI72-M_u3 net116 SN VDD VDD p w=0.685u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net69 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI75 VDD net116 net139 VDD p w=1.37u l=0.18u
MI77 net139 D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFKSNQD2BWP7T SI D SE CP SN Q VDD VSS 
MI112 net93 INCP net105 VSS n w=0.91u l=0.18u
MI135 net87 SI VSS VSS n w=0.42u l=0.18u
MI128 net132 net107 net90 VSS n w=1u l=0.18u
MI29 net105 INCPB net79 VSS n w=0.42u l=0.18u
MI26 net79 net69 VSS VSS n w=0.42u l=0.18u
MI126 net109 INCPB net155 VSS n w=0.91u l=0.18u
MI101 net155 INCP net95 VSS n w=0.42u l=0.18u
MI102 net95 net93 VSS VSS n w=0.42u l=0.18u
MI78 net132 net116 VSS VSS n w=0.42u l=0.18u
MI79 net132 D VSS VSS n w=1u l=0.18u
MI134 net90 SE net87 VSS n w=0.42u l=0.18u
MI48-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI130-M_u2 net109 net90 VSS VSS n w=1u l=0.18u
MI49-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI139-M_u2 net107 SE VSS VSS n w=0.5u l=0.18u
MI42-M_u2 net93 net155 VSS VSS n w=0.54u l=0.18u
MI115-M_u2 net69 net105 VSS VSS n w=0.5u l=0.18u
MI116_0-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI116_1-M_u2 Q net105 VSS VSS n w=1u l=0.18u
MI72-M_u2 net116 SN VSS VSS n w=0.5u l=0.18u
MI48-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI130-M_u3 net109 net90 VDD VDD p w=1.23u l=0.18u
MI49-M_u3 INCP INCPB VDD VDD p w=0.63u l=0.18u
MI139-M_u3 net107 SE VDD VDD p w=0.685u l=0.18u
MI42-M_u3 net93 net155 VDD VDD p w=0.96u l=0.18u
MI115-M_u3 net69 net105 VDD VDD p w=0.685u l=0.18u
MI116_0-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI116_1-M_u3 Q net105 VDD VDD p w=1.37u l=0.18u
MI72-M_u3 net116 SN VDD VDD p w=0.685u l=0.18u
MI28 net105 INCP net168 VDD p w=0.42u l=0.18u
MI129 net132 SE net90 VDD p w=1.15u l=0.18u
MI24 net168 net69 VDD VDD p w=0.42u l=0.18u
MI133 net138 net107 net90 VDD p w=0.42u l=0.18u
MI119 net93 INCPB net105 VDD p w=1.34u l=0.18u
MI127 net109 INCP net155 VDD p w=0.92u l=0.18u
MI99 net155 INCPB net153 VDD p w=0.42u l=0.18u
MI100 net153 net93 VDD VDD p w=0.42u l=0.18u
MI131 VDD SI net138 VDD p w=0.42u l=0.18u
MI75 VDD net116 net139 VDD p w=1.37u l=0.18u
MI77 net139 D net132 VDD p w=1.37u l=0.18u
.ends
.subckt SDFNCND0BWP7T SI D SE CPN CDN Q QN VDD VSS 
MI162 net177 net120 net065 VSS n w=1u l=0.18u
MI150 net62 net101 d2 VSS n w=0.42u l=0.18u
MI149 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI49 net79 d1 VSS VSS n w=0.42u l=0.18u
MI48 net82 CDN net79 VSS n w=0.42u l=0.18u
MI47 d0 INCPB net82 VSS n w=0.42u l=0.18u
MI77 d0 net101 net177 VSS n w=0.97u l=0.18u
MI78 net89 SI VSS VSS n w=0.42u l=0.18u
MI80 net177 SE net89 VSS n w=0.42u l=0.18u
MI81 net065 D VSS VSS n w=1u l=0.18u
MI158-M_u4 XI158-net6 CDN VSS VSS n w=0.97u l=0.18u
MI158-M_u3 d3 d2 XI158-net6 VSS n w=0.97u l=0.18u
MI151-M_u2 QN net62 VSS VSS n w=0.5u l=0.18u
MI152-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI153-M_u2 net62 d3 VSS VSS n w=0.42u l=0.18u
MI85-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI165-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI32-M_u2 net101 INCPB VSS VSS n w=0.5u l=0.18u
MI158-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI158-M_u1 d3 d2 VDD VDD p w=1.31u l=0.18u
MI151-M_u3 QN net62 VDD VDD p w=0.685u l=0.18u
MI152-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI153-M_u3 net62 d3 VDD VDD p w=0.685u l=0.18u
MI85-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI165-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI32-M_u3 net101 INCPB VDD VDD p w=0.685u l=0.18u
MI164 net177 SE net069 VDD p w=1.095u l=0.18u
MI155 net62 INCPB d2 VDD p w=0.42u l=0.18u
MI45 d0 net101 net166 VDD p w=0.42u l=0.18u
MI43 net166 d1 VDD VDD p w=0.42u l=0.18u
MI163 net177 net120 net142 VDD p w=0.42u l=0.18u
MI73 net069 D VDD VDD p w=1.37u l=0.18u
MI74 d0 INCPB net177 VDD p w=0.92u l=0.18u
MI75 net142 SI VDD VDD p w=0.42u l=0.18u
MI44 net166 CDN VDD VDD p w=0.42u l=0.18u
MI154 d1 net101 d2 VDD p w=0.62u l=0.18u
.ends
.subckt SDFNCND1BWP7T SI D SE CPN CDN Q QN VDD VSS 
MI162 net177 net120 net065 VSS n w=1u l=0.18u
MI150 net62 net101 d2 VSS n w=0.42u l=0.18u
MI149 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI49 net79 d1 VSS VSS n w=0.42u l=0.18u
MI48 net82 CDN net79 VSS n w=0.42u l=0.18u
MI47 d0 INCPB net82 VSS n w=0.42u l=0.18u
MI77 d0 net101 net177 VSS n w=0.97u l=0.18u
MI78 net89 SI VSS VSS n w=0.42u l=0.18u
MI80 net177 SE net89 VSS n w=0.42u l=0.18u
MI81 net065 D VSS VSS n w=1u l=0.18u
MI158-M_u4 XI158-net6 CDN VSS VSS n w=0.97u l=0.18u
MI158-M_u3 d3 d2 XI158-net6 VSS n w=1u l=0.18u
MI151-M_u2 QN net62 VSS VSS n w=0.94u l=0.18u
MI152-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI153-M_u2 net62 d3 VSS VSS n w=0.42u l=0.18u
MI85-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI165-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI32-M_u2 net101 INCPB VSS VSS n w=0.5u l=0.18u
MI158-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI158-M_u1 d3 d2 VDD VDD p w=1.37u l=0.18u
MI151-M_u3 QN net62 VDD VDD p w=1.37u l=0.18u
MI152-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI153-M_u3 net62 d3 VDD VDD p w=0.685u l=0.18u
MI85-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI165-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI32-M_u3 net101 INCPB VDD VDD p w=0.685u l=0.18u
MI164 net177 SE net069 VDD p w=1.095u l=0.18u
MI155 net62 INCPB d2 VDD p w=0.42u l=0.18u
MI45 d0 net101 net166 VDD p w=0.42u l=0.18u
MI43 net166 d1 VDD VDD p w=0.42u l=0.18u
MI163 net177 net120 net142 VDD p w=0.42u l=0.18u
MI73 net069 D VDD VDD p w=1.37u l=0.18u
MI74 d0 INCPB net177 VDD p w=0.92u l=0.18u
MI75 net142 SI VDD VDD p w=0.42u l=0.18u
MI44 net166 CDN VDD VDD p w=0.42u l=0.18u
MI154 d1 net101 d2 VDD p w=0.62u l=0.18u
.ends
.subckt SDFNCND2BWP7T SI D SE CPN CDN Q QN VDD VSS 
MI162 net177 net120 net066 VSS n w=1u l=0.18u
MI150 net62 net101 d2 VSS n w=0.42u l=0.18u
MI149 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI49 net79 d1 VSS VSS n w=0.42u l=0.18u
MI48 net82 CDN net79 VSS n w=0.42u l=0.18u
MI47 d0 INCPB net82 VSS n w=0.42u l=0.18u
MI77 d0 net101 net177 VSS n w=0.97u l=0.18u
MI78 net89 SI VSS VSS n w=0.42u l=0.18u
MI80 net177 SE net89 VSS n w=0.42u l=0.18u
MI81 net066 D VSS VSS n w=1u l=0.18u
MI158-M_u4 XI158-net6 CDN VSS VSS n w=0.97u l=0.18u
MI158-M_u3 d3 d2 XI158-net6 VSS n w=0.97u l=0.18u
MI151_0-M_u2 QN net62 VSS VSS n w=1u l=0.18u
MI151_1-M_u2 QN net62 VSS VSS n w=1u l=0.18u
MI152_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI152_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI153-M_u2 net62 d3 VSS VSS n w=0.97u l=0.18u
MI85-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI165-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI32-M_u2 net101 INCPB VSS VSS n w=0.5u l=0.18u
MI158-M_u2 d3 CDN VDD VDD p w=0.42u l=0.18u
MI158-M_u1 d3 d2 VDD VDD p w=1.23u l=0.18u
MI151_0-M_u3 QN net62 VDD VDD p w=1.3u l=0.18u
MI151_1-M_u3 QN net62 VDD VDD p w=1.3u l=0.18u
MI152_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI152_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI153-M_u3 net62 d3 VDD VDD p w=0.97u l=0.18u
MI85-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI165-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI32-M_u3 net101 INCPB VDD VDD p w=0.685u l=0.18u
MI164 net177 SE net069 VDD p w=1.095u l=0.18u
MI155 net62 INCPB d2 VDD p w=0.42u l=0.18u
MI45 d0 net101 net166 VDD p w=0.42u l=0.18u
MI43 net166 d1 VDD VDD p w=0.42u l=0.18u
MI163 net177 net120 net142 VDD p w=0.42u l=0.18u
MI73 net069 D VDD VDD p w=1.37u l=0.18u
MI74 d0 INCPB net177 VDD p w=0.92u l=0.18u
MI75 net142 SI VDD VDD p w=0.42u l=0.18u
MI44 net166 CDN VDD VDD p w=0.42u l=0.18u
MI154 d1 net101 d2 VDD p w=0.62u l=0.18u
.ends
.subckt SDFND0BWP7T SI D SE CPN Q QN VDD VSS 
MI39 net13 net57 net083 VSS n w=1u l=0.18u
MI25 net65 INCPB d2 VSS n w=0.91u l=0.18u
MI13 net28 INCPB net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net55 net89 d2 VSS n w=0.42u l=0.18u
MU65 net28 net89 net13 VSS n w=0.57u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net083 D VSS VSS n w=1u l=0.18u
MI28-M_u2 net55 d3 VSS VSS n w=0.42u l=0.18u
MI30-M_u2 d3 d2 VSS VSS n w=0.5u l=0.18u
MI33-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI34-M_u2 QN net55 VSS VSS n w=0.5u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MI41-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MU85-M_u2 net89 INCPB VSS VSS n w=0.5u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net55 d3 VDD VDD p w=0.685u l=0.18u
MI30-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI33-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI34-M_u3 QN net55 VDD VDD p w=0.685u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MI41-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MU85-M_u3 net89 INCPB VDD VDD p w=0.685u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net55 INCPB d2 VDD p w=0.42u l=0.18u
MI40 net13 SE net110 VDD p w=1.18u l=0.18u
MI36 net65 net89 d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net110 D VDD VDD p w=1.18u l=0.18u
MU62 net28 INCPB net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 net89 net137 VDD p w=0.42u l=0.18u
.ends
.subckt SDFND1BWP7T SI D SE CPN Q QN VDD VSS 
MI39 net13 net57 net083 VSS n w=1u l=0.18u
MI25 net65 INCPB d2 VSS n w=0.91u l=0.18u
MI13 net28 INCPB net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net55 net89 d2 VSS n w=0.42u l=0.18u
MU65 net28 net89 net13 VSS n w=0.57u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net083 D VSS VSS n w=1u l=0.18u
MI28-M_u2 net55 d3 VSS VSS n w=0.42u l=0.18u
MI30-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI33-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI34-M_u2 QN net55 VSS VSS n w=0.94u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MI41-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MU85-M_u2 net89 INCPB VSS VSS n w=0.5u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net55 d3 VDD VDD p w=0.685u l=0.18u
MI30-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI33-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI34-M_u3 QN net55 VDD VDD p w=1.37u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MI41-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MU85-M_u3 net89 INCPB VDD VDD p w=0.685u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net55 INCPB d2 VDD p w=0.42u l=0.18u
MI40 net13 SE net110 VDD p w=1.18u l=0.18u
MI36 net65 net89 d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net110 D VDD VDD p w=1.18u l=0.18u
MU62 net28 INCPB net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 net89 net137 VDD p w=0.42u l=0.18u
.ends
.subckt SDFND2BWP7T SI D SE CPN Q QN VDD VSS 
MI39 net13 net57 net083 VSS n w=1u l=0.18u
MI25 net65 INCPB d2 VSS n w=0.91u l=0.18u
MI13 net28 INCPB net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net069 net89 d2 VSS n w=0.42u l=0.18u
MU65 net28 net89 net13 VSS n w=0.57u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net083 D VSS VSS n w=1u l=0.18u
MI28-M_u2 net069 d3 VSS VSS n w=1u l=0.18u
MI30-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI33_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI33_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI34_0-M_u2 QN net069 VSS VSS n w=1u l=0.18u
MI34_1-M_u2 QN net069 VSS VSS n w=1u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MI41-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MU85-M_u2 net89 INCPB VSS VSS n w=0.5u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net069 d3 VDD VDD p w=1.37u l=0.18u
MI30-M_u3 d3 d2 VDD VDD p w=1.23u l=0.18u
MI33_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI33_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI34_0-M_u3 QN net069 VDD VDD p w=1.3u l=0.18u
MI34_1-M_u3 QN net069 VDD VDD p w=1.3u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MI41-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MU85-M_u3 net89 INCPB VDD VDD p w=0.685u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net069 INCPB d2 VDD p w=0.42u l=0.18u
MI40 net13 SE net110 VDD p w=1.18u l=0.18u
MI36 net65 net89 d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net110 D VDD VDD p w=1.18u l=0.18u
MU62 net28 INCPB net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 net89 net137 VDD p w=0.42u l=0.18u
.ends
.subckt SDFNSND0BWP7T SI D SE CPN SDN Q QN VDD VSS 
MI91 d4 net95 d2 VSS n w=0.42u l=0.18u
MI92 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI101 net177 net120 net76 VSS n w=1u l=0.18u
MI48 net72 d1 VSS VSS n w=0.42u l=0.18u
MI47 net075 INCPB net72 VSS n w=0.42u l=0.18u
MI77 net075 net95 net177 VSS n w=0.91u l=0.18u
MI78 net79 SI VSS VSS n w=0.42u l=0.18u
MI80 net177 SE net79 VSS n w=0.42u l=0.18u
MI81 net76 D VSS VSS n w=1u l=0.18u
MI93-M_u4 XI93-net6 d3 VSS VSS n w=0.5u l=0.18u
MI93-M_u3 d4 SDN XI93-net6 VSS n w=0.5u l=0.18u
MI16-M_u4 XI16-net6 SDN VSS VSS n w=0.54u l=0.18u
MI16-M_u3 d1 net075 XI16-net6 VSS n w=0.54u l=0.18u
MI94-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI96-M_u2 d3 d2 VSS VSS n w=0.5u l=0.18u
MI103-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI32-M_u2 net95 INCPB VSS VSS n w=0.45u l=0.18u
MI95-M_u2 QN d4 VSS VSS n w=0.5u l=0.18u
MI93-M_u2 d4 d3 VDD VDD p w=0.685u l=0.18u
MI93-M_u1 d4 SDN VDD VDD p w=0.685u l=0.18u
MI16-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI16-M_u1 d1 net075 VDD VDD p w=0.97u l=0.18u
MI94-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI96-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI103-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI32-M_u3 net95 INCPB VDD VDD p w=0.685u l=0.18u
MI95-M_u3 QN d4 VDD VDD p w=0.685u l=0.18u
MI102 net177 SE net0108 VDD p w=1.095u l=0.18u
MI45 net075 net95 net126 VDD p w=0.42u l=0.18u
MI43 net126 d1 VDD VDD p w=0.42u l=0.18u
MI71 net177 net120 net131 VDD p w=0.42u l=0.18u
MI73 net0108 D VDD VDD p w=1.37u l=0.18u
MI74 net075 INCPB net177 VDD p w=0.92u l=0.18u
MI75 net131 SI VDD VDD p w=0.42u l=0.18u
MI97 d4 INCPB d2 VDD p w=0.42u l=0.18u
MI98 d1 net95 d2 VDD p w=1.34u l=0.18u
.ends
.subckt SDFNSND1BWP7T SI D SE CPN SDN Q QN VDD VSS 
MI91 d4 net95 d2 VSS n w=0.42u l=0.18u
MI92 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI101 net177 net120 net76 VSS n w=1u l=0.18u
MI48 net72 d1 VSS VSS n w=0.42u l=0.18u
MI47 net075 INCPB net72 VSS n w=0.42u l=0.18u
MI77 net075 net95 net177 VSS n w=0.91u l=0.18u
MI78 net79 SI VSS VSS n w=0.42u l=0.18u
MI80 net177 SE net79 VSS n w=0.42u l=0.18u
MI81 net76 D VSS VSS n w=1u l=0.18u
MI93-M_u4 XI93-net6 d3 VSS VSS n w=0.5u l=0.18u
MI93-M_u3 d4 SDN XI93-net6 VSS n w=0.5u l=0.18u
MI16-M_u4 XI16-net6 SDN VSS VSS n w=0.54u l=0.18u
MI16-M_u3 d1 net075 XI16-net6 VSS n w=0.54u l=0.18u
MI94-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI96-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI103-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI32-M_u2 net95 INCPB VSS VSS n w=0.45u l=0.18u
MI95-M_u2 QN d4 VSS VSS n w=1u l=0.18u
MI93-M_u2 d4 d3 VDD VDD p w=0.685u l=0.18u
MI93-M_u1 d4 SDN VDD VDD p w=0.685u l=0.18u
MI16-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI16-M_u1 d1 net075 VDD VDD p w=0.97u l=0.18u
MI94-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI96-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI103-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI32-M_u3 net95 INCPB VDD VDD p w=0.685u l=0.18u
MI95-M_u3 QN d4 VDD VDD p w=1.37u l=0.18u
MI102 net177 SE net0108 VDD p w=1.095u l=0.18u
MI45 net075 net95 net126 VDD p w=0.42u l=0.18u
MI43 net126 d1 VDD VDD p w=0.42u l=0.18u
MI71 net177 net120 net131 VDD p w=0.42u l=0.18u
MI73 net0108 D VDD VDD p w=1.37u l=0.18u
MI74 net075 INCPB net177 VDD p w=0.92u l=0.18u
MI75 net131 SI VDD VDD p w=0.42u l=0.18u
MI97 d4 INCPB d2 VDD p w=0.42u l=0.18u
MI98 d1 net95 d2 VDD p w=1.34u l=0.18u
.ends
.subckt SDFNSND2BWP7T SI D SE CPN SDN Q QN VDD VSS 
MI91 d4 net95 d2 VSS n w=0.42u l=0.18u
MI92 d1 INCPB d2 VSS n w=0.91u l=0.18u
MI101 net177 net120 net76 VSS n w=1u l=0.18u
MI48 net72 d1 VSS VSS n w=0.42u l=0.18u
MI47 net075 INCPB net72 VSS n w=0.42u l=0.18u
MI77 net075 net95 net177 VSS n w=0.91u l=0.18u
MI78 net79 SI VSS VSS n w=0.42u l=0.18u
MI80 net177 SE net79 VSS n w=0.42u l=0.18u
MI81 net76 D VSS VSS n w=1u l=0.18u
MI93-M_u4 XI93-net6 d3 VSS VSS n w=1u l=0.18u
MI93-M_u3 d4 SDN XI93-net6 VSS n w=1u l=0.18u
MI16-M_u4 XI16-net6 SDN VSS VSS n w=0.54u l=0.18u
MI16-M_u3 d1 net075 XI16-net6 VSS n w=0.54u l=0.18u
MI94_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI94_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI96-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI103-M_u2 INCPB CPN VSS VSS n w=0.5u l=0.18u
MI32-M_u2 net95 INCPB VSS VSS n w=0.45u l=0.18u
MI95_0-M_u2 QN d4 VSS VSS n w=1u l=0.18u
MI95_1-M_u2 QN d4 VSS VSS n w=1u l=0.18u
MI93-M_u2 d4 d3 VDD VDD p w=1.37u l=0.18u
MI93-M_u1 d4 SDN VDD VDD p w=0.535u l=0.18u
MI16-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI16-M_u1 d1 net075 VDD VDD p w=0.97u l=0.18u
MI94_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI94_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI96-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI103-M_u3 INCPB CPN VDD VDD p w=0.685u l=0.18u
MI32-M_u3 net95 INCPB VDD VDD p w=0.685u l=0.18u
MI95_0-M_u3 QN d4 VDD VDD p w=1.37u l=0.18u
MI95_1-M_u3 QN d4 VDD VDD p w=1.37u l=0.18u
MI102 net177 SE net0108 VDD p w=1.095u l=0.18u
MI45 net075 net95 net126 VDD p w=0.42u l=0.18u
MI43 net126 d1 VDD VDD p w=0.42u l=0.18u
MI71 net177 net120 net131 VDD p w=0.42u l=0.18u
MI73 net0108 D VDD VDD p w=1.37u l=0.18u
MI74 net075 INCPB net177 VDD p w=0.92u l=0.18u
MI75 net131 SI VDD VDD p w=0.42u l=0.18u
MI97 d4 INCPB d2 VDD p w=0.42u l=0.18u
MI98 d1 net95 d2 VDD p w=1.34u l=0.18u
.ends
.subckt SDFQD0BWP7T SI D SE CP Q VDD VSS 
MI39 net13 net57 net64 VSS n w=0.855u l=0.18u
MI25 net65 INCP d2 VSS n w=0.91u l=0.18u
MI13 net28 INCP net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net55 INCPB d2 VSS n w=0.42u l=0.18u
MU65 net28 INCPB net13 VSS n w=0.5u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net64 D VSS VSS n w=0.855u l=0.18u
MI28-M_u2 net55 d3 VSS VSS n w=0.42u l=0.18u
MI30-M_u2 d3 d2 VSS VSS n w=0.48u l=0.18u
MI33-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MU84-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net55 d3 VDD VDD p w=0.42u l=0.18u
MI30-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI33-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MU84-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net55 INCP d2 VDD p w=0.42u l=0.18u
MI36 net65 INCPB d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net0126 D VDD VDD p w=1.075u l=0.18u
MU62 net28 INCP net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 INCPB net137 VDD p w=0.42u l=0.18u
MI40 net13 SE net0126 VDD p w=1.075u l=0.18u
.ends
.subckt SDFQD1BWP7T SI D SE CP Q VDD VSS 
MI39 net13 net57 net64 VSS n w=1u l=0.18u
MI25 net65 INCP d2 VSS n w=0.91u l=0.18u
MI13 net28 INCP net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net55 INCPB d2 VSS n w=0.42u l=0.18u
MU65 net28 INCPB net13 VSS n w=0.5u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net64 D VSS VSS n w=1u l=0.18u
MI28-M_u2 net55 d3 VSS VSS n w=0.42u l=0.18u
MI30-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI33-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MU84-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net55 d3 VDD VDD p w=0.42u l=0.18u
MI30-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI33-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MU84-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net55 INCP d2 VDD p w=0.42u l=0.18u
MI36 net65 INCPB d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net0126 D VDD VDD p w=1.18u l=0.18u
MU62 net28 INCP net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 INCPB net137 VDD p w=0.42u l=0.18u
MI40 net13 SE net0126 VDD p w=1.18u l=0.18u
.ends
.subckt SDFQD2BWP7T SI D SE CP Q VDD VSS 
MI39 net13 net57 net64 VSS n w=1u l=0.18u
MI25 net65 INCP d2 VSS n w=0.91u l=0.18u
MI43 net054 d3 VSS VSS n w=0.42u l=0.18u
MI13 net28 INCP net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI42 d2 INCPB net054 VSS n w=0.42u l=0.18u
MU65 net28 INCPB net13 VSS n w=0.5u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net64 D VSS VSS n w=1u l=0.18u
MI30_0-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI30_1-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI33_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI33_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MU84-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI30_0-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI30_1-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI33_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI33_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MU84-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI44 net098 d3 VDD VDD p w=0.42u l=0.18u
MI45 d2 INCP net098 VDD p w=0.42u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI36 net65 INCPB d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net0126 D VDD VDD p w=1.18u l=0.18u
MU62 net28 INCP net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 INCPB net137 VDD p w=0.42u l=0.18u
MI40 net13 SE net0126 VDD p w=1.18u l=0.18u
.ends
.subckt SDFQND0BWP7T SI D SE CP QN VDD VSS 
MI39 net13 net57 net64 VSS n w=1u l=0.18u
MI25 net65 INCP d2 VSS n w=0.91u l=0.18u
MI13 net28 INCP net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net55 INCPB d2 VSS n w=0.42u l=0.18u
MU65 net28 INCPB net13 VSS n w=0.5u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net64 D VSS VSS n w=1u l=0.18u
MI28-M_u2 net55 d3 VSS VSS n w=0.5u l=0.18u
MI30-M_u2 d3 d2 VSS VSS n w=0.5u l=0.18u
MI34-M_u2 QN net55 VSS VSS n w=0.5u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MU84-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net55 d3 VDD VDD p w=0.685u l=0.18u
MI30-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI34-M_u3 QN net55 VDD VDD p w=0.685u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MU84-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net55 INCP d2 VDD p w=0.42u l=0.18u
MI36 net65 INCPB d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net0126 D VDD VDD p w=1.18u l=0.18u
MU62 net28 INCP net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 INCPB net137 VDD p w=0.42u l=0.18u
MI40 net13 SE net0126 VDD p w=1.18u l=0.18u
.ends
.subckt SDFQND1BWP7T SI D SE CP QN VDD VSS 
MI39 net13 net57 net64 VSS n w=1u l=0.18u
MI25 net65 INCP d2 VSS n w=0.91u l=0.18u
MI13 net28 INCP net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net55 INCPB d2 VSS n w=0.42u l=0.18u
MU65 net28 INCPB net13 VSS n w=0.5u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net64 D VSS VSS n w=1u l=0.18u
MI28-M_u2 net55 d3 VSS VSS n w=1u l=0.18u
MI30-M_u2 d3 d2 VSS VSS n w=0.5u l=0.18u
MI34-M_u2 QN net55 VSS VSS n w=1u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MU84-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net55 d3 VDD VDD p w=1.37u l=0.18u
MI30-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI34-M_u3 QN net55 VDD VDD p w=1.37u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MU84-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net55 INCP d2 VDD p w=0.42u l=0.18u
MI36 net65 INCPB d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net0126 D VDD VDD p w=1.18u l=0.18u
MU62 net28 INCP net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 INCPB net137 VDD p w=0.42u l=0.18u
MI40 net13 SE net0126 VDD p w=1.18u l=0.18u
.ends
.subckt SDFQND2BWP7T SI D SE CP QN VDD VSS 
MI39 net13 net57 net64 VSS n w=1u l=0.18u
MI25 net65 INCP d2 VSS n w=0.91u l=0.18u
MI13 net28 INCP net66 VSS n w=0.42u l=0.18u
MI14 net66 net65 VSS VSS n w=0.42u l=0.18u
MI26 net064 INCPB d2 VSS n w=0.42u l=0.18u
MU65 net28 INCPB net13 VSS n w=0.5u l=0.18u
MU67 net83 SI VSS VSS n w=0.42u l=0.18u
MU68 net13 SE net83 VSS n w=0.42u l=0.18u
MU63 net64 D VSS VSS n w=1u l=0.18u
MI28-M_u2 net064 d3 VSS VSS n w=1u l=0.18u
MI30-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI34_0-M_u2 QN net064 VSS VSS n w=1u l=0.18u
MI34_1-M_u2 QN net064 VSS VSS n w=1u l=0.18u
MU71-M_u2 net57 SE VSS VSS n w=0.5u l=0.18u
MU84-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MU72-M_u2 net65 net28 VSS VSS n w=0.54u l=0.18u
MI28-M_u3 net064 d3 VDD VDD p w=1.37u l=0.18u
MI30-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI34_0-M_u3 QN net064 VDD VDD p w=1.37u l=0.18u
MI34_1-M_u3 QN net064 VDD VDD p w=1.37u l=0.18u
MU71-M_u3 net57 SE VDD VDD p w=0.685u l=0.18u
MU84-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MU72-M_u3 net65 net28 VDD VDD p w=0.96u l=0.18u
MI11 net137 net65 VDD VDD p w=0.42u l=0.18u
MI35 net064 INCP d2 VDD p w=0.42u l=0.18u
MI36 net65 INCPB d2 VDD p w=1.34u l=0.18u
MU69 net13 net57 net132 VDD p w=0.42u l=0.18u
MU61 net0126 D VDD VDD p w=1.225u l=0.18u
MU62 net28 INCP net13 VDD p w=0.92u l=0.18u
MU70 net132 SI VDD VDD p w=0.42u l=0.18u
MI10 net28 INCPB net137 VDD p w=0.42u l=0.18u
MI40 net13 SE net0126 VDD p w=1.225u l=0.18u
.ends
.subckt SDFSND0BWP7T SI D SE CP SDN Q QN VDD VSS 
MI91 net063 INCPB d2 VSS n w=0.42u l=0.18u
MI92 d1 INCP d2 VSS n w=0.91u l=0.18u
MI102 net104 net120 net75 VSS n w=1u l=0.18u
MI48 net72 d1 VSS VSS n w=0.42u l=0.18u
MI47 net077 INCP net72 VSS n w=0.42u l=0.18u
MI77 net077 INCPB net104 VSS n w=0.83u l=0.18u
MI78 net79 SI VSS VSS n w=0.42u l=0.18u
MI80 net104 SE net79 VSS n w=0.42u l=0.18u
MI81 net75 D VSS VSS n w=1u l=0.18u
MI93-M_u4 XI93-net6 d3 VSS VSS n w=0.5u l=0.18u
MI93-M_u3 net063 SDN XI93-net6 VSS n w=0.5u l=0.18u
MI16-M_u4 XI16-net6 SDN VSS VSS n w=0.54u l=0.18u
MI16-M_u3 d1 net077 XI16-net6 VSS n w=0.54u l=0.18u
MI104-M_u2 QN net063 VSS VSS n w=0.5u l=0.18u
MI94-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI96-M_u2 d3 d2 VSS VSS n w=0.5u l=0.18u
MI103-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI93-M_u2 net063 d3 VDD VDD p w=0.685u l=0.18u
MI93-M_u1 net063 SDN VDD VDD p w=0.685u l=0.18u
MI16-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI16-M_u1 d1 net077 VDD VDD p w=0.97u l=0.18u
MI104-M_u3 QN net063 VDD VDD p w=0.685u l=0.18u
MI94-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI96-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI103-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI45 net077 INCPB net126 VDD p w=0.42u l=0.18u
MI43 net126 d1 VDD VDD p w=0.42u l=0.18u
MI71 net104 net120 net131 VDD p w=0.42u l=0.18u
MI73 net75 D VDD VDD p w=1.37u l=0.18u
MI74 net077 INCP net104 VDD p w=0.92u l=0.18u
MI75 net131 SI VDD VDD p w=0.42u l=0.18u
MI101 net104 SE net75 VDD p w=1.095u l=0.18u
MI97 net063 INCP d2 VDD p w=0.42u l=0.18u
MI98 d1 INCPB d2 VDD p w=1.34u l=0.18u
.ends
.subckt SDFSND1BWP7T SI D SE CP SDN Q QN VDD VSS 
MI91 net063 INCPB d2 VSS n w=0.42u l=0.18u
MI92 d1 INCP d2 VSS n w=0.91u l=0.18u
MI102 net104 net120 net75 VSS n w=1u l=0.18u
MI48 net72 d1 VSS VSS n w=0.42u l=0.18u
MI47 net077 INCP net72 VSS n w=0.42u l=0.18u
MI77 net077 INCPB net104 VSS n w=0.83u l=0.18u
MI78 net79 SI VSS VSS n w=0.42u l=0.18u
MI80 net104 SE net79 VSS n w=0.42u l=0.18u
MI81 net75 D VSS VSS n w=1u l=0.18u
MI93-M_u4 XI93-net6 d3 VSS VSS n w=0.5u l=0.18u
MI93-M_u3 net063 SDN XI93-net6 VSS n w=0.5u l=0.18u
MI16-M_u4 XI16-net6 SDN VSS VSS n w=0.54u l=0.18u
MI16-M_u3 d1 net077 XI16-net6 VSS n w=0.54u l=0.18u
MI104-M_u2 QN net063 VSS VSS n w=1u l=0.18u
MI94-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI96-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI103-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI93-M_u2 net063 d3 VDD VDD p w=0.685u l=0.18u
MI93-M_u1 net063 SDN VDD VDD p w=0.685u l=0.18u
MI16-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI16-M_u1 d1 net077 VDD VDD p w=0.97u l=0.18u
MI104-M_u3 QN net063 VDD VDD p w=1.37u l=0.18u
MI94-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI96-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI103-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI45 net077 INCPB net126 VDD p w=0.42u l=0.18u
MI43 net126 d1 VDD VDD p w=0.42u l=0.18u
MI71 net104 net120 net131 VDD p w=0.42u l=0.18u
MI73 net75 D VDD VDD p w=1.37u l=0.18u
MI74 net077 INCP net104 VDD p w=0.92u l=0.18u
MI75 net131 SI VDD VDD p w=0.42u l=0.18u
MI101 net104 SE net75 VDD p w=1.095u l=0.18u
MI97 net063 INCP d2 VDD p w=0.42u l=0.18u
MI98 d1 INCPB d2 VDD p w=1.34u l=0.18u
.ends
.subckt SDFSND2BWP7T SI D SE CP SDN Q QN VDD VSS 
MI91 net063 INCPB d2 VSS n w=0.42u l=0.18u
MI92 d1 INCP d2 VSS n w=0.91u l=0.18u
MI102 net104 net120 net75 VSS n w=1u l=0.18u
MI48 net72 d1 VSS VSS n w=0.42u l=0.18u
MI47 net077 INCP net72 VSS n w=0.42u l=0.18u
MI77 net077 INCPB net104 VSS n w=0.83u l=0.18u
MI78 net79 SI VSS VSS n w=0.42u l=0.18u
MI80 net104 SE net79 VSS n w=0.42u l=0.18u
MI81 net75 D VSS VSS n w=1u l=0.18u
MI93-M_u4 XI93-net6 d3 VSS VSS n w=1u l=0.18u
MI93-M_u3 net063 SDN XI93-net6 VSS n w=1u l=0.18u
MI16-M_u4 XI16-net6 SDN VSS VSS n w=0.54u l=0.18u
MI16-M_u3 d1 net077 XI16-net6 VSS n w=0.54u l=0.18u
MI104_0-M_u2 QN net063 VSS VSS n w=1u l=0.18u
MI104_1-M_u2 QN net063 VSS VSS n w=1u l=0.18u
MI94_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI94_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI96-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI103-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI93-M_u2 net063 d3 VDD VDD p w=1.37u l=0.18u
MI93-M_u1 net063 SDN VDD VDD p w=0.685u l=0.18u
MI16-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI16-M_u1 d1 net077 VDD VDD p w=0.97u l=0.18u
MI104_0-M_u3 QN net063 VDD VDD p w=1.37u l=0.18u
MI104_1-M_u3 QN net063 VDD VDD p w=1.37u l=0.18u
MI94_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI94_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI96-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI103-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI45 net077 INCPB net126 VDD p w=0.42u l=0.18u
MI43 net126 d1 VDD VDD p w=0.42u l=0.18u
MI71 net104 net120 net131 VDD p w=0.42u l=0.18u
MI73 net75 D VDD VDD p w=1.37u l=0.18u
MI74 net077 INCP net104 VDD p w=0.92u l=0.18u
MI75 net131 SI VDD VDD p w=0.42u l=0.18u
MI101 net104 SE net75 VDD p w=1.095u l=0.18u
MI97 net063 INCP d2 VDD p w=0.42u l=0.18u
MI98 d1 INCPB d2 VDD p w=1.34u l=0.18u
.ends
.subckt SDFSNQD0BWP7T SI D SE CP SDN Q VDD VSS 
MI91 net063 INCPB d2 VSS n w=0.42u l=0.18u
MI92 d1 INCP d2 VSS n w=0.91u l=0.18u
MI102 net104 net120 net75 VSS n w=1u l=0.18u
MI48 net72 d1 VSS VSS n w=0.42u l=0.18u
MI47 net077 INCP net72 VSS n w=0.42u l=0.18u
MI77 net077 INCPB net104 VSS n w=0.83u l=0.18u
MI78 net79 SI VSS VSS n w=0.42u l=0.18u
MI80 net104 SE net79 VSS n w=0.42u l=0.18u
MI81 net75 D VSS VSS n w=1u l=0.18u
MI93-M_u4 XI93-net6 d3 VSS VSS n w=0.5u l=0.18u
MI93-M_u3 net063 SDN XI93-net6 VSS n w=0.5u l=0.18u
MI16-M_u4 XI16-net6 SDN VSS VSS n w=0.54u l=0.18u
MI16-M_u3 d1 net077 XI16-net6 VSS n w=0.54u l=0.18u
MI94-M_u2 Q d3 VSS VSS n w=0.5u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI96-M_u2 d3 d2 VSS VSS n w=0.5u l=0.18u
MI103-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI93-M_u2 net063 d3 VDD VDD p w=0.685u l=0.18u
MI93-M_u1 net063 SDN VDD VDD p w=0.685u l=0.18u
MI16-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI16-M_u1 d1 net077 VDD VDD p w=0.97u l=0.18u
MI94-M_u3 Q d3 VDD VDD p w=0.685u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI96-M_u3 d3 d2 VDD VDD p w=0.685u l=0.18u
MI103-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI45 net077 INCPB net126 VDD p w=0.42u l=0.18u
MI43 net126 d1 VDD VDD p w=0.42u l=0.18u
MI71 net104 net120 net131 VDD p w=0.42u l=0.18u
MI73 net75 D VDD VDD p w=1.37u l=0.18u
MI74 net077 INCP net104 VDD p w=0.92u l=0.18u
MI75 net131 SI VDD VDD p w=0.42u l=0.18u
MI101 net104 SE net75 VDD p w=1.095u l=0.18u
MI97 net063 INCP d2 VDD p w=0.42u l=0.18u
MI98 d1 INCPB d2 VDD p w=1.34u l=0.18u
.ends
.subckt SDFSNQD1BWP7T SI D SE CP SDN Q VDD VSS 
MI91 net063 INCPB d2 VSS n w=0.42u l=0.18u
MI92 d1 INCP d2 VSS n w=0.91u l=0.18u
MI102 net104 net120 net75 VSS n w=1u l=0.18u
MI48 net72 d1 VSS VSS n w=0.42u l=0.18u
MI47 net077 INCP net72 VSS n w=0.42u l=0.18u
MI77 net077 INCPB net104 VSS n w=0.83u l=0.18u
MI78 net79 SI VSS VSS n w=0.42u l=0.18u
MI80 net104 SE net79 VSS n w=0.42u l=0.18u
MI81 net75 D VSS VSS n w=1u l=0.18u
MI93-M_u4 XI93-net6 d3 VSS VSS n w=0.5u l=0.18u
MI93-M_u3 net063 SDN XI93-net6 VSS n w=0.5u l=0.18u
MI16-M_u4 XI16-net6 SDN VSS VSS n w=0.54u l=0.18u
MI16-M_u3 d1 net077 XI16-net6 VSS n w=0.54u l=0.18u
MI94-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI96-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI103-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI93-M_u2 net063 d3 VDD VDD p w=0.685u l=0.18u
MI93-M_u1 net063 SDN VDD VDD p w=0.685u l=0.18u
MI16-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI16-M_u1 d1 net077 VDD VDD p w=0.97u l=0.18u
MI94-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI96-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI103-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI45 net077 INCPB net126 VDD p w=0.42u l=0.18u
MI43 net126 d1 VDD VDD p w=0.42u l=0.18u
MI71 net104 net120 net131 VDD p w=0.42u l=0.18u
MI73 net75 D VDD VDD p w=1.37u l=0.18u
MI74 net077 INCP net104 VDD p w=0.92u l=0.18u
MI75 net131 SI VDD VDD p w=0.42u l=0.18u
MI101 net104 SE net75 VDD p w=1.095u l=0.18u
MI97 net063 INCP d2 VDD p w=0.42u l=0.18u
MI98 d1 INCPB d2 VDD p w=1.34u l=0.18u
.ends
.subckt SDFSNQD2BWP7T SI D SE CP SDN Q VDD VSS 
MI91 net063 INCPB d2 VSS n w=0.42u l=0.18u
MI92 d1 INCP d2 VSS n w=0.91u l=0.18u
MI102 net104 net120 net75 VSS n w=1u l=0.18u
MI48 net72 d1 VSS VSS n w=0.42u l=0.18u
MI47 net077 INCP net72 VSS n w=0.42u l=0.18u
MI77 net077 INCPB net104 VSS n w=0.83u l=0.18u
MI78 net79 SI VSS VSS n w=0.42u l=0.18u
MI80 net104 SE net79 VSS n w=0.42u l=0.18u
MI81 net75 D VSS VSS n w=1u l=0.18u
MI93-M_u4 XI93-net6 d3 VSS VSS n w=0.42u l=0.18u
MI93-M_u3 net063 SDN XI93-net6 VSS n w=0.42u l=0.18u
MI16-M_u4 XI16-net6 SDN VSS VSS n w=0.54u l=0.18u
MI16-M_u3 d1 net077 XI16-net6 VSS n w=0.54u l=0.18u
MI94_0-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI94_1-M_u2 Q d3 VSS VSS n w=1u l=0.18u
MI82-M_u2 net120 SE VSS VSS n w=0.5u l=0.18u
MI96-M_u2 d3 d2 VSS VSS n w=1u l=0.18u
MI103-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI32-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI93-M_u2 net063 d3 VDD VDD p w=0.685u l=0.18u
MI93-M_u1 net063 SDN VDD VDD p w=0.685u l=0.18u
MI16-M_u2 d1 SDN VDD VDD p w=0.42u l=0.18u
MI16-M_u1 d1 net077 VDD VDD p w=0.97u l=0.18u
MI94_0-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI94_1-M_u3 Q d3 VDD VDD p w=1.37u l=0.18u
MI82-M_u3 net120 SE VDD VDD p w=0.685u l=0.18u
MI96-M_u3 d3 d2 VDD VDD p w=1.37u l=0.18u
MI103-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI32-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI45 net077 INCPB net126 VDD p w=0.42u l=0.18u
MI43 net126 d1 VDD VDD p w=0.42u l=0.18u
MI71 net104 net120 net131 VDD p w=0.42u l=0.18u
MI73 net75 D VDD VDD p w=1.37u l=0.18u
MI74 net077 INCP net104 VDD p w=0.92u l=0.18u
MI75 net131 SI VDD VDD p w=0.42u l=0.18u
MI101 net104 SE net75 VDD p w=1.095u l=0.18u
MI97 net063 INCP d2 VDD p w=0.42u l=0.18u
MI98 d1 INCPB d2 VDD p w=1.34u l=0.18u
.ends
.subckt SDFXD0BWP7T DA DB SA SI SE CP Q QN VDD VSS 
MI178 d1 INCP net69 VSS n w=0.91u l=0.18u
MI179 net67 INCPB net69 VSS n w=0.42u l=0.18u
MI189 net163 net318 net0112 VSS n w=1u l=0.18u
MI119 net79 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net79 VSS n w=0.42u l=0.18u
MI162 net112 SI VSS VSS n w=0.42u l=0.18u
MI168 net250 net0124 net95 VSS n w=1u l=0.18u
MI167 net95 DB VSS VSS n w=1u l=0.18u
MI166 net250 SA net101 VSS n w=0.52u l=0.18u
MI165 net101 DA VSS VSS n w=0.52u l=0.18u
MI164 d0 INCPB net163 VSS n w=0.91u l=0.18u
MI160 net0112 net314 VSS VSS n w=1u l=0.18u
MI161 net163 SE net112 VSS n w=0.42u l=0.18u
MI180-M_u2 net67 net107 VSS VSS n w=0.42u l=0.18u
MI181-M_u2 net107 net69 VSS VSS n w=0.5u l=0.18u
MI182-M_u2 Q net107 VSS VSS n w=0.5u l=0.18u
MI183-M_u2 QN net67 VSS VSS n w=0.5u l=0.18u
MI171-M_u2 net314 net250 VSS VSS n w=1u l=0.18u
MI170-M_u2 net0124 SA VSS VSS n w=0.5u l=0.18u
MI169-M_u2 net318 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI190-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI123-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI180-M_u3 net67 net107 VDD VDD p w=0.685u l=0.18u
MI181-M_u3 net107 net69 VDD VDD p w=0.685u l=0.18u
MI182-M_u3 Q net107 VDD VDD p w=0.685u l=0.18u
MI183-M_u3 QN net67 VDD VDD p w=0.685u l=0.18u
MI171-M_u3 net314 net250 VDD VDD p w=1.36u l=0.18u
MI170-M_u3 net0124 SA VDD VDD p w=0.685u l=0.18u
MI169-M_u3 net318 SE VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI190-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI123-M_u3 d1 d0 VDD VDD p w=0.96u l=0.18u
MI184 net67 INCP net69 VDD p w=0.42u l=0.18u
MI185 d1 INCPB net69 VDD p w=1.34u l=0.18u
MI188 net163 SE net208 VDD p w=1.095u l=0.18u
MI102 net144 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net144 VDD p w=0.42u l=0.18u
MI149 net167 SI VDD VDD p w=0.42u l=0.18u
MI150 net208 net314 VDD VDD p w=1.23u l=0.18u
MI157 net250 net0124 net161 VDD p w=0.725u l=0.18u
MI152 net163 net318 net167 VDD p w=0.42u l=0.18u
MI153 d0 INCP net163 VDD p w=0.92u l=0.18u
MI154 net250 SA net173 VDD p w=1.095u l=0.18u
MI155 net161 DA VDD VDD p w=0.725u l=0.18u
MI156 net173 DB VDD VDD p w=1.36u l=0.18u
.ends
.subckt SDFXD1BWP7T DA DB SA SI SE CP Q QN VDD VSS 
MI178 d1 INCP net69 VSS n w=0.91u l=0.18u
MI179 net67 INCPB net69 VSS n w=0.42u l=0.18u
MI189 net163 net318 net0112 VSS n w=1u l=0.18u
MI119 net79 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net79 VSS n w=0.42u l=0.18u
MI162 net112 SI VSS VSS n w=0.42u l=0.18u
MI168 net250 net0124 net95 VSS n w=1u l=0.18u
MI167 net95 DB VSS VSS n w=1u l=0.18u
MI166 net250 SA net101 VSS n w=0.52u l=0.18u
MI165 net101 DA VSS VSS n w=0.52u l=0.18u
MI164 d0 INCPB net163 VSS n w=0.91u l=0.18u
MI160 net0112 net314 VSS VSS n w=1u l=0.18u
MI161 net163 SE net112 VSS n w=0.42u l=0.18u
MI180-M_u2 net67 net107 VSS VSS n w=0.42u l=0.18u
MI181-M_u2 net107 net69 VSS VSS n w=1u l=0.18u
MI182-M_u2 Q net107 VSS VSS n w=1u l=0.18u
MI183-M_u2 QN net67 VSS VSS n w=0.94u l=0.18u
MI171-M_u2 net314 net250 VSS VSS n w=1u l=0.18u
MI170-M_u2 net0124 SA VSS VSS n w=0.5u l=0.18u
MI169-M_u2 net318 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI190-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI123-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI180-M_u3 net67 net107 VDD VDD p w=0.685u l=0.18u
MI181-M_u3 net107 net69 VDD VDD p w=1.37u l=0.18u
MI182-M_u3 Q net107 VDD VDD p w=1.37u l=0.18u
MI183-M_u3 QN net67 VDD VDD p w=1.37u l=0.18u
MI171-M_u3 net314 net250 VDD VDD p w=1.36u l=0.18u
MI170-M_u3 net0124 SA VDD VDD p w=0.685u l=0.18u
MI169-M_u3 net318 SE VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI190-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI123-M_u3 d1 d0 VDD VDD p w=0.96u l=0.18u
MI184 net67 INCP net69 VDD p w=0.42u l=0.18u
MI185 d1 INCPB net69 VDD p w=1.34u l=0.18u
MI188 net163 SE net208 VDD p w=1.095u l=0.18u
MI102 net144 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net144 VDD p w=0.42u l=0.18u
MI149 net167 SI VDD VDD p w=0.42u l=0.18u
MI150 net208 net314 VDD VDD p w=1.23u l=0.18u
MI157 net250 net0124 net161 VDD p w=0.725u l=0.18u
MI152 net163 net318 net167 VDD p w=0.42u l=0.18u
MI153 d0 INCP net163 VDD p w=0.92u l=0.18u
MI154 net250 SA net173 VDD p w=1.095u l=0.18u
MI155 net161 DA VDD VDD p w=0.725u l=0.18u
MI156 net173 DB VDD VDD p w=1.36u l=0.18u
.ends
.subckt SDFXD2BWP7T DA DB SA SI SE CP Q QN VDD VSS 
MI178 d1 INCP net69 VSS n w=0.91u l=0.18u
MI179 net67 INCPB net69 VSS n w=0.42u l=0.18u
MI189 net163 net318 net0112 VSS n w=1u l=0.18u
MI119 net79 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net79 VSS n w=0.42u l=0.18u
MI162 net112 SI VSS VSS n w=0.42u l=0.18u
MI168 net250 net0124 net95 VSS n w=1u l=0.18u
MI167 net95 DB VSS VSS n w=1u l=0.18u
MI166 net250 SA net101 VSS n w=0.52u l=0.18u
MI165 net101 DA VSS VSS n w=0.52u l=0.18u
MI164 d0 INCPB net163 VSS n w=0.91u l=0.18u
MI160 net0112 net314 VSS VSS n w=1u l=0.18u
MI161 net163 SE net112 VSS n w=0.42u l=0.18u
MI180-M_u2 net67 net0117 VSS VSS n w=1u l=0.18u
MI181-M_u2 net0117 net69 VSS VSS n w=1u l=0.18u
MI182_0-M_u2 Q net0117 VSS VSS n w=1u l=0.18u
MI182_1-M_u2 Q net0117 VSS VSS n w=1u l=0.18u
MI183_0-M_u2 QN net67 VSS VSS n w=1u l=0.18u
MI183_1-M_u2 QN net67 VSS VSS n w=1u l=0.18u
MI171-M_u2 net314 net250 VSS VSS n w=1u l=0.18u
MI170-M_u2 net0124 SA VSS VSS n w=0.5u l=0.18u
MI169-M_u2 net318 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI190-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI123-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI180-M_u3 net67 net0117 VDD VDD p w=1.37u l=0.18u
MI181-M_u3 net0117 net69 VDD VDD p w=1.23u l=0.18u
MI182_0-M_u3 Q net0117 VDD VDD p w=1.37u l=0.18u
MI182_1-M_u3 Q net0117 VDD VDD p w=1.37u l=0.18u
MI183_0-M_u3 QN net67 VDD VDD p w=1.3u l=0.18u
MI183_1-M_u3 QN net67 VDD VDD p w=1.3u l=0.18u
MI171-M_u3 net314 net250 VDD VDD p w=1.36u l=0.18u
MI170-M_u3 net0124 SA VDD VDD p w=0.685u l=0.18u
MI169-M_u3 net318 SE VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI190-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI123-M_u3 d1 d0 VDD VDD p w=0.96u l=0.18u
MI184 net67 INCP net69 VDD p w=0.42u l=0.18u
MI185 d1 INCPB net69 VDD p w=1.34u l=0.18u
MI188 net163 SE net208 VDD p w=1.095u l=0.18u
MI102 net144 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net144 VDD p w=0.42u l=0.18u
MI149 net167 SI VDD VDD p w=0.42u l=0.18u
MI150 net208 net314 VDD VDD p w=1.23u l=0.18u
MI157 net250 net0124 net161 VDD p w=0.725u l=0.18u
MI152 net163 net318 net167 VDD p w=0.42u l=0.18u
MI153 d0 INCP net163 VDD p w=0.92u l=0.18u
MI154 net250 SA net173 VDD p w=1.095u l=0.18u
MI155 net161 DA VDD VDD p w=0.725u l=0.18u
MI156 net173 DB VDD VDD p w=1.36u l=0.18u
.ends
.subckt SDFXQD0BWP7T DA DB SA SI SE CP Q VDD VSS 
MI178 d1 INCP net69 VSS n w=0.91u l=0.18u
MI179 net67 INCPB net69 VSS n w=0.42u l=0.18u
MI189 net163 net318 net0112 VSS n w=1u l=0.18u
MI119 net79 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net79 VSS n w=0.42u l=0.18u
MI162 net112 SI VSS VSS n w=0.42u l=0.18u
MI168 net250 net0124 net95 VSS n w=1u l=0.18u
MI167 net95 DB VSS VSS n w=1u l=0.18u
MI166 net250 SA net101 VSS n w=0.52u l=0.18u
MI165 net101 DA VSS VSS n w=0.52u l=0.18u
MI164 d0 INCPB net163 VSS n w=0.91u l=0.18u
MI160 net0112 net314 VSS VSS n w=1u l=0.18u
MI161 net163 SE net112 VSS n w=0.42u l=0.18u
MI180-M_u2 net67 net107 VSS VSS n w=0.42u l=0.18u
MI181-M_u2 net107 net69 VSS VSS n w=0.5u l=0.18u
MI182-M_u2 Q net107 VSS VSS n w=0.5u l=0.18u
MI171-M_u2 net314 net250 VSS VSS n w=1u l=0.18u
MI170-M_u2 net0124 SA VSS VSS n w=0.5u l=0.18u
MI169-M_u2 net318 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI190-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI123-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI180-M_u3 net67 net107 VDD VDD p w=0.42u l=0.18u
MI181-M_u3 net107 net69 VDD VDD p w=0.685u l=0.18u
MI182-M_u3 Q net107 VDD VDD p w=0.685u l=0.18u
MI171-M_u3 net314 net250 VDD VDD p w=1.36u l=0.18u
MI170-M_u3 net0124 SA VDD VDD p w=0.685u l=0.18u
MI169-M_u3 net318 SE VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI190-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI123-M_u3 d1 d0 VDD VDD p w=0.96u l=0.18u
MI184 net67 INCP net69 VDD p w=0.42u l=0.18u
MI185 d1 INCPB net69 VDD p w=1.34u l=0.18u
MI188 net163 SE net208 VDD p w=1.095u l=0.18u
MI102 net144 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net144 VDD p w=0.42u l=0.18u
MI149 net167 SI VDD VDD p w=0.42u l=0.18u
MI150 net208 net314 VDD VDD p w=1.23u l=0.18u
MI157 net250 net0124 net161 VDD p w=0.725u l=0.18u
MI152 net163 net318 net167 VDD p w=0.42u l=0.18u
MI153 d0 INCP net163 VDD p w=0.92u l=0.18u
MI154 net250 SA net173 VDD p w=1.095u l=0.18u
MI155 net161 DA VDD VDD p w=0.725u l=0.18u
MI156 net173 DB VDD VDD p w=1.36u l=0.18u
.ends
.subckt SDFXQD1BWP7T DA DB SA SI SE CP Q VDD VSS 
MI178 d1 INCP net69 VSS n w=0.91u l=0.18u
MI179 net67 INCPB net69 VSS n w=0.42u l=0.18u
MI189 net163 net318 net0112 VSS n w=1u l=0.18u
MI119 net79 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net79 VSS n w=0.42u l=0.18u
MI162 net112 SI VSS VSS n w=0.42u l=0.18u
MI168 net250 net0124 net95 VSS n w=1u l=0.18u
MI167 net95 DB VSS VSS n w=1u l=0.18u
MI166 net250 SA net101 VSS n w=0.52u l=0.18u
MI165 net101 DA VSS VSS n w=0.52u l=0.18u
MI164 d0 INCPB net163 VSS n w=0.91u l=0.18u
MI160 net0112 net314 VSS VSS n w=1u l=0.18u
MI161 net163 SE net112 VSS n w=0.42u l=0.18u
MI180-M_u2 net67 net107 VSS VSS n w=0.42u l=0.18u
MI181-M_u2 net107 net69 VSS VSS n w=1u l=0.18u
MI182-M_u2 Q net107 VSS VSS n w=1u l=0.18u
MI171-M_u2 net314 net250 VSS VSS n w=1u l=0.18u
MI170-M_u2 net0124 SA VSS VSS n w=0.5u l=0.18u
MI169-M_u2 net318 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI190-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI123-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI180-M_u3 net67 net107 VDD VDD p w=0.42u l=0.18u
MI181-M_u3 net107 net69 VDD VDD p w=1.37u l=0.18u
MI182-M_u3 Q net107 VDD VDD p w=1.37u l=0.18u
MI171-M_u3 net314 net250 VDD VDD p w=1.36u l=0.18u
MI170-M_u3 net0124 SA VDD VDD p w=0.685u l=0.18u
MI169-M_u3 net318 SE VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI190-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI123-M_u3 d1 d0 VDD VDD p w=0.96u l=0.18u
MI184 net67 INCP net69 VDD p w=0.42u l=0.18u
MI185 d1 INCPB net69 VDD p w=1.34u l=0.18u
MI188 net163 SE net208 VDD p w=1.095u l=0.18u
MI102 net144 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net144 VDD p w=0.42u l=0.18u
MI149 net167 SI VDD VDD p w=0.42u l=0.18u
MI150 net208 net314 VDD VDD p w=1.23u l=0.18u
MI157 net250 net0124 net161 VDD p w=0.725u l=0.18u
MI152 net163 net318 net167 VDD p w=0.42u l=0.18u
MI153 d0 INCP net163 VDD p w=0.92u l=0.18u
MI154 net250 SA net173 VDD p w=1.095u l=0.18u
MI155 net161 DA VDD VDD p w=0.725u l=0.18u
MI156 net173 DB VDD VDD p w=1.36u l=0.18u
.ends
.subckt SDFXQD2BWP7T DA DB SA SI SE CP Q VDD VSS 
MI178 d1 INCP net69 VSS n w=0.91u l=0.18u
MI189 net163 net318 net0112 VSS n w=1u l=0.18u
MI192 net075 net0117 VSS VSS n w=0.42u l=0.18u
MI119 net79 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net79 VSS n w=0.42u l=0.18u
MI193 net69 INCPB net075 VSS n w=0.42u l=0.18u
MI162 net112 SI VSS VSS n w=0.42u l=0.18u
MI168 net250 net0124 net95 VSS n w=1u l=0.18u
MI167 net95 DB VSS VSS n w=1u l=0.18u
MI166 net250 SA net101 VSS n w=0.52u l=0.18u
MI165 net101 DA VSS VSS n w=0.52u l=0.18u
MI164 d0 INCPB net163 VSS n w=0.91u l=0.18u
MI160 net0112 net314 VSS VSS n w=1u l=0.18u
MI161 net163 SE net112 VSS n w=0.42u l=0.18u
MI181_0-M_u2 net0117 net69 VSS VSS n w=1u l=0.18u
MI181_1-M_u2 net0117 net69 VSS VSS n w=1u l=0.18u
MI182_0-M_u2 Q net0117 VSS VSS n w=1u l=0.18u
MI182_1-M_u2 Q net0117 VSS VSS n w=1u l=0.18u
MI171-M_u2 net314 net250 VSS VSS n w=1u l=0.18u
MI170-M_u2 net0124 SA VSS VSS n w=0.5u l=0.18u
MI169-M_u2 net318 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI190-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI123-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI181_0-M_u3 net0117 net69 VDD VDD p w=1.37u l=0.18u
MI181_1-M_u3 net0117 net69 VDD VDD p w=1.37u l=0.18u
MI182_0-M_u3 Q net0117 VDD VDD p w=1.37u l=0.18u
MI182_1-M_u3 Q net0117 VDD VDD p w=1.37u l=0.18u
MI171-M_u3 net314 net250 VDD VDD p w=1.36u l=0.18u
MI170-M_u3 net0124 SA VDD VDD p w=0.685u l=0.18u
MI169-M_u3 net318 SE VDD VDD p w=0.685u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI190-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI123-M_u3 d1 d0 VDD VDD p w=0.96u l=0.18u
MI195 net69 INCP net0135 VDD p w=0.42u l=0.18u
MI194 net0135 net0117 VDD VDD p w=0.42u l=0.18u
MI185 d1 INCPB net69 VDD p w=1.34u l=0.18u
MI188 net163 SE net208 VDD p w=1.095u l=0.18u
MI102 net144 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net144 VDD p w=0.42u l=0.18u
MI149 net167 SI VDD VDD p w=0.42u l=0.18u
MI150 net208 net314 VDD VDD p w=1.23u l=0.18u
MI157 net250 net0124 net161 VDD p w=0.725u l=0.18u
MI152 net163 net318 net167 VDD p w=0.42u l=0.18u
MI153 d0 INCP net163 VDD p w=0.92u l=0.18u
MI154 net250 SA net173 VDD p w=1.095u l=0.18u
MI155 net161 DA VDD VDD p w=0.725u l=0.18u
MI156 net173 DB VDD VDD p w=1.36u l=0.18u
.ends
.subckt SEDFCND0BWP7T E SE CP SI D CDN Q QN VDD VSS 
MI239 net080 net083 net079 VSS n w=0.52u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net92 d1 VSS VSS n w=0.42u l=0.18u
MI119 net95 CDN net92 VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net083 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.52u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI183-M_u4 XI183-net6 CDN VSS VSS n w=0.93u l=0.18u
MI183-M_u3 d2 net084 XI183-net6 VSS n w=1u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI189-M_u2 QN net083 VSS VSS n w=0.5u l=0.18u
MI175-M_u2 Q d2 VSS VSS n w=0.5u l=0.18u
MI177-M_u2 net083 d2 VSS VSS n w=0.42u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI183-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI183-M_u1 d2 net084 VDD VDD p w=1.03u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI189-M_u3 QN net083 VDD VDD p w=0.685u l=0.18u
MI175-M_u3 Q d2 VDD VDD p w=0.685u l=0.18u
MI177-M_u3 net083 d2 VDD VDD p w=0.685u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.42u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI101 net83 CDN VDD VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net083 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=0.62u l=0.18u
MI233 net0147 net083 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.78u l=0.18u
.ends
.subckt SEDFCND1BWP7T E SE CP SI D CDN Q QN VDD VSS 
MI239 net080 net083 net079 VSS n w=0.52u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net92 d1 VSS VSS n w=0.42u l=0.18u
MI119 net95 CDN net92 VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net083 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.52u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI183-M_u4 XI183-net6 CDN VSS VSS n w=0.93u l=0.18u
MI183-M_u3 d2 net084 XI183-net6 VSS n w=1u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI189-M_u2 QN net083 VSS VSS n w=0.94u l=0.18u
MI175-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI177-M_u2 net083 d2 VSS VSS n w=0.42u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI183-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI183-M_u1 d2 net084 VDD VDD p w=1.03u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI189-M_u3 QN net083 VDD VDD p w=1.37u l=0.18u
MI175-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI177-M_u3 net083 d2 VDD VDD p w=0.685u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.42u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI101 net83 CDN VDD VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net083 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=0.62u l=0.18u
MI233 net0147 net083 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.78u l=0.18u
.ends
.subckt SEDFCND2BWP7T E SE CP SI D CDN Q QN VDD VSS 
MI239 net080 net090 net079 VSS n w=0.52u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net92 d1 VSS VSS n w=0.42u l=0.18u
MI119 net95 CDN net92 VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net090 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.52u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI183-M_u4 XI183-net6 CDN VSS VSS n w=0.97u l=0.18u
MI183-M_u3 d2 net084 XI183-net6 VSS n w=0.97u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI189_0-M_u2 QN net090 VSS VSS n w=1u l=0.18u
MI189_1-M_u2 QN net090 VSS VSS n w=1u l=0.18u
MI175_0-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI175_1-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI177-M_u2 net090 d2 VSS VSS n w=0.97u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI183-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI183-M_u1 d2 net084 VDD VDD p w=1.23u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI189_0-M_u3 QN net090 VDD VDD p w=1.3u l=0.18u
MI189_1-M_u3 QN net090 VDD VDD p w=1.3u l=0.18u
MI175_0-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI175_1-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI177-M_u3 net090 d2 VDD VDD p w=0.97u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.42u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0151 VDD p w=0.42u l=0.18u
MI101 net83 CDN VDD VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net090 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=0.62u l=0.18u
MI233 net0147 net090 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0151 VDD p w=0.87u l=0.18u
MI231 net0151 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.78u l=0.18u
.ends
.subckt SEDFCNQD0BWP7T E SE CP SI D CDN Q VDD VSS 
MI239 net080 net083 net079 VSS n w=0.52u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net92 d1 VSS VSS n w=0.42u l=0.18u
MI119 net95 CDN net92 VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net083 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.52u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI183-M_u4 XI183-net6 CDN VSS VSS n w=1u l=0.18u
MI183-M_u3 d2 net084 XI183-net6 VSS n w=1u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI175-M_u2 Q d2 VSS VSS n w=0.5u l=0.18u
MI177-M_u2 net083 d2 VSS VSS n w=0.42u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI183-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI183-M_u1 d2 net084 VDD VDD p w=1.035u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI175-M_u3 Q d2 VDD VDD p w=0.685u l=0.18u
MI177-M_u3 net083 d2 VDD VDD p w=0.42u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.42u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI101 net83 CDN VDD VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net083 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=0.62u l=0.18u
MI233 net0147 net083 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.78u l=0.18u
.ends
.subckt SEDFCNQD1BWP7T E SE CP SI D CDN Q VDD VSS 
MI239 net080 net083 net079 VSS n w=0.52u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net92 d1 VSS VSS n w=0.42u l=0.18u
MI119 net95 CDN net92 VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net083 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.52u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI183-M_u4 XI183-net6 CDN VSS VSS n w=1u l=0.18u
MI183-M_u3 d2 net084 XI183-net6 VSS n w=1u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI175-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI177-M_u2 net083 d2 VSS VSS n w=0.42u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI183-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI183-M_u1 d2 net084 VDD VDD p w=1.035u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI175-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI177-M_u3 net083 d2 VDD VDD p w=0.42u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.42u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI101 net83 CDN VDD VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net083 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=0.62u l=0.18u
MI233 net0147 net083 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.78u l=0.18u
.ends
.subckt SEDFCNQD2BWP7T E SE CP SI D CDN Q VDD VSS 
MI239 net080 net090 net079 VSS n w=0.52u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net92 d1 VSS VSS n w=0.42u l=0.18u
MI119 net95 CDN net92 VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net090 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.52u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI183-M_u4 XI183-net6 CDN VSS VSS n w=1u l=0.18u
MI183-M_u3 d2 net084 XI183-net6 VSS n w=1u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI175_0-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI175_1-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI177-M_u2 net090 d2 VSS VSS n w=0.42u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI183-M_u2 d2 CDN VDD VDD p w=0.42u l=0.18u
MI183-M_u1 d2 net084 VDD VDD p w=1.035u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.62u l=0.18u
MI175_0-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI175_1-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI177-M_u3 net090 d2 VDD VDD p w=0.42u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.42u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0151 VDD p w=0.42u l=0.18u
MI101 net83 CDN VDD VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net090 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=0.62u l=0.18u
MI233 net0147 net090 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0151 VDD p w=0.87u l=0.18u
MI231 net0151 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.78u l=0.18u
.ends
.subckt SEDFD0BWP7T E SE CP SI D Q QN VDD VSS 
MI239 net080 net087 net079 VSS n w=0.42u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net95 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net087 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.42u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI189-M_u2 QN net087 VSS VSS n w=0.5u l=0.18u
MI175-M_u2 Q d2 VSS VSS n w=0.5u l=0.18u
MI177-M_u2 net087 d2 VSS VSS n w=0.42u l=0.18u
MI190-M_u2 d2 net084 VSS VSS n w=0.5u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.84u l=0.18u
MI189-M_u3 QN net087 VDD VDD p w=0.685u l=0.18u
MI175-M_u3 Q d2 VDD VDD p w=0.685u l=0.18u
MI177-M_u3 net087 d2 VDD VDD p w=0.685u l=0.18u
MI190-M_u3 d2 net084 VDD VDD p w=0.685u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net087 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=1.34u l=0.18u
MI233 net0147 net087 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.62u l=0.18u
.ends
.subckt SEDFD1BWP7T E SE CP SI D Q QN VDD VSS 
MI239 net080 net087 net079 VSS n w=0.42u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net95 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net087 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.42u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI189-M_u2 QN net087 VSS VSS n w=0.94u l=0.18u
MI175-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI177-M_u2 net087 d2 VSS VSS n w=0.42u l=0.18u
MI190-M_u2 d2 net084 VSS VSS n w=1u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.84u l=0.18u
MI189-M_u3 QN net087 VDD VDD p w=1.37u l=0.18u
MI175-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI177-M_u3 net087 d2 VDD VDD p w=0.685u l=0.18u
MI190-M_u3 d2 net084 VDD VDD p w=1.37u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net087 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=1.34u l=0.18u
MI233 net0147 net087 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.62u l=0.18u
.ends
.subckt SEDFD2BWP7T E SE CP SI D Q QN VDD VSS 
MI239 net080 net087 net079 VSS n w=0.42u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net95 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net087 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.42u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI189_0-M_u2 QN net087 VSS VSS n w=1u l=0.18u
MI189_1-M_u2 QN net087 VSS VSS n w=1u l=0.18u
MI175_0-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI175_1-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI177-M_u2 net087 d2 VSS VSS n w=1u l=0.18u
MI190-M_u2 d2 net084 VSS VSS n w=1u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.84u l=0.18u
MI189_0-M_u3 QN net087 VDD VDD p w=1.3u l=0.18u
MI189_1-M_u3 QN net087 VDD VDD p w=1.3u l=0.18u
MI175_0-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI175_1-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI177-M_u3 net087 d2 VDD VDD p w=1.37u l=0.18u
MI190-M_u3 d2 net084 VDD VDD p w=1.23u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net087 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=1.34u l=0.18u
MI233 net0147 net087 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.62u l=0.18u
.ends
.subckt SEDFKCND0BWP7T SI D E SE CP CN Q QN VDD VSS 
MI188 net170 net171 net169 VSS n w=0.42u l=0.18u
MI187 net112 net136 net170 VSS n w=0.42u l=0.18u
MI189 net169 CN net176 VSS n w=0.57u l=0.18u
MI190 net151 net165 VSS VSS n w=0.42u l=0.18u
MI197 net165 INCP net142 VSS n w=0.91u l=0.18u
MI192 net154 D net169 VSS n w=0.57u l=0.18u
MI191 net171 INCPB net142 VSS n w=0.42u l=0.18u
MI194 d0 INCP net151 VSS n w=0.42u l=0.18u
MI196 net112 SE net145 VSS n w=0.42u l=0.18u
MI193 net112 E net154 VSS n w=0.94u l=0.18u
MI185 net145 SI VSS VSS n w=0.42u l=0.18u
MI186 net176 net138 VSS VSS n w=0.57u l=0.18u
MI195 d0 INCPB net112 VSS n w=0.91u l=0.18u
MI177-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI184-M_u2 net124 net142 VSS VSS n w=0.5u l=0.18u
MI181-M_u2 net171 net124 VSS VSS n w=0.42u l=0.18u
MI178-M_u2 net138 SE VSS VSS n w=0.5u l=0.18u
MI183-M_u2 net165 d0 VSS VSS n w=0.54u l=0.18u
MI180-M_u2 Q net124 VSS VSS n w=0.5u l=0.18u
MI179-M_u2 net136 E VSS VSS n w=0.5u l=0.18u
MI218-M_u2 QN net171 VSS VSS n w=0.5u l=0.18u
MI182-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI177-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI184-M_u3 net124 net142 VDD VDD p w=0.685u l=0.18u
MI181-M_u3 net171 net124 VDD VDD p w=0.685u l=0.18u
MI178-M_u3 net138 SE VDD VDD p w=0.65u l=0.18u
MI183-M_u3 net165 d0 VDD VDD p w=0.84u l=0.18u
MI180-M_u3 Q net124 VDD VDD p w=0.685u l=0.18u
MI179-M_u3 net136 E VDD VDD p w=0.685u l=0.18u
MI218-M_u3 QN net171 VDD VDD p w=0.685u l=0.18u
MI182-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI168 net96 SE VDD VDD p w=0.75u l=0.18u
MI166 net165 INCPB net142 VDD p w=1.34u l=0.18u
MI162 net120 net165 VDD VDD p w=0.42u l=0.18u
MI176 net112 CN net96 VDD p w=0.42u l=0.18u
MI172 net112 net136 net91 VDD p w=0.685u l=0.18u
MI171 net100 SI VDD VDD p w=0.42u l=0.18u
MI170 net112 net171 net105 VDD p w=0.42u l=0.18u
MI175 d0 INCP net112 VDD p w=0.62u l=0.18u
MI169 net171 INCP net142 VDD p w=0.42u l=0.18u
MI167 net112 net138 net100 VDD p w=0.42u l=0.18u
MI173 net105 E net96 VDD p w=0.42u l=0.18u
MI174 net91 D net96 VDD p w=0.75u l=0.18u
MI165 d0 INCPB net120 VDD p w=0.42u l=0.18u
.ends
.subckt SEDFKCND1BWP7T SI D E SE CP CN Q QN VDD VSS 
MI188 net170 net171 net169 VSS n w=0.42u l=0.18u
MI187 net112 net136 net170 VSS n w=0.42u l=0.18u
MI189 net169 CN net176 VSS n w=0.57u l=0.18u
MI190 net151 net165 VSS VSS n w=0.42u l=0.18u
MI197 net165 INCP net142 VSS n w=0.91u l=0.18u
MI192 net154 D net169 VSS n w=0.57u l=0.18u
MI191 net171 INCPB net142 VSS n w=0.42u l=0.18u
MI194 d0 INCP net151 VSS n w=0.42u l=0.18u
MI196 net112 SE net145 VSS n w=0.42u l=0.18u
MI193 net112 E net154 VSS n w=0.94u l=0.18u
MI185 net145 SI VSS VSS n w=0.42u l=0.18u
MI186 net176 net138 VSS VSS n w=0.57u l=0.18u
MI195 d0 INCPB net112 VSS n w=0.91u l=0.18u
MI177-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI184-M_u2 net124 net142 VSS VSS n w=1u l=0.18u
MI181-M_u2 net171 net124 VSS VSS n w=0.42u l=0.18u
MI178-M_u2 net138 SE VSS VSS n w=0.5u l=0.18u
MI183-M_u2 net165 d0 VSS VSS n w=0.54u l=0.18u
MI180-M_u2 Q net124 VSS VSS n w=1u l=0.18u
MI179-M_u2 net136 E VSS VSS n w=0.5u l=0.18u
MI218-M_u2 QN net171 VSS VSS n w=0.94u l=0.18u
MI182-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI177-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI184-M_u3 net124 net142 VDD VDD p w=1.37u l=0.18u
MI181-M_u3 net171 net124 VDD VDD p w=0.685u l=0.18u
MI178-M_u3 net138 SE VDD VDD p w=0.65u l=0.18u
MI183-M_u3 net165 d0 VDD VDD p w=0.84u l=0.18u
MI180-M_u3 Q net124 VDD VDD p w=1.37u l=0.18u
MI179-M_u3 net136 E VDD VDD p w=0.685u l=0.18u
MI218-M_u3 QN net171 VDD VDD p w=1.37u l=0.18u
MI182-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI168 net96 SE VDD VDD p w=0.75u l=0.18u
MI166 net165 INCPB net142 VDD p w=1.34u l=0.18u
MI162 net120 net165 VDD VDD p w=0.42u l=0.18u
MI176 net112 CN net96 VDD p w=0.42u l=0.18u
MI172 net112 net136 net91 VDD p w=0.685u l=0.18u
MI171 net100 SI VDD VDD p w=0.42u l=0.18u
MI170 net112 net171 net105 VDD p w=0.42u l=0.18u
MI175 d0 INCP net112 VDD p w=0.62u l=0.18u
MI169 net171 INCP net142 VDD p w=0.42u l=0.18u
MI167 net112 net138 net100 VDD p w=0.42u l=0.18u
MI173 net105 E net96 VDD p w=0.42u l=0.18u
MI174 net91 D net96 VDD p w=0.75u l=0.18u
MI165 d0 INCPB net120 VDD p w=0.42u l=0.18u
.ends
.subckt SEDFKCND2BWP7T SI D E SE CP CN Q QN VDD VSS 
MI188 net170 net171 net169 VSS n w=0.42u l=0.18u
MI187 net112 net136 net170 VSS n w=0.42u l=0.18u
MI189 net169 CN net176 VSS n w=0.57u l=0.18u
MI190 net151 net165 VSS VSS n w=0.42u l=0.18u
MI197 net165 INCP net142 VSS n w=0.91u l=0.18u
MI192 net154 D net169 VSS n w=0.57u l=0.18u
MI191 net171 INCPB net142 VSS n w=0.42u l=0.18u
MI194 d0 INCP net151 VSS n w=0.42u l=0.18u
MI196 net112 SE net145 VSS n w=0.42u l=0.18u
MI193 net112 E net154 VSS n w=0.94u l=0.18u
MI185 net145 SI VSS VSS n w=0.42u l=0.18u
MI186 net176 net138 VSS VSS n w=0.57u l=0.18u
MI195 d0 INCPB net112 VSS n w=0.91u l=0.18u
MI177-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI184-M_u2 net124 net142 VSS VSS n w=1u l=0.18u
MI181-M_u2 net171 net124 VSS VSS n w=1u l=0.18u
MI178-M_u2 net138 SE VSS VSS n w=0.5u l=0.18u
MI183-M_u2 net165 d0 VSS VSS n w=0.54u l=0.18u
MI180_0-M_u2 Q net124 VSS VSS n w=1u l=0.18u
MI180_1-M_u2 Q net124 VSS VSS n w=1u l=0.18u
MI179-M_u2 net136 E VSS VSS n w=0.5u l=0.18u
MI218-M_u2 QN net171 VSS VSS n w=2u l=0.18u
MI182-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI177-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI184-M_u3 net124 net142 VDD VDD p w=1.235u l=0.18u
MI181-M_u3 net171 net124 VDD VDD p w=1.37u l=0.18u
MI178-M_u3 net138 SE VDD VDD p w=0.65u l=0.18u
MI183-M_u3 net165 d0 VDD VDD p w=0.84u l=0.18u
MI180_0-M_u3 Q net124 VDD VDD p w=1.37u l=0.18u
MI180_1-M_u3 Q net124 VDD VDD p w=1.37u l=0.18u
MI179-M_u3 net136 E VDD VDD p w=0.685u l=0.18u
MI218-M_u3 QN net171 VDD VDD p w=2.605u l=0.18u
MI182-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI168 net96 SE VDD VDD p w=0.75u l=0.18u
MI166 net165 INCPB net142 VDD p w=1.34u l=0.18u
MI162 net120 net165 VDD VDD p w=0.42u l=0.18u
MI176 net112 CN net96 VDD p w=0.42u l=0.18u
MI172 net112 net136 net91 VDD p w=0.685u l=0.18u
MI171 net100 SI VDD VDD p w=0.42u l=0.18u
MI170 net112 net171 net105 VDD p w=0.42u l=0.18u
MI175 d0 INCP net112 VDD p w=0.62u l=0.18u
MI169 net171 INCP net142 VDD p w=0.42u l=0.18u
MI167 net112 net138 net100 VDD p w=0.42u l=0.18u
MI173 net105 E net96 VDD p w=0.42u l=0.18u
MI174 net91 D net96 VDD p w=0.75u l=0.18u
MI165 d0 INCPB net120 VDD p w=0.42u l=0.18u
.ends
.subckt SEDFKCNQD0BWP7T SI D E SE CP CN Q VDD VSS 
MI188 net170 net171 net169 VSS n w=0.42u l=0.18u
MI187 net112 net136 net170 VSS n w=0.42u l=0.18u
MI189 net169 CN net176 VSS n w=0.57u l=0.18u
MI190 net151 net165 VSS VSS n w=0.42u l=0.18u
MI197 net165 INCP net142 VSS n w=0.91u l=0.18u
MI192 net154 D net169 VSS n w=0.57u l=0.18u
MI191 net171 INCPB net142 VSS n w=0.42u l=0.18u
MI194 d0 INCP net151 VSS n w=0.42u l=0.18u
MI196 net112 SE net145 VSS n w=0.42u l=0.18u
MI193 net112 E net154 VSS n w=0.94u l=0.18u
MI185 net145 SI VSS VSS n w=0.42u l=0.18u
MI186 net176 net138 VSS VSS n w=0.57u l=0.18u
MI195 d0 INCPB net112 VSS n w=0.91u l=0.18u
MI177-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI184-M_u2 net124 net142 VSS VSS n w=0.5u l=0.18u
MI181-M_u2 net171 net124 VSS VSS n w=0.42u l=0.18u
MI178-M_u2 net138 SE VSS VSS n w=0.5u l=0.18u
MI183-M_u2 net165 d0 VSS VSS n w=0.54u l=0.18u
MI180-M_u2 Q net124 VSS VSS n w=0.5u l=0.18u
MI179-M_u2 net136 E VSS VSS n w=0.5u l=0.18u
MI182-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI177-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI184-M_u3 net124 net142 VDD VDD p w=0.685u l=0.18u
MI181-M_u3 net171 net124 VDD VDD p w=0.42u l=0.18u
MI178-M_u3 net138 SE VDD VDD p w=0.65u l=0.18u
MI183-M_u3 net165 d0 VDD VDD p w=0.84u l=0.18u
MI180-M_u3 Q net124 VDD VDD p w=0.685u l=0.18u
MI179-M_u3 net136 E VDD VDD p w=0.685u l=0.18u
MI182-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI168 net96 SE VDD VDD p w=0.75u l=0.18u
MI166 net165 INCPB net142 VDD p w=1.34u l=0.18u
MI162 net120 net165 VDD VDD p w=0.42u l=0.18u
MI176 net112 CN net96 VDD p w=0.42u l=0.18u
MI172 net112 net136 net91 VDD p w=0.685u l=0.18u
MI171 net100 SI VDD VDD p w=0.42u l=0.18u
MI170 net112 net171 net105 VDD p w=0.42u l=0.18u
MI175 d0 INCP net112 VDD p w=0.62u l=0.18u
MI169 net171 INCP net142 VDD p w=0.42u l=0.18u
MI167 net112 net138 net100 VDD p w=0.42u l=0.18u
MI173 net105 E net96 VDD p w=0.42u l=0.18u
MI174 net91 D net96 VDD p w=0.75u l=0.18u
MI165 d0 INCPB net120 VDD p w=0.42u l=0.18u
.ends
.subckt SEDFKCNQD1BWP7T SI D E SE CP CN Q VDD VSS 
MI188 net170 net171 net169 VSS n w=0.42u l=0.18u
MI187 net112 net136 net170 VSS n w=0.42u l=0.18u
MI189 net169 CN net176 VSS n w=0.57u l=0.18u
MI190 net151 net165 VSS VSS n w=0.42u l=0.18u
MI197 net165 INCP net142 VSS n w=0.91u l=0.18u
MI192 net154 D net169 VSS n w=0.57u l=0.18u
MI191 net171 INCPB net142 VSS n w=0.42u l=0.18u
MI194 d0 INCP net151 VSS n w=0.42u l=0.18u
MI196 net112 SE net145 VSS n w=0.42u l=0.18u
MI193 net112 E net154 VSS n w=0.94u l=0.18u
MI185 net145 SI VSS VSS n w=0.42u l=0.18u
MI186 net176 net138 VSS VSS n w=0.57u l=0.18u
MI195 d0 INCPB net112 VSS n w=0.91u l=0.18u
MI177-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI184-M_u2 net124 net142 VSS VSS n w=1u l=0.18u
MI181-M_u2 net171 net124 VSS VSS n w=0.42u l=0.18u
MI178-M_u2 net138 SE VSS VSS n w=0.5u l=0.18u
MI183-M_u2 net165 d0 VSS VSS n w=0.54u l=0.18u
MI180-M_u2 Q net124 VSS VSS n w=1u l=0.18u
MI179-M_u2 net136 E VSS VSS n w=0.5u l=0.18u
MI182-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI177-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI184-M_u3 net124 net142 VDD VDD p w=1.37u l=0.18u
MI181-M_u3 net171 net124 VDD VDD p w=0.42u l=0.18u
MI178-M_u3 net138 SE VDD VDD p w=0.65u l=0.18u
MI183-M_u3 net165 d0 VDD VDD p w=0.84u l=0.18u
MI180-M_u3 Q net124 VDD VDD p w=1.37u l=0.18u
MI179-M_u3 net136 E VDD VDD p w=0.685u l=0.18u
MI182-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI168 net96 SE VDD VDD p w=0.75u l=0.18u
MI166 net165 INCPB net142 VDD p w=1.34u l=0.18u
MI162 net120 net165 VDD VDD p w=0.42u l=0.18u
MI176 net112 CN net96 VDD p w=0.42u l=0.18u
MI172 net112 net136 net91 VDD p w=0.685u l=0.18u
MI171 net100 SI VDD VDD p w=0.42u l=0.18u
MI170 net112 net171 net105 VDD p w=0.42u l=0.18u
MI175 d0 INCP net112 VDD p w=0.62u l=0.18u
MI169 net171 INCP net142 VDD p w=0.42u l=0.18u
MI167 net112 net138 net100 VDD p w=0.42u l=0.18u
MI173 net105 E net96 VDD p w=0.42u l=0.18u
MI174 net91 D net96 VDD p w=0.75u l=0.18u
MI165 d0 INCPB net120 VDD p w=0.42u l=0.18u
.ends
.subckt SEDFKCNQD2BWP7T SI D E SE CP CN Q VDD VSS 
MI188 net170 net171 net169 VSS n w=0.42u l=0.18u
MI187 net112 net136 net170 VSS n w=0.42u l=0.18u
MI189 net169 CN net176 VSS n w=0.57u l=0.18u
MI190 net151 net165 VSS VSS n w=0.42u l=0.18u
MI197 net165 INCP net142 VSS n w=0.91u l=0.18u
MI192 net154 D net169 VSS n w=0.57u l=0.18u
MI191 net171 INCPB net142 VSS n w=0.42u l=0.18u
MI194 d0 INCP net151 VSS n w=0.42u l=0.18u
MI196 net112 SE net145 VSS n w=0.42u l=0.18u
MI193 net112 E net154 VSS n w=0.94u l=0.18u
MI185 net145 SI VSS VSS n w=0.42u l=0.18u
MI186 net176 net138 VSS VSS n w=0.57u l=0.18u
MI195 d0 INCPB net112 VSS n w=0.91u l=0.18u
MI177-M_u2 INCP INCPB VSS VSS n w=0.5u l=0.18u
MI184-M_u2 net124 net142 VSS VSS n w=1u l=0.18u
MI181-M_u2 net171 net124 VSS VSS n w=0.42u l=0.18u
MI178-M_u2 net138 SE VSS VSS n w=0.5u l=0.18u
MI183-M_u2 net165 d0 VSS VSS n w=0.54u l=0.18u
MI180_0-M_u2 Q net124 VSS VSS n w=1u l=0.18u
MI180_1-M_u2 Q net124 VSS VSS n w=1u l=0.18u
MI179-M_u2 net136 E VSS VSS n w=0.5u l=0.18u
MI182-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI177-M_u3 INCP INCPB VDD VDD p w=0.685u l=0.18u
MI184-M_u3 net124 net142 VDD VDD p w=1.37u l=0.18u
MI181-M_u3 net171 net124 VDD VDD p w=0.42u l=0.18u
MI178-M_u3 net138 SE VDD VDD p w=0.65u l=0.18u
MI183-M_u3 net165 d0 VDD VDD p w=0.84u l=0.18u
MI180_0-M_u3 Q net124 VDD VDD p w=1.37u l=0.18u
MI180_1-M_u3 Q net124 VDD VDD p w=1.37u l=0.18u
MI179-M_u3 net136 E VDD VDD p w=0.685u l=0.18u
MI182-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI168 net96 SE VDD VDD p w=0.75u l=0.18u
MI166 net165 INCPB net142 VDD p w=1.34u l=0.18u
MI162 net120 net165 VDD VDD p w=0.42u l=0.18u
MI176 net112 CN net96 VDD p w=0.42u l=0.18u
MI172 net112 net136 net91 VDD p w=0.685u l=0.18u
MI171 net100 SI VDD VDD p w=0.42u l=0.18u
MI170 net112 net171 net105 VDD p w=0.42u l=0.18u
MI175 d0 INCP net112 VDD p w=0.62u l=0.18u
MI169 net171 INCP net142 VDD p w=0.42u l=0.18u
MI167 net112 net138 net100 VDD p w=0.42u l=0.18u
MI173 net105 E net96 VDD p w=0.42u l=0.18u
MI174 net91 D net96 VDD p w=0.75u l=0.18u
MI165 d0 INCPB net120 VDD p w=0.42u l=0.18u
.ends
.subckt SEDFQD0BWP7T E SE CP SI D Q VDD VSS 
MI239 net080 net090 net079 VSS n w=0.42u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net95 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net090 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.42u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI175-M_u2 Q d2 VSS VSS n w=0.5u l=0.18u
MI177-M_u2 net090 d2 VSS VSS n w=0.42u l=0.18u
MI190-M_u2 d2 net084 VSS VSS n w=0.5u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.84u l=0.18u
MI175-M_u3 Q d2 VDD VDD p w=0.685u l=0.18u
MI177-M_u3 net090 d2 VDD VDD p w=0.42u l=0.18u
MI190-M_u3 d2 net084 VDD VDD p w=0.685u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net090 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=1.34u l=0.18u
MI233 net0147 net090 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.62u l=0.18u
.ends
.subckt SEDFQD1BWP7T E SE CP SI D Q VDD VSS 
MI239 net080 net090 net079 VSS n w=0.42u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net95 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net090 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.42u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI175-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI177-M_u2 net090 d2 VSS VSS n w=0.42u l=0.18u
MI190-M_u2 d2 net084 VSS VSS n w=1u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.84u l=0.18u
MI175-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI177-M_u3 net090 d2 VDD VDD p w=0.42u l=0.18u
MI190-M_u3 d2 net084 VDD VDD p w=1.37u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net090 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=1.34u l=0.18u
MI233 net0147 net090 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.62u l=0.18u
.ends
.subckt SEDFQD2BWP7T E SE CP SI D Q VDD VSS 
MI239 net080 net090 net079 VSS n w=0.42u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net95 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net090 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.42u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI175_0-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI175_1-M_u2 Q d2 VSS VSS n w=1u l=0.18u
MI177-M_u2 net090 d2 VSS VSS n w=0.42u l=0.18u
MI190-M_u2 d2 net084 VSS VSS n w=1u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.84u l=0.18u
MI175_0-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI175_1-M_u3 Q d2 VDD VDD p w=1.37u l=0.18u
MI177-M_u3 net090 d2 VDD VDD p w=0.42u l=0.18u
MI190-M_u3 d2 net084 VDD VDD p w=1.37u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net090 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=1.34u l=0.18u
MI233 net0147 net090 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.62u l=0.18u
.ends
.subckt SEDFQND0BWP7T E SE CP SI D QN VDD VSS 
MI239 net080 net087 net079 VSS n w=0.42u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net95 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net087 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.42u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI189-M_u2 QN net087 VSS VSS n w=0.5u l=0.18u
MI177-M_u2 net087 net077 VSS VSS n w=0.42u l=0.18u
MI190-M_u2 net077 net084 VSS VSS n w=0.5u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.84u l=0.18u
MI189-M_u3 QN net087 VDD VDD p w=0.685u l=0.18u
MI177-M_u3 net087 net077 VDD VDD p w=0.685u l=0.18u
MI190-M_u3 net077 net084 VDD VDD p w=0.685u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net087 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=1.34u l=0.18u
MI233 net0147 net087 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.62u l=0.18u
.ends
.subckt SEDFQND1BWP7T E SE CP SI D QN VDD VSS 
MI239 net080 net087 net079 VSS n w=0.42u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net95 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net087 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.42u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI189-M_u2 QN net087 VSS VSS n w=1u l=0.18u
MI177-M_u2 net087 net077 VSS VSS n w=0.42u l=0.18u
MI190-M_u2 net077 net084 VSS VSS n w=0.665u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.84u l=0.18u
MI189-M_u3 QN net087 VDD VDD p w=1.37u l=0.18u
MI177-M_u3 net087 net077 VDD VDD p w=1.37u l=0.18u
MI190-M_u3 net077 net084 VDD VDD p w=1.37u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net087 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=1.34u l=0.18u
MI233 net0147 net087 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.62u l=0.18u
.ends
.subckt SEDFQND2BWP7T E SE CP SI D QN VDD VSS 
MI239 net080 net085 net079 VSS n w=0.42u l=0.18u
MI174 d1 INCP net084 VSS n w=0.91u l=0.18u
MI118 net95 d1 VSS VSS n w=0.42u l=0.18u
MI120 d0 INCP net95 VSS n w=0.42u l=0.18u
MI173 net085 INCPB net084 VSS n w=0.42u l=0.18u
MI237 net0147 SE net0113 VSS n w=0.42u l=0.18u
MI163 net074 D net079 VSS n w=0.64u l=0.18u
MI238 net0147 net0128 net080 VSS n w=0.42u l=0.18u
MI160 net0147 E net074 VSS n w=0.64u l=0.18u
MI164 d0 INCPB net0147 VSS n w=0.42u l=0.18u
MI236 net0113 SI VSS VSS n w=0.42u l=0.18u
MI240 net079 net0126 VSS VSS n w=0.57u l=0.18u
MI188-M_u2 d1 d0 VSS VSS n w=0.54u l=0.18u
MI189_0-M_u2 QN net085 VSS VSS n w=1u l=0.18u
MI189_1-M_u2 QN net085 VSS VSS n w=1u l=0.18u
MI177-M_u2 net085 net077 VSS VSS n w=0.42u l=0.18u
MI190-M_u2 net077 net084 VSS VSS n w=0.66u l=0.18u
MI229-M_u2 net0128 E VSS VSS n w=0.5u l=0.18u
MI230-M_u2 net0126 SE VSS VSS n w=0.5u l=0.18u
MU85-M_u2 INCP INCPB VSS VSS n w=0.9u l=0.18u
MI181-M_u2 INCPB CP VSS VSS n w=0.5u l=0.18u
MI188-M_u3 d1 d0 VDD VDD p w=0.84u l=0.18u
MI189_0-M_u3 QN net085 VDD VDD p w=1.37u l=0.18u
MI189_1-M_u3 QN net085 VDD VDD p w=1.37u l=0.18u
MI177-M_u3 net085 net077 VDD VDD p w=1.37u l=0.18u
MI190-M_u3 net077 net084 VDD VDD p w=1.37u l=0.18u
MI229-M_u3 net0128 E VDD VDD p w=0.685u l=0.18u
MI230-M_u3 net0126 SE VDD VDD p w=0.65u l=0.18u
MU85-M_u3 INCP INCPB VDD VDD p w=0.6u l=0.18u
MI181-M_u3 INCPB CP VDD VDD p w=0.685u l=0.18u
MI150 net0147 net0128 net0134 VDD p w=0.87u l=0.18u
MI232 net0158 E net0137 VDD p w=0.42u l=0.18u
MI102 net83 d1 VDD VDD p w=0.42u l=0.18u
MI103 d0 INCPB net83 VDD p w=0.42u l=0.18u
MI234 net0147 net0126 net0165 VDD p w=0.42u l=0.18u
MI178 net085 INCP net084 VDD p w=0.42u l=0.18u
MI179 d1 INCPB net084 VDD p w=1.34u l=0.18u
MI233 net0147 net085 net0158 VDD p w=0.42u l=0.18u
MI151 net0134 D net0137 VDD p w=0.87u l=0.18u
MI231 net0137 SE VDD VDD p w=0.75u l=0.18u
MI235 net0165 SI VDD VDD p w=0.42u l=0.18u
MI153 d0 INCP net0147 VDD p w=0.62u l=0.18u
.ends
.subckt TIEHBWP7T Z VDD VSS 
M_u2 net6 net6 VSS VSS n w=1u l=0.18u
M_u1 Z net6 VDD VDD p w=1.37u l=0.18u
.ends
.subckt TIELBWP7T ZN VDD VSS 
M_u2 ZN net6 VSS VSS n w=1u l=0.18u
M_u1 net6 net6 VDD VDD p w=1.37u l=0.18u
.ends
.subckt XNR2D0BWP7T A1 A2 ZN VDD VSS 
MI0-M_u2 net4 A1 net14 VSS n w=0.5u l=0.18u
M_u7-M_u2 net6 net10 net14 VSS n w=0.5u l=0.18u
M_u2-M_u2 net4 A2 VSS VSS n w=0.5u l=0.18u
M_u5-M_u2 net6 net4 VSS VSS n w=0.5u l=0.18u
M_u4-M_u2 ZN net14 VSS VSS n w=0.5u l=0.18u
M_u8-M_u2 net10 A1 VSS VSS n w=0.5u l=0.18u
MI0-M_u3 net4 net10 net14 VDD p w=0.685u l=0.18u
M_u7-M_u3 net6 A1 net14 VDD p w=0.685u l=0.18u
M_u2-M_u3 net4 A2 VDD VDD p w=0.685u l=0.18u
M_u5-M_u3 net6 net4 VDD VDD p w=0.685u l=0.18u
M_u4-M_u3 ZN net14 VDD VDD p w=0.685u l=0.18u
M_u8-M_u3 net10 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XNR2D1BWP7T A1 A2 ZN VDD VSS 
MI9 net025 net4 VSS VSS n w=0.5u l=0.18u
MI10 net14 net10 net025 VSS n w=0.5u l=0.18u
M_u6-M_u2 net4 A1 net14 VSS n w=0.5u l=0.18u
M_u2-M_u2 net4 A2 VSS VSS n w=1u l=0.18u
M_u4-M_u2 ZN net14 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net10 A1 VSS VSS n w=0.5u l=0.18u
MI6 net016 net4 VDD VDD p w=0.685u l=0.18u
MI7 net14 A1 net016 VDD p w=0.685u l=0.18u
M_u6-M_u3 net4 net10 net14 VDD p w=0.685u l=0.18u
M_u2-M_u3 net4 A2 VDD VDD p w=1.37u l=0.18u
M_u4-M_u3 ZN net14 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net10 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XNR2D2BWP7T A1 A2 ZN VDD VSS 
M_u6-M_u2 net4 A1 net14 VSS n w=0.5u l=0.18u
M_u7-M_u2 net6 net10 net14 VSS n w=0.5u l=0.18u
M_u2-M_u2 net4 A2 VSS VSS n w=1u l=0.18u
M_u5-M_u2 net6 net4 VSS VSS n w=1u l=0.18u
M_u4_0-M_u2 ZN net14 VSS VSS n w=1u l=0.18u
M_u4_1-M_u2 ZN net14 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net10 A1 VSS VSS n w=0.5u l=0.18u
M_u6-M_u3 net4 net10 net14 VDD p w=0.685u l=0.18u
M_u7-M_u3 net6 A1 net14 VDD p w=0.685u l=0.18u
M_u2-M_u3 net4 A2 VDD VDD p w=1.37u l=0.18u
M_u5-M_u3 net6 net4 VDD VDD p w=1.37u l=0.18u
M_u4_0-M_u3 ZN net14 VDD VDD p w=1.37u l=0.18u
M_u4_1-M_u3 ZN net14 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net10 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XNR3D0BWP7T A1 A2 A3 ZN VDD VSS 
MI3-M_u2 net11 A2 net17 VSS n w=0.5u l=0.18u
MU11-M_u2 net5 net17 net21 VSS n w=0.5u l=0.18u
MI5-M_u2 net5 A3 VSS VSS n w=0.5u l=0.18u
MU22-M_u2 ZN net21 VSS VSS n w=0.5u l=0.18u
M_u8-M_u2 net16 A2 VSS VSS n w=0.5u l=0.18u
MI4-M_u2 net11 A1 VSS VSS n w=0.705u l=0.18u
MI6-M_u2 net13 net17 VSS VSS n w=0.5u l=0.18u
MI2-MU3 net17 net16 XI2-net16 VSS n w=0.5u l=0.18u
MI2-MU4 XI2-net16 net11 VSS VSS n w=0.5u l=0.18u
MU21-MU3 net21 net13 XU21-net16 VSS n w=0.5u l=0.18u
MU21-MU4 XU21-net16 net5 VSS VSS n w=0.5u l=0.18u
MI3-M_u3 net11 net16 net17 VDD p w=0.685u l=0.18u
MU11-M_u3 net5 net13 net21 VDD p w=0.685u l=0.18u
MI5-M_u3 net5 A3 VDD VDD p w=0.685u l=0.18u
MU22-M_u3 ZN net21 VDD VDD p w=0.685u l=0.18u
M_u8-M_u3 net16 A2 VDD VDD p w=0.685u l=0.18u
MI4-M_u3 net11 A1 VDD VDD p w=0.685u l=0.18u
MI6-M_u3 net13 net17 VDD VDD p w=0.685u l=0.18u
MI2-MU2 net17 A2 XI2-net6 VDD p w=0.685u l=0.18u
MI2-MU1 XI2-net6 net11 VDD VDD p w=0.685u l=0.18u
MU21-MU2 net21 net17 XU21-net6 VDD p w=0.685u l=0.18u
MU21-MU1 XU21-net6 net5 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XNR3D1BWP7T A1 A2 A3 ZN VDD VSS 
M_u6-M_u2 net11 A2 net17 VSS n w=0.5u l=0.18u
MU11-M_u2 net5 net17 net21 VSS n w=0.5u l=0.18u
MI1-M_u2 net5 A3 VSS VSS n w=1u l=0.18u
MU22-M_u2 ZN net21 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net16 A2 VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net11 A1 VSS VSS n w=1u l=0.18u
MU12-M_u2 net13 net17 VSS VSS n w=0.5u l=0.18u
MI0-MU3 net17 net16 XI0-net16 VSS n w=0.5u l=0.18u
MI0-MU4 XI0-net16 net11 VSS VSS n w=0.5u l=0.18u
MU21-MU3 net21 net13 XU21-net16 VSS n w=0.5u l=0.18u
MU21-MU4 XU21-net16 net5 VSS VSS n w=0.5u l=0.18u
M_u6-M_u3 net11 net16 net17 VDD p w=0.68u l=0.18u
MU11-M_u3 net5 net13 net21 VDD p w=0.685u l=0.18u
MI1-M_u3 net5 A3 VDD VDD p w=1.37u l=0.18u
MU22-M_u3 ZN net21 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net16 A2 VDD VDD p w=0.685u l=0.18u
M_u2-M_u3 net11 A1 VDD VDD p w=1.37u l=0.18u
MU12-M_u3 net13 net17 VDD VDD p w=0.685u l=0.18u
MI0-MU2 net17 A2 XI0-net6 VDD p w=0.68u l=0.18u
MI0-MU1 XI0-net6 net11 VDD VDD p w=0.68u l=0.18u
MU21-MU2 net21 net17 XU21-net6 VDD p w=0.685u l=0.18u
MU21-MU1 XU21-net6 net5 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XNR3D2BWP7T A1 A2 A3 ZN VDD VSS 
M_u6-M_u2 net11 A2 net17 VSS n w=0.5u l=0.18u
MU11-M_u2 net5 net17 net21 VSS n w=0.5u l=0.18u
MI1-M_u2 net5 A3 VSS VSS n w=1u l=0.18u
MU22_0-M_u2 ZN net21 VSS VSS n w=1u l=0.18u
MU22_1-M_u2 ZN net21 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net16 A2 VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net11 A1 VSS VSS n w=1u l=0.18u
MU12-M_u2 net13 net17 VSS VSS n w=0.64u l=0.18u
MI0-MU3 net17 net16 XI0-net16 VSS n w=0.5u l=0.18u
MI0-MU4 XI0-net16 net11 VSS VSS n w=0.5u l=0.18u
MU21-MU3 net21 net13 XU21-net16 VSS n w=0.57u l=0.18u
MU21-MU4 XU21-net16 net5 VSS VSS n w=0.57u l=0.18u
M_u6-M_u3 net11 net16 net17 VDD p w=0.685u l=0.18u
MU11-M_u3 net5 net13 net21 VDD p w=0.865u l=0.18u
MI1-M_u3 net5 A3 VDD VDD p w=1.37u l=0.18u
MU22_0-M_u3 ZN net21 VDD VDD p w=1.37u l=0.18u
MU22_1-M_u3 ZN net21 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net16 A2 VDD VDD p w=0.685u l=0.18u
M_u2-M_u3 net11 A1 VDD VDD p w=1.37u l=0.18u
MU12-M_u3 net13 net17 VDD VDD p w=0.825u l=0.18u
MI0-MU2 net17 A2 XI0-net6 VDD p w=0.685u l=0.18u
MI0-MU1 XI0-net6 net11 VDD VDD p w=1.37u l=0.18u
MU21-MU2 net21 net17 XU21-net6 VDD p w=0.8u l=0.18u
MU21-MU1 XU21-net6 net5 VDD VDD p w=0.935u l=0.18u
.ends
.subckt XNR4D0BWP7T A1 A2 A3 A4 ZN VDD VSS 
MU21-MU3 net24 A1 XU21-net16 VSS n w=0.5u l=0.18u
MU21-MU4 XU21-net16 net32 VSS VSS n w=0.5u l=0.18u
MI21-MU3 net20 A4 XI21-net16 VSS n w=0.5u l=0.18u
MI21-MU4 XI21-net16 net077 VSS VSS n w=0.5u l=0.18u
MI20-MU3 net044 net20 XI20-net16 VSS n w=0.5u l=0.18u
MI20-MU4 XI20-net16 net24 VSS VSS n w=0.5u l=0.18u
MI22-M_u2 net20 net064 net077 VSS n w=0.5u l=0.18u
MI8-M_u2 net24 net30 net32 VSS n w=0.5u l=0.18u
MI17-M_u2 net044 net40 net24 VSS n w=0.5u l=0.18u
MI24-M_u2 net064 A4 VSS VSS n w=0.5u l=0.18u
MI18-M_u2 net32 A2 VSS VSS n w=0.5u l=0.18u
M_u8-M_u2 net30 A1 VSS VSS n w=0.5u l=0.18u
MI23-M_u2 net077 A3 VSS VSS n w=0.5u l=0.18u
MU20-M_u2 ZN net044 VSS VSS n w=0.5u l=0.18u
MU14-M_u2 net40 net20 VSS VSS n w=0.5u l=0.18u
MU21-MU2 net24 net30 XU21-net6 VDD p w=0.685u l=0.18u
MU21-MU1 XU21-net6 net32 VDD VDD p w=0.685u l=0.18u
MI21-MU2 net20 net064 XI21-net6 VDD p w=0.685u l=0.18u
MI21-MU1 XI21-net6 net077 VDD VDD p w=0.685u l=0.18u
MI20-MU2 net044 net40 XI20-net6 VDD p w=0.685u l=0.18u
MI20-MU1 XI20-net6 net24 VDD VDD p w=0.685u l=0.18u
MI22-M_u3 net20 A4 net077 VDD p w=0.685u l=0.18u
MI8-M_u3 net24 A1 net32 VDD p w=0.685u l=0.18u
MI17-M_u3 net044 net20 net24 VDD p w=0.685u l=0.18u
MI24-M_u3 net064 A4 VDD VDD p w=0.685u l=0.18u
MI18-M_u3 net32 A2 VDD VDD p w=0.685u l=0.18u
M_u8-M_u3 net30 A1 VDD VDD p w=0.685u l=0.18u
MI23-M_u3 net077 A3 VDD VDD p w=0.685u l=0.18u
MU20-M_u3 ZN net044 VDD VDD p w=0.685u l=0.18u
MU14-M_u3 net40 net20 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XNR4D1BWP7T A1 A2 A3 A4 ZN VDD VSS 
MU21-MU3 net24 A1 XU21-net16 VSS n w=0.5u l=0.18u
MU21-MU4 XU21-net16 net32 VSS VSS n w=0.5u l=0.18u
MI21-MU3 net20 A4 XI21-net16 VSS n w=0.5u l=0.18u
MI21-MU4 XI21-net16 net077 VSS VSS n w=0.5u l=0.18u
MI20-MU3 net044 net20 XI20-net16 VSS n w=0.5u l=0.18u
MI20-MU4 XI20-net16 net24 VSS VSS n w=0.5u l=0.18u
MI22-M_u2 net20 net064 net077 VSS n w=0.5u l=0.18u
MI8-M_u2 net24 net30 net32 VSS n w=0.5u l=0.18u
MI17-M_u2 net044 net40 net24 VSS n w=0.5u l=0.18u
MI24-M_u2 net064 A4 VSS VSS n w=0.5u l=0.18u
MI18-M_u2 net32 A2 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net30 A1 VSS VSS n w=0.5u l=0.18u
MI23-M_u2 net077 A3 VSS VSS n w=1u l=0.18u
MU20-M_u2 ZN net044 VSS VSS n w=1u l=0.18u
MU14-M_u2 net40 net20 VSS VSS n w=0.5u l=0.18u
MU21-MU2 net24 net30 XU21-net6 VDD p w=0.685u l=0.18u
MU21-MU1 XU21-net6 net32 VDD VDD p w=0.685u l=0.18u
MI21-MU2 net20 net064 XI21-net6 VDD p w=0.685u l=0.18u
MI21-MU1 XI21-net6 net077 VDD VDD p w=0.685u l=0.18u
MI20-MU2 net044 net40 XI20-net6 VDD p w=0.685u l=0.18u
MI20-MU1 XI20-net6 net24 VDD VDD p w=0.685u l=0.18u
MI22-M_u3 net20 A4 net077 VDD p w=0.685u l=0.18u
MI8-M_u3 net24 A1 net32 VDD p w=0.685u l=0.18u
MI17-M_u3 net044 net20 net24 VDD p w=0.685u l=0.18u
MI24-M_u3 net064 A4 VDD VDD p w=0.685u l=0.18u
MI18-M_u3 net32 A2 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net30 A1 VDD VDD p w=0.685u l=0.18u
MI23-M_u3 net077 A3 VDD VDD p w=1.37u l=0.18u
MU20-M_u3 ZN net044 VDD VDD p w=1.31u l=0.18u
MU14-M_u3 net40 net20 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XNR4D2BWP7T A1 A2 A3 A4 ZN VDD VSS 
MU21-MU3 net24 A1 XU21-net16 VSS n w=0.5u l=0.18u
MU21-MU4 XU21-net16 net32 VSS VSS n w=0.5u l=0.18u
MI21-MU3 net20 A4 XI21-net16 VSS n w=0.5u l=0.18u
MI21-MU4 XI21-net16 net077 VSS VSS n w=0.5u l=0.18u
MI20-MU3 net044 net20 XI20-net16 VSS n w=0.5u l=0.18u
MI20-MU4 XI20-net16 net24 VSS VSS n w=0.5u l=0.18u
MI22-M_u2 net20 net064 net077 VSS n w=0.5u l=0.18u
MI8-M_u2 net24 net30 net32 VSS n w=0.5u l=0.18u
MI17-M_u2 net044 net40 net24 VSS n w=0.5u l=0.18u
MI24-M_u2 net064 A4 VSS VSS n w=0.5u l=0.18u
MI18-M_u2 net32 A2 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net30 A1 VSS VSS n w=0.5u l=0.18u
MI23-M_u2 net077 A3 VSS VSS n w=1u l=0.18u
MU20_0-M_u2 ZN net044 VSS VSS n w=1u l=0.18u
MU20_1-M_u2 ZN net044 VSS VSS n w=1u l=0.18u
MU14-M_u2 net40 net20 VSS VSS n w=0.5u l=0.18u
MU21-MU2 net24 net30 XU21-net6 VDD p w=0.685u l=0.18u
MU21-MU1 XU21-net6 net32 VDD VDD p w=0.685u l=0.18u
MI21-MU2 net20 net064 XI21-net6 VDD p w=0.685u l=0.18u
MI21-MU1 XI21-net6 net077 VDD VDD p w=0.685u l=0.18u
MI20-MU2 net044 net40 XI20-net6 VDD p w=0.685u l=0.18u
MI20-MU1 XI20-net6 net24 VDD VDD p w=0.685u l=0.18u
MI22-M_u3 net20 A4 net077 VDD p w=0.685u l=0.18u
MI8-M_u3 net24 A1 net32 VDD p w=0.685u l=0.18u
MI17-M_u3 net044 net20 net24 VDD p w=0.685u l=0.18u
MI24-M_u3 net064 A4 VDD VDD p w=0.685u l=0.18u
MI18-M_u3 net32 A2 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net30 A1 VDD VDD p w=0.685u l=0.18u
MI23-M_u3 net077 A3 VDD VDD p w=1.37u l=0.18u
MU20_0-M_u3 ZN net044 VDD VDD p w=1.37u l=0.18u
MU20_1-M_u3 ZN net044 VDD VDD p w=1.37u l=0.18u
MU14-M_u3 net40 net20 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XOR2D0BWP7T A1 A2 Z VDD VSS 
M_u6-M_u2 net4 net10 net14 VSS n w=0.5u l=0.18u
MI3-M_u2 net6 A1 net14 VSS n w=0.5u l=0.18u
MI1-M_u2 net4 A2 VSS VSS n w=0.5u l=0.18u
M_u5-M_u2 net6 net4 VSS VSS n w=0.5u l=0.18u
M_u4-M_u2 Z net14 VSS VSS n w=0.5u l=0.18u
MI2-M_u2 net10 A1 VSS VSS n w=0.5u l=0.18u
M_u6-M_u3 net4 A1 net14 VDD p w=0.685u l=0.18u
MI3-M_u3 net6 net10 net14 VDD p w=0.685u l=0.18u
MI1-M_u3 net4 A2 VDD VDD p w=0.685u l=0.18u
M_u5-M_u3 net6 net4 VDD VDD p w=0.685u l=0.18u
M_u4-M_u3 Z net14 VDD VDD p w=0.685u l=0.18u
MI2-M_u3 net10 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XOR2D1BWP7T A1 A2 Z VDD VSS 
M_u6-M_u2 net4 net10 net14 VSS n w=0.5u l=0.18u
MI0-M_u2 net6 A1 net14 VSS n w=0.5u l=0.18u
M_u2-M_u2 net4 A2 VSS VSS n w=1u l=0.18u
M_u5-M_u2 net6 net4 VSS VSS n w=0.5u l=0.18u
M_u4-M_u2 Z net14 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net10 A1 VSS VSS n w=0.685u l=0.18u
M_u6-M_u3 net4 A1 net14 VDD p w=0.685u l=0.18u
MI0-M_u3 net6 net10 net14 VDD p w=0.685u l=0.18u
M_u2-M_u3 net4 A2 VDD VDD p w=1.37u l=0.18u
M_u5-M_u3 net6 net4 VDD VDD p w=0.685u l=0.18u
M_u4-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net10 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XOR2D2BWP7T A1 A2 Z VDD VSS 
M_u6-M_u2 net4 net10 net14 VSS n w=0.81u l=0.18u
MI0-M_u2 net6 A1 net14 VSS n w=0.81u l=0.18u
M_u2-M_u2 net4 A2 VSS VSS n w=1u l=0.18u
M_u5-M_u2 net6 net4 VSS VSS n w=1u l=0.18u
M_u4_0-M_u2 Z net14 VSS VSS n w=1u l=0.18u
M_u4_1-M_u2 Z net14 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net10 A1 VSS VSS n w=0.5u l=0.18u
M_u6-M_u3 net4 A1 net14 VDD p w=0.73u l=0.18u
MI0-M_u3 net6 net10 net14 VDD p w=0.73u l=0.18u
M_u2-M_u3 net4 A2 VDD VDD p w=1.37u l=0.18u
M_u5-M_u3 net6 net4 VDD VDD p w=1.37u l=0.18u
M_u4_0-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
M_u4_1-M_u3 Z net14 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net10 A1 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XOR3D0BWP7T A1 A2 A3 Z VDD VSS 
M_u6-M_u2 net19 net17 net25 VSS n w=0.5u l=0.18u
MU18-M_u2 net13 net25 net29 VSS n w=0.5u l=0.18u
MI1-M_u2 Z net29 VSS VSS n w=0.5u l=0.18u
MI3-M_u2 net13 A3 VSS VSS n w=0.5u l=0.18u
MI4-M_u2 net17 A2 VSS VSS n w=0.5u l=0.18u
MI2-M_u2 net19 A1 VSS VSS n w=0.5u l=0.18u
M_u4-M_u2 net21 net25 VSS VSS n w=0.5u l=0.18u
MU33-MU3 net29 net21 XU33-net16 VSS n w=0.5u l=0.18u
MU33-MU4 XU33-net16 net13 VSS VSS n w=0.5u l=0.18u
MI5-MU3 net25 A2 XI5-net16 VSS n w=0.5u l=0.18u
MI5-MU4 XI5-net16 net19 VSS VSS n w=0.5u l=0.18u
M_u6-M_u3 net19 A2 net25 VDD p w=0.685u l=0.18u
MU18-M_u3 net13 net21 net29 VDD p w=0.685u l=0.18u
MI1-M_u3 Z net29 VDD VDD p w=0.685u l=0.18u
MI3-M_u3 net13 A3 VDD VDD p w=0.685u l=0.18u
MI4-M_u3 net17 A2 VDD VDD p w=0.685u l=0.18u
MI2-M_u3 net19 A1 VDD VDD p w=0.685u l=0.18u
M_u4-M_u3 net21 net25 VDD VDD p w=0.685u l=0.18u
MU33-MU2 net29 net25 XU33-net6 VDD p w=0.685u l=0.18u
MU33-MU1 XU33-net6 net13 VDD VDD p w=0.685u l=0.18u
MI5-MU2 net25 net17 XI5-net6 VDD p w=0.685u l=0.18u
MI5-MU1 XI5-net6 net19 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XOR3D1BWP7T A1 A2 A3 Z VDD VSS 
M_u6-M_u2 net19 net17 net25 VSS n w=0.5u l=0.18u
MU18-M_u2 net13 net25 net29 VSS n w=0.5u l=0.18u
MU13-M_u2 net13 A3 VSS VSS n w=1u l=0.18u
MU14-M_u2 Z net29 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net17 A2 VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net19 A1 VSS VSS n w=1u l=0.18u
M_u4-M_u2 net21 net25 VSS VSS n w=0.5u l=0.18u
MU33-MU3 net29 net21 XU33-net16 VSS n w=0.5u l=0.18u
MU33-MU4 XU33-net16 net13 VSS VSS n w=0.5u l=0.18u
MI0-MU3 net25 A2 XI0-net16 VSS n w=0.5u l=0.18u
MI0-MU4 XI0-net16 net19 VSS VSS n w=0.5u l=0.18u
M_u6-M_u3 net19 A2 net25 VDD p w=0.685u l=0.18u
MU18-M_u3 net13 net21 net29 VDD p w=0.685u l=0.18u
MU13-M_u3 net13 A3 VDD VDD p w=1.37u l=0.18u
MU14-M_u3 Z net29 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net17 A2 VDD VDD p w=0.685u l=0.18u
M_u2-M_u3 net19 A1 VDD VDD p w=1.37u l=0.18u
M_u4-M_u3 net21 net25 VDD VDD p w=0.685u l=0.18u
MU33-MU2 net29 net25 XU33-net6 VDD p w=0.685u l=0.18u
MU33-MU1 XU33-net6 net13 VDD VDD p w=0.685u l=0.18u
MI0-MU2 net25 net17 XI0-net6 VDD p w=0.685u l=0.18u
MI0-MU1 XI0-net6 net19 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XOR3D2BWP7T A1 A2 A3 Z VDD VSS 
M_u6-M_u2 net19 net17 net25 VSS n w=0.5u l=0.18u
MU18-M_u2 net13 net25 net032 VSS n w=0.5u l=0.18u
MU13-M_u2 net13 A3 VSS VSS n w=1u l=0.18u
MU14_0-M_u2 Z net032 VSS VSS n w=1u l=0.18u
MU14_1-M_u2 Z net032 VSS VSS n w=1u l=0.18u
M_u8-M_u2 net17 A2 VSS VSS n w=0.5u l=0.18u
M_u2-M_u2 net19 A1 VSS VSS n w=1u l=0.18u
M_u4-M_u2 net21 net25 VSS VSS n w=0.5u l=0.18u
MU33-MU3 net032 net21 XU33-net16 VSS n w=0.5u l=0.18u
MU33-MU4 XU33-net16 net13 VSS VSS n w=0.57u l=0.18u
MI0-MU3 net25 A2 XI0-net16 VSS n w=0.5u l=0.18u
MI0-MU4 XI0-net16 net19 VSS VSS n w=0.5u l=0.18u
M_u6-M_u3 net19 A2 net25 VDD p w=0.74u l=0.18u
MU18-M_u3 net13 net21 net032 VDD p w=0.71u l=0.18u
MU13-M_u3 net13 A3 VDD VDD p w=1.37u l=0.18u
MU14_0-M_u3 Z net032 VDD VDD p w=1.37u l=0.18u
MU14_1-M_u3 Z net032 VDD VDD p w=1.37u l=0.18u
M_u8-M_u3 net17 A2 VDD VDD p w=0.685u l=0.18u
M_u2-M_u3 net19 A1 VDD VDD p w=1.37u l=0.18u
M_u4-M_u3 net21 net25 VDD VDD p w=0.685u l=0.18u
MU33-MU2 net032 net25 XU33-net6 VDD p w=0.685u l=0.18u
MU33-MU1 XU33-net6 net13 VDD VDD p w=1.37u l=0.18u
MI0-MU2 net25 net17 XI0-net6 VDD p w=0.74u l=0.18u
MI0-MU1 XI0-net6 net19 VDD VDD p w=1.37u l=0.18u
.ends
.subckt XOR4D0BWP7T A1 A2 A3 A4 Z VDD VSS 
MI30-M_u2 net61 net59 VSS VSS n w=0.5u l=0.18u
MI26-M_u2 net48 A4 VSS VSS n w=0.5u l=0.18u
MI18-M_u2 net46 A2 VSS VSS n w=0.5u l=0.18u
MI27-M_u2 net44 A1 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net054 A3 VSS VSS n w=0.5u l=0.18u
MI29-M_u2 Z net63 VSS VSS n w=0.5u l=0.18u
MI24-M_u2 net59 net48 net054 VSS n w=0.5u l=0.18u
MI25-M_u2 net55 net44 net46 VSS n w=0.5u l=0.18u
MI23-M_u2 net63 net59 net55 VSS n w=0.5u l=0.18u
MI21-MU3 net59 A4 XI21-net16 VSS n w=0.5u l=0.18u
MI21-MU4 XI21-net16 net054 VSS VSS n w=0.5u l=0.18u
MI22-MU3 net63 net61 XI22-net16 VSS n w=0.5u l=0.18u
MI22-MU4 XI22-net16 net55 VSS VSS n w=0.5u l=0.18u
MU21-MU3 net55 A1 XU21-net16 VSS n w=0.5u l=0.18u
MU21-MU4 XU21-net16 net46 VSS VSS n w=0.5u l=0.18u
MI30-M_u3 net61 net59 VDD VDD p w=0.685u l=0.18u
MI26-M_u3 net48 A4 VDD VDD p w=0.685u l=0.18u
MI18-M_u3 net46 A2 VDD VDD p w=0.685u l=0.18u
MI27-M_u3 net44 A1 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net054 A3 VDD VDD p w=0.685u l=0.18u
MI29-M_u3 Z net63 VDD VDD p w=0.685u l=0.18u
MI24-M_u3 net59 A4 net054 VDD p w=0.685u l=0.18u
MI25-M_u3 net55 A1 net46 VDD p w=0.685u l=0.18u
MI23-M_u3 net63 net61 net55 VDD p w=0.685u l=0.18u
MI21-MU2 net59 net48 XI21-net6 VDD p w=0.685u l=0.18u
MI21-MU1 XI21-net6 net054 VDD VDD p w=0.685u l=0.18u
MI22-MU2 net63 net59 XI22-net6 VDD p w=0.685u l=0.18u
MI22-MU1 XI22-net6 net55 VDD VDD p w=0.685u l=0.18u
MU21-MU2 net55 net44 XU21-net6 VDD p w=0.685u l=0.18u
MU21-MU1 XU21-net6 net46 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XOR4D1BWP7T A1 A2 A3 A4 Z VDD VSS 
MI30-M_u2 net61 net59 VSS VSS n w=0.5u l=0.18u
MI26-M_u2 net48 A4 VSS VSS n w=0.5u l=0.18u
MI18-M_u2 net46 A2 VSS VSS n w=1u l=0.18u
MI27-M_u2 net44 A1 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net054 A3 VSS VSS n w=1u l=0.18u
MI29-M_u2 Z net63 VSS VSS n w=1u l=0.18u
MI24-M_u2 net59 net48 net054 VSS n w=0.5u l=0.18u
MI25-M_u2 net55 net44 net46 VSS n w=0.5u l=0.18u
MI23-M_u2 net63 net59 net55 VSS n w=0.5u l=0.18u
MI21-MU3 net59 A4 XI21-net16 VSS n w=0.5u l=0.18u
MI21-MU4 XI21-net16 net054 VSS VSS n w=0.5u l=0.18u
MI22-MU3 net63 net61 XI22-net16 VSS n w=0.5u l=0.18u
MI22-MU4 XI22-net16 net55 VSS VSS n w=0.5u l=0.18u
MU21-MU3 net55 A1 XU21-net16 VSS n w=0.5u l=0.18u
MU21-MU4 XU21-net16 net46 VSS VSS n w=0.5u l=0.18u
MI30-M_u3 net61 net59 VDD VDD p w=0.685u l=0.18u
MI26-M_u3 net48 A4 VDD VDD p w=0.685u l=0.18u
MI18-M_u3 net46 A2 VDD VDD p w=1.37u l=0.18u
MI27-M_u3 net44 A1 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net054 A3 VDD VDD p w=1.37u l=0.18u
MI29-M_u3 Z net63 VDD VDD p w=1.31u l=0.18u
MI24-M_u3 net59 A4 net054 VDD p w=0.685u l=0.18u
MI25-M_u3 net55 A1 net46 VDD p w=0.685u l=0.18u
MI23-M_u3 net63 net61 net55 VDD p w=0.685u l=0.18u
MI21-MU2 net59 net48 XI21-net6 VDD p w=0.685u l=0.18u
MI21-MU1 XI21-net6 net054 VDD VDD p w=0.685u l=0.18u
MI22-MU2 net63 net59 XI22-net6 VDD p w=0.685u l=0.18u
MI22-MU1 XI22-net6 net55 VDD VDD p w=0.685u l=0.18u
MU21-MU2 net55 net44 XU21-net6 VDD p w=0.685u l=0.18u
MU21-MU1 XU21-net6 net46 VDD VDD p w=0.685u l=0.18u
.ends
.subckt XOR4D2BWP7T A1 A2 A3 A4 Z VDD VSS 
MI30-M_u2 net61 net59 VSS VSS n w=0.5u l=0.18u
MI26-M_u2 net48 A4 VSS VSS n w=0.5u l=0.18u
MI18-M_u2 net46 A2 VSS VSS n w=1u l=0.18u
MI27-M_u2 net44 A1 VSS VSS n w=0.5u l=0.18u
MI28-M_u2 net054 A3 VSS VSS n w=1u l=0.18u
MI29_0-M_u2 Z net63 VSS VSS n w=1u l=0.18u
MI29_1-M_u2 Z net63 VSS VSS n w=1u l=0.18u
MI24-M_u2 net59 net48 net054 VSS n w=0.5u l=0.18u
MI25-M_u2 net55 net44 net46 VSS n w=0.5u l=0.18u
MI23-M_u2 net63 net59 net55 VSS n w=0.5u l=0.18u
MI21-MU3 net59 A4 XI21-net16 VSS n w=0.5u l=0.18u
MI21-MU4 XI21-net16 net054 VSS VSS n w=0.5u l=0.18u
MI22-MU3 net63 net61 XI22-net16 VSS n w=0.5u l=0.18u
MI22-MU4 XI22-net16 net55 VSS VSS n w=0.5u l=0.18u
MU21-MU3 net55 A1 XU21-net16 VSS n w=0.5u l=0.18u
MU21-MU4 XU21-net16 net46 VSS VSS n w=0.5u l=0.18u
MI30-M_u3 net61 net59 VDD VDD p w=0.685u l=0.18u
MI26-M_u3 net48 A4 VDD VDD p w=0.685u l=0.18u
MI18-M_u3 net46 A2 VDD VDD p w=1.37u l=0.18u
MI27-M_u3 net44 A1 VDD VDD p w=0.685u l=0.18u
MI28-M_u3 net054 A3 VDD VDD p w=1.37u l=0.18u
MI29_0-M_u3 Z net63 VDD VDD p w=1.37u l=0.18u
MI29_1-M_u3 Z net63 VDD VDD p w=1.37u l=0.18u
MI24-M_u3 net59 A4 net054 VDD p w=0.685u l=0.18u
MI25-M_u3 net55 A1 net46 VDD p w=0.685u l=0.18u
MI23-M_u3 net63 net61 net55 VDD p w=0.685u l=0.18u
MI21-MU2 net59 net48 XI21-net6 VDD p w=0.685u l=0.18u
MI21-MU1 XI21-net6 net054 VDD VDD p w=0.685u l=0.18u
MI22-MU2 net63 net59 XI22-net6 VDD p w=0.685u l=0.18u
MI22-MU1 XI22-net6 net55 VDD VDD p w=0.685u l=0.18u
MU21-MU2 net55 net44 XU21-net6 VDD p w=0.685u l=0.18u
MU21-MU1 XU21-net6 net46 VDD VDD p w=0.685u l=0.18u
.ends
